magic
tech sky130A
magscale 1 2
timestamp 1647613226
<< metal1 >>
rect 201494 703332 201500 703384
rect 201552 703372 201558 703384
rect 202782 703372 202788 703384
rect 201552 703344 202788 703372
rect 201552 703332 201558 703344
rect 202782 703332 202788 703344
rect 202840 703332 202846 703384
rect 77938 703264 77944 703316
rect 77996 703304 78002 703316
rect 267642 703304 267648 703316
rect 77996 703276 267648 703304
rect 77996 703264 78002 703276
rect 267642 703264 267648 703276
rect 267700 703264 267706 703316
rect 95142 703196 95148 703248
rect 95200 703236 95206 703248
rect 332502 703236 332508 703248
rect 95200 703208 332508 703236
rect 95200 703196 95206 703208
rect 332502 703196 332508 703208
rect 332560 703196 332566 703248
rect 109678 703128 109684 703180
rect 109736 703168 109742 703180
rect 348786 703168 348792 703180
rect 109736 703140 348792 703168
rect 109736 703128 109742 703140
rect 348786 703128 348792 703140
rect 348844 703128 348850 703180
rect 111058 703060 111064 703112
rect 111116 703100 111122 703112
rect 397454 703100 397460 703112
rect 111116 703072 397460 703100
rect 111116 703060 111122 703072
rect 397454 703060 397460 703072
rect 397512 703060 397518 703112
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 76558 702992 76564 703044
rect 76616 703032 76622 703044
rect 364978 703032 364984 703044
rect 76616 703004 364984 703032
rect 76616 702992 76622 703004
rect 364978 702992 364984 703004
rect 365036 702992 365042 703044
rect 104802 702924 104808 702976
rect 104860 702964 104866 702976
rect 413646 702964 413652 702976
rect 104860 702936 413652 702964
rect 104860 702924 104866 702936
rect 413646 702924 413652 702936
rect 413704 702924 413710 702976
rect 115842 702856 115848 702908
rect 115900 702896 115906 702908
rect 462314 702896 462320 702908
rect 115900 702868 462320 702896
rect 115900 702856 115906 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 75178 702788 75184 702840
rect 75236 702828 75242 702840
rect 429194 702828 429200 702840
rect 75236 702800 429200 702828
rect 75236 702788 75242 702800
rect 429194 702788 429200 702800
rect 429252 702828 429258 702840
rect 429838 702828 429844 702840
rect 429252 702800 429844 702828
rect 429252 702788 429258 702800
rect 429838 702788 429844 702800
rect 429896 702788 429902 702840
rect 117222 702720 117228 702772
rect 117280 702760 117286 702772
rect 478506 702760 478512 702772
rect 117280 702732 478512 702760
rect 117280 702720 117286 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 113082 702652 113088 702704
rect 113140 702692 113146 702704
rect 453942 702692 453948 702704
rect 113140 702664 453948 702692
rect 113140 702652 113146 702664
rect 453942 702652 453948 702664
rect 454000 702652 454006 702704
rect 492582 702652 492588 702704
rect 492640 702692 492646 702704
rect 494790 702692 494796 702704
rect 492640 702664 494796 702692
rect 492640 702652 492646 702664
rect 494790 702652 494796 702664
rect 494848 702652 494854 702704
rect 79318 702584 79324 702636
rect 79376 702624 79382 702636
rect 527174 702624 527180 702636
rect 79376 702596 527180 702624
rect 79376 702584 79382 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 108942 702516 108948 702568
rect 109000 702556 109006 702568
rect 511902 702556 511908 702568
rect 109000 702528 511908 702556
rect 109000 702516 109006 702528
rect 511902 702516 511908 702528
rect 511960 702516 511966 702568
rect 550542 702516 550548 702568
rect 550600 702556 550606 702568
rect 559650 702556 559656 702568
rect 550600 702528 559656 702556
rect 550600 702516 550606 702528
rect 559650 702516 559656 702528
rect 559708 702516 559714 702568
rect 68922 702448 68928 702500
rect 68980 702488 68986 702500
rect 543458 702488 543464 702500
rect 68980 702460 543464 702488
rect 68980 702448 68986 702460
rect 543458 702448 543464 702460
rect 543516 702448 543522 702500
rect 364978 701700 364984 701752
rect 365036 701740 365042 701752
rect 483658 701740 483664 701752
rect 365036 701712 483664 701740
rect 365036 701700 365042 701712
rect 483658 701700 483664 701712
rect 483716 701700 483722 701752
rect 71038 700340 71044 700392
rect 71096 700380 71102 700392
rect 154114 700380 154120 700392
rect 71096 700352 154120 700380
rect 71096 700340 71102 700352
rect 154114 700340 154120 700352
rect 154172 700340 154178 700392
rect 162118 700340 162124 700392
rect 162176 700380 162182 700392
rect 218974 700380 218980 700392
rect 162176 700352 218980 700380
rect 162176 700340 162182 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 62022 700272 62028 700324
rect 62080 700312 62086 700324
rect 235166 700312 235172 700324
rect 62080 700284 235172 700312
rect 62080 700272 62086 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 238018 700272 238024 700324
rect 238076 700312 238082 700324
rect 283834 700312 283840 700324
rect 238076 700284 283840 700312
rect 238076 700272 238082 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 450538 700272 450544 700324
rect 450596 700312 450602 700324
rect 453942 700312 453948 700324
rect 450596 700284 453948 700312
rect 450596 700272 450602 700284
rect 453942 700272 453948 700284
rect 454000 700312 454006 700324
rect 492582 700312 492588 700324
rect 454000 700284 492588 700312
rect 454000 700272 454006 700284
rect 492582 700272 492588 700284
rect 492640 700272 492646 700324
rect 511902 700272 511908 700324
rect 511960 700312 511966 700324
rect 550542 700312 550548 700324
rect 511960 700284 550548 700312
rect 511960 700272 511966 700284
rect 550542 700272 550548 700284
rect 550600 700272 550606 700324
rect 511258 699660 511264 699712
rect 511316 699700 511322 699712
rect 511902 699700 511908 699712
rect 511316 699672 511908 699700
rect 511316 699660 511322 699672
rect 511902 699660 511908 699672
rect 511960 699660 511966 699712
rect 24302 698912 24308 698964
rect 24360 698952 24366 698964
rect 106274 698952 106280 698964
rect 24360 698924 106280 698952
rect 24360 698912 24366 698924
rect 106274 698912 106280 698924
rect 106332 698912 106338 698964
rect 57882 697552 57888 697604
rect 57940 697592 57946 697604
rect 170306 697592 170312 697604
rect 57940 697564 170312 697592
rect 57940 697552 57946 697564
rect 170306 697552 170312 697564
rect 170364 697552 170370 697604
rect 69014 696940 69020 696992
rect 69072 696980 69078 696992
rect 580166 696980 580172 696992
rect 69072 696952 580172 696980
rect 69072 696940 69078 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 159358 683136 159364 683188
rect 159416 683176 159422 683188
rect 580166 683176 580172 683188
rect 159416 683148 580172 683176
rect 159416 683136 159422 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 15838 670732 15844 670744
rect 3568 670704 15844 670732
rect 3568 670692 3574 670704
rect 15838 670692 15844 670704
rect 15896 670692 15902 670744
rect 90358 670692 90364 670744
rect 90416 670732 90422 670744
rect 580902 670732 580908 670744
rect 90416 670704 580908 670732
rect 90416 670692 90422 670704
rect 580902 670692 580908 670704
rect 580960 670692 580966 670744
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 11698 656928 11704 656940
rect 3568 656900 11704 656928
rect 3568 656888 3574 656900
rect 11698 656888 11704 656900
rect 11756 656888 11762 656940
rect 3510 632068 3516 632120
rect 3568 632108 3574 632120
rect 58618 632108 58624 632120
rect 3568 632080 58624 632108
rect 3568 632068 3574 632080
rect 58618 632068 58624 632080
rect 58676 632068 58682 632120
rect 119338 630640 119344 630692
rect 119396 630680 119402 630692
rect 580166 630680 580172 630692
rect 119396 630652 580172 630680
rect 119396 630640 119402 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3510 618264 3516 618316
rect 3568 618304 3574 618316
rect 93118 618304 93124 618316
rect 3568 618276 93124 618304
rect 3568 618264 3574 618276
rect 93118 618264 93124 618276
rect 93176 618264 93182 618316
rect 425698 616088 425704 616140
rect 425756 616128 425762 616140
rect 580166 616128 580172 616140
rect 425756 616100 580172 616128
rect 425756 616088 425762 616100
rect 580166 616088 580172 616100
rect 580224 616088 580230 616140
rect 6914 598204 6920 598256
rect 6972 598244 6978 598256
rect 46842 598244 46848 598256
rect 6972 598216 46848 598244
rect 6972 598204 6978 598216
rect 46842 598204 46848 598216
rect 46900 598204 46906 598256
rect 46842 597524 46848 597576
rect 46900 597564 46906 597576
rect 85574 597564 85580 597576
rect 46900 597536 85580 597564
rect 46900 597524 46906 597536
rect 85574 597524 85580 597536
rect 85632 597524 85638 597576
rect 68830 596776 68836 596828
rect 68888 596816 68894 596828
rect 238018 596816 238024 596828
rect 68888 596788 238024 596816
rect 68888 596776 68894 596788
rect 238018 596776 238024 596788
rect 238076 596776 238082 596828
rect 3418 595416 3424 595468
rect 3476 595456 3482 595468
rect 42794 595456 42800 595468
rect 3476 595428 42800 595456
rect 3476 595416 3482 595428
rect 42794 595416 42800 595428
rect 42852 595416 42858 595468
rect 42794 594804 42800 594856
rect 42852 594844 42858 594856
rect 44082 594844 44088 594856
rect 42852 594816 44088 594844
rect 42852 594804 42858 594816
rect 44082 594804 44088 594816
rect 44140 594844 44146 594856
rect 71866 594844 71872 594856
rect 44140 594816 71872 594844
rect 44140 594804 44146 594816
rect 71866 594804 71872 594816
rect 71924 594804 71930 594856
rect 3510 594056 3516 594108
rect 3568 594096 3574 594108
rect 106458 594096 106464 594108
rect 3568 594068 106464 594096
rect 3568 594056 3574 594068
rect 106458 594056 106464 594068
rect 106516 594056 106522 594108
rect 68646 592628 68652 592680
rect 68704 592668 68710 592680
rect 136634 592668 136640 592680
rect 68704 592640 136640 592668
rect 68704 592628 68710 592640
rect 136634 592628 136640 592640
rect 136692 592628 136698 592680
rect 82078 591268 82084 591320
rect 82136 591308 82142 591320
rect 90358 591308 90364 591320
rect 82136 591280 90364 591308
rect 82136 591268 82142 591280
rect 90358 591268 90364 591280
rect 90416 591268 90422 591320
rect 40034 590656 40040 590708
rect 40092 590696 40098 590708
rect 48222 590696 48228 590708
rect 40092 590668 48228 590696
rect 40092 590656 40098 590668
rect 48222 590656 48228 590668
rect 48280 590696 48286 590708
rect 74626 590696 74632 590708
rect 48280 590668 74632 590696
rect 48280 590656 48286 590668
rect 74626 590656 74632 590668
rect 74684 590656 74690 590708
rect 556798 590656 556804 590708
rect 556856 590696 556862 590708
rect 579798 590696 579804 590708
rect 556856 590668 579804 590696
rect 556856 590656 556862 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 11698 588548 11704 588600
rect 11756 588588 11762 588600
rect 87322 588588 87328 588600
rect 11756 588560 87328 588588
rect 11756 588548 11762 588560
rect 87322 588548 87328 588560
rect 87380 588548 87386 588600
rect 88334 588548 88340 588600
rect 88392 588588 88398 588600
rect 117406 588588 117412 588600
rect 88392 588560 117412 588588
rect 88392 588548 88398 588560
rect 117406 588548 117412 588560
rect 117464 588548 117470 588600
rect 103514 586712 103520 586764
rect 103572 586752 103578 586764
rect 104802 586752 104808 586764
rect 103572 586724 104808 586752
rect 103572 586712 103578 586724
rect 104802 586712 104808 586724
rect 104860 586752 104866 586764
rect 131298 586752 131304 586764
rect 104860 586724 131304 586752
rect 104860 586712 104866 586724
rect 131298 586712 131304 586724
rect 131356 586712 131362 586764
rect 85298 586644 85304 586696
rect 85356 586684 85362 586696
rect 113266 586684 113272 586696
rect 85356 586656 113272 586684
rect 85356 586644 85362 586656
rect 113266 586644 113272 586656
rect 113324 586644 113330 586696
rect 49602 586576 49608 586628
rect 49660 586616 49666 586628
rect 79318 586616 79324 586628
rect 49660 586588 79324 586616
rect 49660 586576 49666 586588
rect 79318 586576 79324 586588
rect 79376 586576 79382 586628
rect 91002 586576 91008 586628
rect 91060 586616 91066 586628
rect 123018 586616 123024 586628
rect 91060 586588 123024 586616
rect 91060 586576 91066 586588
rect 123018 586576 123024 586588
rect 123076 586576 123082 586628
rect 52362 586508 52368 586560
rect 52420 586548 52426 586560
rect 84286 586548 84292 586560
rect 52420 586520 84292 586548
rect 52420 586508 52426 586520
rect 84286 586508 84292 586520
rect 84344 586508 84350 586560
rect 94866 586508 94872 586560
rect 94924 586548 94930 586560
rect 128446 586548 128452 586560
rect 94924 586520 128452 586548
rect 94924 586508 94930 586520
rect 128446 586508 128452 586520
rect 128504 586508 128510 586560
rect 112070 585760 112076 585812
rect 112128 585800 112134 585812
rect 162118 585800 162124 585812
rect 112128 585772 162124 585800
rect 112128 585760 112134 585772
rect 162118 585760 162124 585772
rect 162176 585760 162182 585812
rect 93118 585352 93124 585404
rect 93176 585392 93182 585404
rect 95878 585392 95884 585404
rect 93176 585364 95884 585392
rect 93176 585352 93182 585364
rect 95878 585352 95884 585364
rect 95936 585392 95942 585404
rect 115934 585392 115940 585404
rect 95936 585364 115940 585392
rect 95936 585352 95942 585364
rect 115934 585352 115940 585364
rect 115992 585352 115998 585404
rect 61930 585284 61936 585336
rect 61988 585324 61994 585336
rect 80606 585324 80612 585336
rect 61988 585296 80612 585324
rect 61988 585284 61994 585296
rect 80606 585284 80612 585296
rect 80664 585284 80670 585336
rect 95142 585284 95148 585336
rect 95200 585324 95206 585336
rect 120074 585324 120080 585336
rect 95200 585296 120080 585324
rect 95200 585284 95206 585296
rect 120074 585284 120080 585296
rect 120132 585284 120138 585336
rect 50706 585216 50712 585268
rect 50764 585256 50770 585268
rect 76558 585256 76564 585268
rect 50764 585228 76564 585256
rect 50764 585216 50770 585228
rect 76558 585216 76564 585228
rect 76616 585216 76622 585268
rect 87322 585216 87328 585268
rect 87380 585256 87386 585268
rect 87506 585256 87512 585268
rect 87380 585228 87512 585256
rect 87380 585216 87386 585228
rect 87506 585216 87512 585228
rect 87564 585256 87570 585268
rect 118786 585256 118792 585268
rect 87564 585228 118792 585256
rect 87564 585216 87570 585228
rect 118786 585216 118792 585228
rect 118844 585216 118850 585268
rect 49510 585148 49516 585200
rect 49568 585188 49574 585200
rect 78030 585188 78036 585200
rect 49568 585160 78036 585188
rect 49568 585148 49574 585160
rect 78030 585148 78036 585160
rect 78088 585148 78094 585200
rect 97902 585148 97908 585200
rect 97960 585188 97966 585200
rect 131114 585188 131120 585200
rect 97960 585160 131120 585188
rect 97960 585148 97966 585160
rect 131114 585148 131120 585160
rect 131172 585148 131178 585200
rect 88242 584196 88248 584248
rect 88300 584236 88306 584248
rect 105630 584236 105636 584248
rect 88300 584208 105636 584236
rect 88300 584196 88306 584208
rect 105630 584196 105636 584208
rect 105688 584196 105694 584248
rect 98730 584128 98736 584180
rect 98788 584168 98794 584180
rect 101398 584168 101404 584180
rect 98788 584140 101404 584168
rect 98788 584128 98794 584140
rect 101398 584128 101404 584140
rect 101456 584128 101462 584180
rect 77846 584100 77852 584112
rect 64846 584072 77852 584100
rect 39850 583992 39856 584044
rect 39908 584032 39914 584044
rect 64846 584032 64874 584072
rect 77846 584060 77852 584072
rect 77904 584100 77910 584112
rect 79226 584100 79232 584112
rect 77904 584072 79232 584100
rect 77904 584060 77910 584072
rect 79226 584060 79232 584072
rect 79284 584060 79290 584112
rect 99282 584060 99288 584112
rect 99340 584100 99346 584112
rect 129826 584100 129832 584112
rect 99340 584072 129832 584100
rect 99340 584060 99346 584072
rect 129826 584060 129832 584072
rect 129884 584060 129890 584112
rect 39908 584004 64874 584032
rect 39908 583992 39914 584004
rect 66162 583992 66168 584044
rect 66220 584032 66226 584044
rect 70946 584032 70952 584044
rect 66220 584004 70952 584032
rect 66220 583992 66226 584004
rect 70946 583992 70952 584004
rect 71004 583992 71010 584044
rect 96522 583992 96528 584044
rect 96580 584032 96586 584044
rect 110414 584032 110420 584044
rect 96580 584004 110420 584032
rect 96580 583992 96586 584004
rect 110414 583992 110420 584004
rect 110472 583992 110478 584044
rect 56502 583924 56508 583976
rect 56560 583964 56566 583976
rect 70394 583964 70400 583976
rect 56560 583936 70400 583964
rect 56560 583924 56566 583936
rect 70394 583924 70400 583936
rect 70452 583924 70458 583976
rect 101306 583924 101312 583976
rect 101364 583964 101370 583976
rect 116026 583964 116032 583976
rect 101364 583936 116032 583964
rect 101364 583924 101370 583936
rect 116026 583924 116032 583936
rect 116084 583924 116090 583976
rect 41230 583856 41236 583908
rect 41288 583896 41294 583908
rect 73338 583896 73344 583908
rect 41288 583868 73344 583896
rect 41288 583856 41294 583868
rect 73338 583856 73344 583868
rect 73396 583856 73402 583908
rect 101858 583856 101864 583908
rect 101916 583896 101922 583908
rect 113358 583896 113364 583908
rect 101916 583868 113364 583896
rect 101916 583856 101922 583868
rect 113358 583856 113364 583868
rect 113416 583856 113422 583908
rect 59170 583788 59176 583840
rect 59228 583828 59234 583840
rect 96706 583828 96712 583840
rect 59228 583800 96712 583828
rect 59228 583788 59234 583800
rect 96706 583788 96712 583800
rect 96764 583788 96770 583840
rect 104434 583788 104440 583840
rect 104492 583828 104498 583840
rect 125686 583828 125692 583840
rect 104492 583800 125692 583828
rect 104492 583788 104498 583800
rect 125686 583788 125692 583800
rect 125744 583788 125750 583840
rect 70302 583720 70308 583772
rect 70360 583760 70366 583772
rect 83366 583760 83372 583772
rect 70360 583732 83372 583760
rect 70360 583720 70366 583732
rect 83366 583720 83372 583732
rect 83424 583720 83430 583772
rect 88978 583720 88984 583772
rect 89036 583760 89042 583772
rect 102134 583760 102140 583772
rect 89036 583732 102140 583760
rect 89036 583720 89042 583732
rect 102134 583720 102140 583732
rect 102192 583720 102198 583772
rect 105262 583720 105268 583772
rect 105320 583760 105326 583772
rect 114554 583760 114560 583772
rect 105320 583732 114560 583760
rect 105320 583720 105326 583732
rect 114554 583720 114560 583732
rect 114612 583720 114618 583772
rect 59998 582972 60004 583024
rect 60056 583012 60062 583024
rect 71774 583012 71780 583024
rect 60056 582984 71780 583012
rect 60056 582972 60062 582984
rect 71774 582972 71780 582984
rect 71832 582972 71838 583024
rect 102134 582972 102140 583024
rect 102192 583012 102198 583024
rect 121454 583012 121460 583024
rect 102192 582984 121460 583012
rect 102192 582972 102198 582984
rect 121454 582972 121460 582984
rect 121512 582972 121518 583024
rect 92842 582632 92848 582684
rect 92900 582672 92906 582684
rect 109034 582672 109040 582684
rect 92900 582644 109040 582672
rect 92900 582632 92906 582644
rect 109034 582632 109040 582644
rect 109092 582632 109098 582684
rect 83274 582564 83280 582616
rect 83332 582604 83338 582616
rect 110506 582604 110512 582616
rect 83332 582576 110512 582604
rect 83332 582564 83338 582576
rect 110506 582564 110512 582576
rect 110564 582564 110570 582616
rect 54478 582496 54484 582548
rect 54536 582536 54542 582548
rect 76742 582536 76748 582548
rect 54536 582508 76748 582536
rect 54536 582496 54542 582508
rect 76742 582496 76748 582508
rect 76800 582496 76806 582548
rect 91554 582496 91560 582548
rect 91612 582536 91618 582548
rect 120166 582536 120172 582548
rect 91612 582508 120172 582536
rect 91612 582496 91618 582508
rect 120166 582496 120172 582508
rect 120224 582496 120230 582548
rect 57790 582428 57796 582480
rect 57848 582468 57854 582480
rect 84470 582468 84476 582480
rect 57848 582440 84476 582468
rect 57848 582428 57854 582440
rect 84470 582428 84476 582440
rect 84528 582428 84534 582480
rect 89622 582428 89628 582480
rect 89680 582468 89686 582480
rect 122834 582468 122840 582480
rect 89680 582440 122840 582468
rect 89680 582428 89686 582440
rect 122834 582428 122840 582440
rect 122892 582428 122898 582480
rect 14458 582360 14464 582412
rect 14516 582400 14522 582412
rect 107654 582400 107660 582412
rect 14516 582372 107660 582400
rect 14516 582360 14522 582372
rect 107654 582360 107660 582372
rect 107712 582360 107718 582412
rect 68462 581952 68468 582004
rect 68520 581992 68526 582004
rect 71038 581992 71044 582004
rect 68520 581964 71044 581992
rect 68520 581952 68526 581964
rect 71038 581952 71044 581964
rect 71096 581952 71102 582004
rect 65518 581748 65524 581800
rect 65576 581788 65582 581800
rect 75454 581788 75460 581800
rect 65576 581760 75460 581788
rect 65576 581748 65582 581760
rect 75454 581748 75460 581760
rect 75512 581748 75518 581800
rect 72234 581680 72240 581732
rect 72292 581680 72298 581732
rect 78674 581720 78680 581732
rect 74506 581692 78680 581720
rect 53098 581204 53104 581256
rect 53156 581244 53162 581256
rect 67634 581244 67640 581256
rect 53156 581216 67640 581244
rect 53156 581204 53162 581216
rect 67634 581204 67640 581216
rect 67692 581204 67698 581256
rect 50798 581136 50804 581188
rect 50856 581176 50862 581188
rect 72252 581176 72280 581680
rect 50856 581148 72280 581176
rect 50856 581136 50862 581148
rect 48038 581068 48044 581120
rect 48096 581108 48102 581120
rect 74506 581108 74534 581692
rect 78674 581680 78680 581692
rect 78732 581680 78738 581732
rect 90266 581680 90272 581732
rect 90324 581720 90330 581732
rect 90324 581692 93854 581720
rect 90324 581680 90330 581692
rect 48096 581080 74534 581108
rect 48096 581068 48102 581080
rect 35802 581000 35808 581052
rect 35860 581040 35866 581052
rect 65518 581040 65524 581052
rect 35860 581012 65524 581040
rect 35860 581000 35866 581012
rect 65518 581000 65524 581012
rect 65576 581000 65582 581052
rect 93826 581040 93854 581692
rect 100570 581680 100576 581732
rect 100628 581720 100634 581732
rect 100628 581692 103514 581720
rect 100628 581680 100634 581692
rect 103486 581176 103514 581692
rect 104986 581680 104992 581732
rect 105044 581720 105050 581732
rect 108942 581720 108948 581732
rect 105044 581692 108948 581720
rect 105044 581680 105050 581692
rect 108942 581680 108948 581692
rect 109000 581680 109006 581732
rect 117314 581176 117320 581188
rect 103486 581148 117320 581176
rect 117314 581136 117320 581148
rect 117372 581136 117378 581188
rect 108942 581068 108948 581120
rect 109000 581108 109006 581120
rect 127066 581108 127072 581120
rect 109000 581080 127072 581108
rect 109000 581068 109006 581080
rect 127066 581068 127072 581080
rect 127124 581068 127130 581120
rect 122926 581040 122932 581052
rect 93826 581012 122932 581040
rect 122926 581000 122932 581012
rect 122984 581000 122990 581052
rect 65518 579640 65524 579692
rect 65576 579680 65582 579692
rect 68646 579680 68652 579692
rect 65576 579652 68652 579680
rect 65576 579640 65582 579652
rect 68646 579640 68652 579652
rect 68704 579640 68710 579692
rect 108206 579640 108212 579692
rect 108264 579680 108270 579692
rect 111794 579680 111800 579692
rect 108264 579652 111800 579680
rect 108264 579640 108270 579652
rect 111794 579640 111800 579652
rect 111852 579640 111858 579692
rect 64598 578280 64604 578332
rect 64656 578320 64662 578332
rect 67726 578320 67732 578332
rect 64656 578292 67732 578320
rect 64656 578280 64662 578292
rect 67726 578280 67732 578292
rect 67784 578280 67790 578332
rect 108850 578280 108856 578332
rect 108908 578320 108914 578332
rect 133138 578320 133144 578332
rect 108908 578292 133144 578320
rect 108908 578280 108914 578292
rect 133138 578280 133144 578292
rect 133196 578280 133202 578332
rect 53650 578212 53656 578264
rect 53708 578252 53714 578264
rect 67634 578252 67640 578264
rect 53708 578224 67640 578252
rect 53708 578212 53714 578224
rect 67634 578212 67640 578224
rect 67692 578212 67698 578264
rect 108942 578212 108948 578264
rect 109000 578252 109006 578264
rect 135254 578252 135260 578264
rect 109000 578224 135260 578252
rect 109000 578212 109006 578224
rect 135254 578212 135260 578224
rect 135312 578212 135318 578264
rect 69106 576988 69112 577040
rect 69164 577028 69170 577040
rect 69750 577028 69756 577040
rect 69164 577000 69756 577028
rect 69164 576988 69170 577000
rect 69750 576988 69756 577000
rect 69808 576988 69814 577040
rect 64506 576852 64512 576904
rect 64564 576892 64570 576904
rect 67634 576892 67640 576904
rect 64564 576864 67640 576892
rect 64564 576852 64570 576864
rect 67634 576852 67640 576864
rect 67692 576852 67698 576904
rect 105630 576104 105636 576156
rect 105688 576144 105694 576156
rect 118878 576144 118884 576156
rect 105688 576116 118884 576144
rect 105688 576104 105694 576116
rect 118878 576104 118884 576116
rect 118936 576104 118942 576156
rect 37182 575492 37188 575544
rect 37240 575532 37246 575544
rect 67634 575532 67640 575544
rect 37240 575504 67640 575532
rect 37240 575492 37246 575504
rect 67634 575492 67640 575504
rect 67692 575492 67698 575544
rect 108942 575492 108948 575544
rect 109000 575532 109006 575544
rect 122742 575532 122748 575544
rect 109000 575504 122748 575532
rect 109000 575492 109006 575504
rect 122742 575492 122748 575504
rect 122800 575532 122806 575544
rect 431218 575532 431224 575544
rect 122800 575504 431224 575532
rect 122800 575492 122806 575504
rect 431218 575492 431224 575504
rect 431276 575492 431282 575544
rect 61746 574132 61752 574184
rect 61804 574172 61810 574184
rect 67726 574172 67732 574184
rect 61804 574144 67732 574172
rect 61804 574132 61810 574144
rect 67726 574132 67732 574144
rect 67784 574132 67790 574184
rect 56318 574064 56324 574116
rect 56376 574104 56382 574116
rect 67634 574104 67640 574116
rect 56376 574076 67640 574104
rect 56376 574064 56382 574076
rect 67634 574064 67640 574076
rect 67692 574064 67698 574116
rect 108942 574064 108948 574116
rect 109000 574104 109006 574116
rect 137278 574104 137284 574116
rect 109000 574076 137284 574104
rect 109000 574064 109006 574076
rect 137278 574064 137284 574076
rect 137336 574064 137342 574116
rect 122098 573996 122104 574048
rect 122156 574036 122162 574048
rect 159358 574036 159364 574048
rect 122156 574008 159364 574036
rect 122156 573996 122162 574008
rect 159358 573996 159364 574008
rect 159416 573996 159422 574048
rect 108942 573316 108948 573368
rect 109000 573356 109006 573368
rect 122098 573356 122104 573368
rect 109000 573328 122104 573356
rect 109000 573316 109006 573328
rect 122098 573316 122104 573328
rect 122156 573316 122162 573368
rect 108666 572976 108672 573028
rect 108724 573016 108730 573028
rect 113174 573016 113180 573028
rect 108724 572988 113180 573016
rect 108724 572976 108730 572988
rect 113174 572976 113180 572988
rect 113232 572976 113238 573028
rect 34422 572772 34428 572824
rect 34480 572812 34486 572824
rect 67634 572812 67640 572824
rect 34480 572784 67640 572812
rect 34480 572772 34486 572784
rect 67634 572772 67640 572784
rect 67692 572772 67698 572824
rect 105630 572772 105636 572824
rect 105688 572812 105694 572824
rect 110598 572812 110604 572824
rect 105688 572784 110604 572812
rect 105688 572772 105694 572784
rect 110598 572772 110604 572784
rect 110656 572772 110662 572824
rect 108942 572704 108948 572756
rect 109000 572744 109006 572756
rect 128630 572744 128636 572756
rect 109000 572716 128636 572744
rect 109000 572704 109006 572716
rect 128630 572704 128636 572716
rect 128688 572704 128694 572756
rect 66070 571548 66076 571600
rect 66128 571588 66134 571600
rect 68278 571588 68284 571600
rect 66128 571560 68284 571588
rect 66128 571548 66134 571560
rect 68278 571548 68284 571560
rect 68336 571548 68342 571600
rect 108942 571344 108948 571396
rect 109000 571384 109006 571396
rect 140774 571384 140780 571396
rect 109000 571356 140780 571384
rect 109000 571344 109006 571356
rect 140774 571344 140780 571356
rect 140832 571344 140838 571396
rect 66162 571276 66168 571328
rect 66220 571316 66226 571328
rect 68278 571316 68284 571328
rect 66220 571288 68284 571316
rect 66220 571276 66226 571288
rect 68278 571276 68284 571288
rect 68336 571276 68342 571328
rect 63218 569916 63224 569968
rect 63276 569956 63282 569968
rect 67634 569956 67640 569968
rect 63276 569928 67640 569956
rect 63276 569916 63282 569928
rect 67634 569916 67640 569928
rect 67692 569916 67698 569968
rect 108942 569916 108948 569968
rect 109000 569956 109006 569968
rect 142154 569956 142160 569968
rect 109000 569928 142160 569956
rect 109000 569916 109006 569928
rect 142154 569916 142160 569928
rect 142212 569916 142218 569968
rect 107654 568624 107660 568676
rect 107712 568664 107718 568676
rect 109770 568664 109776 568676
rect 107712 568636 109776 568664
rect 107712 568624 107718 568636
rect 109770 568624 109776 568636
rect 109828 568624 109834 568676
rect 66162 568556 66168 568608
rect 66220 568596 66226 568608
rect 67634 568596 67640 568608
rect 66220 568568 67640 568596
rect 66220 568556 66226 568568
rect 67634 568556 67640 568568
rect 67692 568556 67698 568608
rect 108942 567536 108948 567588
rect 109000 567576 109006 567588
rect 114738 567576 114744 567588
rect 109000 567548 114744 567576
rect 109000 567536 109006 567548
rect 114738 567536 114744 567548
rect 114796 567536 114802 567588
rect 64690 567264 64696 567316
rect 64748 567304 64754 567316
rect 67634 567304 67640 567316
rect 64748 567276 67640 567304
rect 64748 567264 64754 567276
rect 67634 567264 67640 567276
rect 67692 567264 67698 567316
rect 63310 567196 63316 567248
rect 63368 567236 63374 567248
rect 67726 567236 67732 567248
rect 63368 567208 67732 567236
rect 63368 567196 63374 567208
rect 67726 567196 67732 567208
rect 67784 567196 67790 567248
rect 108942 567196 108948 567248
rect 109000 567236 109006 567248
rect 117958 567236 117964 567248
rect 109000 567208 117964 567236
rect 109000 567196 109006 567208
rect 117958 567196 117964 567208
rect 118016 567196 118022 567248
rect 108850 565904 108856 565956
rect 108908 565944 108914 565956
rect 125778 565944 125784 565956
rect 108908 565916 125784 565944
rect 108908 565904 108914 565916
rect 125778 565904 125784 565916
rect 125836 565904 125842 565956
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 25498 565876 25504 565888
rect 3292 565848 25504 565876
rect 3292 565836 3298 565848
rect 25498 565836 25504 565848
rect 25556 565836 25562 565888
rect 63126 565836 63132 565888
rect 63184 565876 63190 565888
rect 67634 565876 67640 565888
rect 63184 565848 67640 565876
rect 63184 565836 63190 565848
rect 67634 565836 67640 565848
rect 67692 565836 67698 565888
rect 108942 565836 108948 565888
rect 109000 565876 109006 565888
rect 142246 565876 142252 565888
rect 109000 565848 142252 565876
rect 109000 565836 109006 565848
rect 142246 565836 142252 565848
rect 142304 565836 142310 565888
rect 431218 565088 431224 565140
rect 431276 565128 431282 565140
rect 497458 565128 497464 565140
rect 431276 565100 497464 565128
rect 431276 565088 431282 565100
rect 497458 565088 497464 565100
rect 497516 565128 497522 565140
rect 504358 565128 504364 565140
rect 497516 565100 504364 565128
rect 497516 565088 497522 565100
rect 504358 565088 504364 565100
rect 504416 565088 504422 565140
rect 57698 564408 57704 564460
rect 57756 564448 57762 564460
rect 67634 564448 67640 564460
rect 57756 564420 67640 564448
rect 57756 564408 57762 564420
rect 67634 564408 67640 564420
rect 67692 564408 67698 564460
rect 108850 564408 108856 564460
rect 108908 564448 108914 564460
rect 133874 564448 133880 564460
rect 108908 564420 133880 564448
rect 108908 564408 108914 564420
rect 133874 564408 133880 564420
rect 133932 564448 133938 564460
rect 204898 564448 204904 564460
rect 133932 564420 204904 564448
rect 133932 564408 133938 564420
rect 204898 564408 204904 564420
rect 204956 564408 204962 564460
rect 108942 564340 108948 564392
rect 109000 564380 109006 564392
rect 117222 564380 117228 564392
rect 109000 564352 117228 564380
rect 109000 564340 109006 564352
rect 117222 564340 117228 564352
rect 117280 564380 117286 564392
rect 124306 564380 124312 564392
rect 117280 564352 124312 564380
rect 117280 564340 117286 564352
rect 124306 564340 124312 564352
rect 124364 564340 124370 564392
rect 504358 563660 504364 563712
rect 504416 563700 504422 563712
rect 580166 563700 580172 563712
rect 504416 563672 580172 563700
rect 504416 563660 504422 563672
rect 580166 563660 580172 563672
rect 580224 563660 580230 563712
rect 60458 563116 60464 563168
rect 60516 563156 60522 563168
rect 67634 563156 67640 563168
rect 60516 563128 67640 563156
rect 60516 563116 60522 563128
rect 67634 563116 67640 563128
rect 67692 563116 67698 563168
rect 52270 563048 52276 563100
rect 52328 563088 52334 563100
rect 67726 563088 67732 563100
rect 52328 563060 67732 563088
rect 52328 563048 52334 563060
rect 67726 563048 67732 563060
rect 67784 563048 67790 563100
rect 60734 562300 60740 562352
rect 60792 562340 60798 562352
rect 62022 562340 62028 562352
rect 60792 562312 62028 562340
rect 60792 562300 60798 562312
rect 62022 562300 62028 562312
rect 62080 562340 62086 562352
rect 67634 562340 67640 562352
rect 62080 562312 67640 562340
rect 62080 562300 62086 562312
rect 67634 562300 67640 562312
rect 67692 562300 67698 562352
rect 61838 561688 61844 561740
rect 61896 561728 61902 561740
rect 67634 561728 67640 561740
rect 61896 561700 67640 561728
rect 61896 561688 61902 561700
rect 67634 561688 67640 561700
rect 67692 561688 67698 561740
rect 108942 561688 108948 561740
rect 109000 561728 109006 561740
rect 130010 561728 130016 561740
rect 109000 561700 130016 561728
rect 109000 561688 109006 561700
rect 130010 561688 130016 561700
rect 130068 561688 130074 561740
rect 52178 560940 52184 560992
rect 52236 560980 52242 560992
rect 60734 560980 60740 560992
rect 52236 560952 60740 560980
rect 52236 560940 52242 560952
rect 60734 560940 60740 560952
rect 60792 560940 60798 560992
rect 106918 560940 106924 560992
rect 106976 560980 106982 560992
rect 116118 560980 116124 560992
rect 106976 560952 116124 560980
rect 106976 560940 106982 560952
rect 116118 560940 116124 560952
rect 116176 560940 116182 560992
rect 59262 560328 59268 560380
rect 59320 560368 59326 560380
rect 67726 560368 67732 560380
rect 59320 560340 67732 560368
rect 59320 560328 59326 560340
rect 67726 560328 67732 560340
rect 67784 560328 67790 560380
rect 107654 560328 107660 560380
rect 107712 560368 107718 560380
rect 138106 560368 138112 560380
rect 107712 560340 138112 560368
rect 107712 560328 107718 560340
rect 138106 560328 138112 560340
rect 138164 560328 138170 560380
rect 50982 560260 50988 560312
rect 51040 560300 51046 560312
rect 67634 560300 67640 560312
rect 51040 560272 67640 560300
rect 51040 560260 51046 560272
rect 67634 560260 67640 560272
rect 67692 560260 67698 560312
rect 108942 560260 108948 560312
rect 109000 560300 109006 560312
rect 139486 560300 139492 560312
rect 109000 560272 139492 560300
rect 109000 560260 109006 560272
rect 139486 560260 139492 560272
rect 139544 560260 139550 560312
rect 136818 559512 136824 559564
rect 136876 559552 136882 559564
rect 201494 559552 201500 559564
rect 136876 559524 201500 559552
rect 136876 559512 136882 559524
rect 201494 559512 201500 559524
rect 201552 559512 201558 559564
rect 108942 558968 108948 559020
rect 109000 559008 109006 559020
rect 124214 559008 124220 559020
rect 109000 558980 124220 559008
rect 109000 558968 109006 558980
rect 124214 558968 124220 558980
rect 124272 558968 124278 559020
rect 42702 558900 42708 558952
rect 42760 558940 42766 558952
rect 67634 558940 67640 558952
rect 42760 558912 67640 558940
rect 42760 558900 42766 558912
rect 67634 558900 67640 558912
rect 67692 558900 67698 558952
rect 108850 558900 108856 558952
rect 108908 558940 108914 558952
rect 136818 558940 136824 558952
rect 108908 558912 136824 558940
rect 108908 558900 108914 558912
rect 136818 558900 136824 558912
rect 136876 558900 136882 558952
rect 37090 558152 37096 558204
rect 37148 558192 37154 558204
rect 68830 558192 68836 558204
rect 37148 558164 68836 558192
rect 37148 558152 37154 558164
rect 68830 558152 68836 558164
rect 68888 558152 68894 558204
rect 108942 557744 108948 557796
rect 109000 557784 109006 557796
rect 114646 557784 114652 557796
rect 109000 557756 114652 557784
rect 109000 557744 109006 557756
rect 114646 557744 114652 557756
rect 114704 557744 114710 557796
rect 30282 557540 30288 557592
rect 30340 557580 30346 557592
rect 67634 557580 67640 557592
rect 30340 557552 67640 557580
rect 30340 557540 30346 557552
rect 67634 557540 67640 557552
rect 67692 557540 67698 557592
rect 48130 556248 48136 556300
rect 48188 556288 48194 556300
rect 67634 556288 67640 556300
rect 48188 556260 67640 556288
rect 48188 556248 48194 556260
rect 67634 556248 67640 556260
rect 67692 556248 67698 556300
rect 43898 556180 43904 556232
rect 43956 556220 43962 556232
rect 67726 556220 67732 556232
rect 43956 556192 67732 556220
rect 43956 556180 43962 556192
rect 67726 556180 67732 556192
rect 67784 556180 67790 556232
rect 108942 556180 108948 556232
rect 109000 556220 109006 556232
rect 127618 556220 127624 556232
rect 109000 556192 127624 556220
rect 109000 556180 109006 556192
rect 127618 556180 127624 556192
rect 127676 556180 127682 556232
rect 108850 556112 108856 556164
rect 108908 556152 108914 556164
rect 110598 556152 110604 556164
rect 108908 556124 110604 556152
rect 108908 556112 108914 556124
rect 110598 556112 110604 556124
rect 110656 556112 110662 556164
rect 110598 555432 110604 555484
rect 110656 555472 110662 555484
rect 119430 555472 119436 555484
rect 110656 555444 119436 555472
rect 110656 555432 110662 555444
rect 119430 555432 119436 555444
rect 119488 555432 119494 555484
rect 57974 554820 57980 554872
rect 58032 554860 58038 554872
rect 67634 554860 67640 554872
rect 58032 554832 67640 554860
rect 58032 554820 58038 554832
rect 67634 554820 67640 554832
rect 67692 554820 67698 554872
rect 35710 554752 35716 554804
rect 35768 554792 35774 554804
rect 67726 554792 67732 554804
rect 35768 554764 67732 554792
rect 35768 554752 35774 554764
rect 67726 554752 67732 554764
rect 67784 554752 67790 554804
rect 3510 554684 3516 554736
rect 3568 554724 3574 554736
rect 14458 554724 14464 554736
rect 3568 554696 14464 554724
rect 3568 554684 3574 554696
rect 14458 554684 14464 554696
rect 14516 554684 14522 554736
rect 141510 554004 141516 554056
rect 141568 554044 141574 554056
rect 556798 554044 556804 554056
rect 141568 554016 556804 554044
rect 141568 554004 141574 554016
rect 556798 554004 556804 554016
rect 556856 554004 556862 554056
rect 65610 553392 65616 553444
rect 65668 553432 65674 553444
rect 67634 553432 67640 553444
rect 65668 553404 67640 553432
rect 65668 553392 65674 553404
rect 67634 553392 67640 553404
rect 67692 553392 67698 553444
rect 108942 553392 108948 553444
rect 109000 553432 109006 553444
rect 140958 553432 140964 553444
rect 109000 553404 140964 553432
rect 109000 553392 109006 553404
rect 140958 553392 140964 553404
rect 141016 553432 141022 553444
rect 141510 553432 141516 553444
rect 141016 553404 141516 553432
rect 141016 553392 141022 553404
rect 141510 553392 141516 553404
rect 141568 553392 141574 553444
rect 55030 552032 55036 552084
rect 55088 552072 55094 552084
rect 67634 552072 67640 552084
rect 55088 552044 67640 552072
rect 55088 552032 55094 552044
rect 67634 552032 67640 552044
rect 67692 552032 67698 552084
rect 108942 552032 108948 552084
rect 109000 552072 109006 552084
rect 138014 552072 138020 552084
rect 109000 552044 138020 552072
rect 109000 552032 109006 552044
rect 138014 552032 138020 552044
rect 138072 552032 138078 552084
rect 107654 550672 107660 550724
rect 107712 550712 107718 550724
rect 110690 550712 110696 550724
rect 107712 550684 110696 550712
rect 107712 550672 107718 550684
rect 110690 550672 110696 550684
rect 110748 550672 110754 550724
rect 46750 550604 46756 550656
rect 46808 550644 46814 550656
rect 67634 550644 67640 550656
rect 46808 550616 67640 550644
rect 46808 550604 46814 550616
rect 67634 550604 67640 550616
rect 67692 550604 67698 550656
rect 108942 550604 108948 550656
rect 109000 550644 109006 550656
rect 125594 550644 125600 550656
rect 109000 550616 125600 550644
rect 109000 550604 109006 550616
rect 125594 550604 125600 550616
rect 125652 550604 125658 550656
rect 108850 549312 108856 549364
rect 108908 549352 108914 549364
rect 135438 549352 135444 549364
rect 108908 549324 135444 549352
rect 108908 549312 108914 549324
rect 135438 549312 135444 549324
rect 135496 549312 135502 549364
rect 41138 549244 41144 549296
rect 41196 549284 41202 549296
rect 67634 549284 67640 549296
rect 41196 549256 67640 549284
rect 41196 549244 41202 549256
rect 67634 549244 67640 549256
rect 67692 549244 67698 549296
rect 108942 549244 108948 549296
rect 109000 549284 109006 549296
rect 139578 549284 139584 549296
rect 109000 549256 139584 549284
rect 109000 549244 109006 549256
rect 139578 549244 139584 549256
rect 139636 549244 139642 549296
rect 64782 547952 64788 548004
rect 64840 547992 64846 548004
rect 67634 547992 67640 548004
rect 64840 547964 67640 547992
rect 64840 547952 64846 547964
rect 67634 547952 67640 547964
rect 67692 547952 67698 548004
rect 56410 547884 56416 547936
rect 56468 547924 56474 547936
rect 67726 547924 67732 547936
rect 56468 547896 67732 547924
rect 56468 547884 56474 547896
rect 67726 547884 67732 547896
rect 67784 547884 67790 547936
rect 61654 546524 61660 546576
rect 61712 546564 61718 546576
rect 67726 546564 67732 546576
rect 61712 546536 67732 546564
rect 61712 546524 61718 546536
rect 67726 546524 67732 546536
rect 67784 546524 67790 546576
rect 60550 546456 60556 546508
rect 60608 546496 60614 546508
rect 67634 546496 67640 546508
rect 60608 546468 67640 546496
rect 60608 546456 60614 546468
rect 67634 546456 67640 546468
rect 67692 546456 67698 546508
rect 108942 546456 108948 546508
rect 109000 546496 109006 546508
rect 132586 546496 132592 546508
rect 109000 546468 132592 546496
rect 109000 546456 109006 546468
rect 132586 546456 132592 546468
rect 132644 546456 132650 546508
rect 108942 545708 108948 545760
rect 109000 545748 109006 545760
rect 112346 545748 112352 545760
rect 109000 545720 112352 545748
rect 109000 545708 109006 545720
rect 112346 545708 112352 545720
rect 112404 545708 112410 545760
rect 33042 545096 33048 545148
rect 33100 545136 33106 545148
rect 68094 545136 68100 545148
rect 33100 545108 68100 545136
rect 33100 545096 33106 545108
rect 68094 545096 68100 545108
rect 68152 545096 68158 545148
rect 108942 545096 108948 545148
rect 109000 545136 109006 545148
rect 134242 545136 134248 545148
rect 109000 545108 134248 545136
rect 109000 545096 109006 545108
rect 134242 545096 134248 545108
rect 134300 545096 134306 545148
rect 25498 544348 25504 544400
rect 25556 544388 25562 544400
rect 68002 544388 68008 544400
rect 25556 544360 68008 544388
rect 25556 544348 25562 544360
rect 68002 544348 68008 544360
rect 68060 544348 68066 544400
rect 108942 544348 108948 544400
rect 109000 544388 109006 544400
rect 115842 544388 115848 544400
rect 109000 544360 115848 544388
rect 109000 544348 109006 544360
rect 115842 544348 115848 544360
rect 115900 544388 115906 544400
rect 116210 544388 116216 544400
rect 115900 544360 116216 544388
rect 115900 544348 115906 544360
rect 116210 544348 116216 544360
rect 116268 544348 116274 544400
rect 108942 543736 108948 543788
rect 109000 543776 109006 543788
rect 140866 543776 140872 543788
rect 109000 543748 140872 543776
rect 109000 543736 109006 543748
rect 140866 543736 140872 543748
rect 140924 543736 140930 543788
rect 63402 542444 63408 542496
rect 63460 542484 63466 542496
rect 67634 542484 67640 542496
rect 63460 542456 67640 542484
rect 63460 542444 63466 542456
rect 67634 542444 67640 542456
rect 67692 542444 67698 542496
rect 45462 542376 45468 542428
rect 45520 542416 45526 542428
rect 68002 542416 68008 542428
rect 45520 542388 68008 542416
rect 45520 542376 45526 542388
rect 68002 542376 68008 542388
rect 68060 542376 68066 542428
rect 107838 542376 107844 542428
rect 107896 542416 107902 542428
rect 134150 542416 134156 542428
rect 107896 542388 134156 542416
rect 107896 542376 107902 542388
rect 134150 542376 134156 542388
rect 134208 542376 134214 542428
rect 61930 541628 61936 541680
rect 61988 541668 61994 541680
rect 69658 541668 69664 541680
rect 61988 541640 69664 541668
rect 61988 541628 61994 541640
rect 69658 541628 69664 541640
rect 69716 541628 69722 541680
rect 60642 540948 60648 541000
rect 60700 540988 60706 541000
rect 67634 540988 67640 541000
rect 60700 540960 67640 540988
rect 60700 540948 60706 540960
rect 67634 540948 67640 540960
rect 67692 540948 67698 541000
rect 108298 540744 108304 540796
rect 108356 540784 108362 540796
rect 109678 540784 109684 540796
rect 108356 540756 109684 540784
rect 108356 540744 108362 540756
rect 109678 540744 109684 540756
rect 109736 540744 109742 540796
rect 62022 539588 62028 539640
rect 62080 539628 62086 539640
rect 67634 539628 67640 539640
rect 62080 539600 67640 539628
rect 62080 539588 62086 539600
rect 67634 539588 67640 539600
rect 67692 539588 67698 539640
rect 106826 539588 106832 539640
rect 106884 539628 106890 539640
rect 142430 539628 142436 539640
rect 106884 539600 142436 539628
rect 106884 539588 106890 539600
rect 142430 539588 142436 539600
rect 142488 539588 142494 539640
rect 3418 539520 3424 539572
rect 3476 539560 3482 539572
rect 98362 539560 98368 539572
rect 3476 539532 98368 539560
rect 3476 539520 3482 539532
rect 98362 539520 98368 539532
rect 98420 539520 98426 539572
rect 425054 539520 425060 539572
rect 425112 539560 425118 539572
rect 425698 539560 425704 539572
rect 425112 539532 425704 539560
rect 425112 539520 425118 539532
rect 425698 539520 425704 539532
rect 425756 539520 425762 539572
rect 58618 539452 58624 539504
rect 58676 539492 58682 539504
rect 99006 539492 99012 539504
rect 58676 539464 99012 539492
rect 58676 539452 58682 539464
rect 99006 539452 99012 539464
rect 99064 539452 99070 539504
rect 70302 539044 70308 539096
rect 70360 539084 70366 539096
rect 71958 539084 71964 539096
rect 70360 539056 71964 539084
rect 70360 539044 70366 539056
rect 71958 539044 71964 539056
rect 72016 539044 72022 539096
rect 95142 538976 95148 539028
rect 95200 539016 95206 539028
rect 109126 539016 109132 539028
rect 95200 538988 109132 539016
rect 95200 538976 95206 538988
rect 109126 538976 109132 538988
rect 109184 538976 109190 539028
rect 99282 538908 99288 538960
rect 99340 538948 99346 538960
rect 121546 538948 121552 538960
rect 99340 538920 121552 538948
rect 99340 538908 99346 538920
rect 121546 538908 121552 538920
rect 121604 538908 121610 538960
rect 99006 538840 99012 538892
rect 99064 538880 99070 538892
rect 129918 538880 129924 538892
rect 99064 538852 129924 538880
rect 99064 538840 99070 538852
rect 129918 538840 129924 538852
rect 129976 538840 129982 538892
rect 41322 538228 41328 538280
rect 41380 538268 41386 538280
rect 59998 538268 60004 538280
rect 41380 538240 60004 538268
rect 41380 538228 41386 538240
rect 59998 538228 60004 538240
rect 60056 538268 60062 538280
rect 60056 538240 60688 538268
rect 60056 538228 60062 538240
rect 60660 538200 60688 538240
rect 109678 538228 109684 538280
rect 109736 538268 109742 538280
rect 123478 538268 123484 538280
rect 109736 538240 123484 538268
rect 109736 538228 109742 538240
rect 123478 538228 123484 538240
rect 123536 538268 123542 538280
rect 425054 538268 425060 538280
rect 123536 538240 425060 538268
rect 123536 538228 123542 538240
rect 425054 538228 425060 538240
rect 425112 538228 425118 538280
rect 73890 538200 73896 538212
rect 60660 538172 73896 538200
rect 73890 538160 73896 538172
rect 73948 538160 73954 538212
rect 80330 538160 80336 538212
rect 80388 538200 80394 538212
rect 111058 538200 111064 538212
rect 80388 538172 111064 538200
rect 80388 538160 80394 538172
rect 111058 538160 111064 538172
rect 111116 538160 111122 538212
rect 204898 538160 204904 538212
rect 204956 538200 204962 538212
rect 580166 538200 580172 538212
rect 204956 538172 580172 538200
rect 204956 538160 204962 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 100938 538092 100944 538144
rect 100996 538132 101002 538144
rect 119338 538132 119344 538144
rect 100996 538104 119344 538132
rect 100996 538092 101002 538104
rect 119338 538092 119344 538104
rect 119396 538092 119402 538144
rect 53742 537684 53748 537736
rect 53800 537724 53806 537736
rect 82906 537724 82912 537736
rect 53800 537696 82912 537724
rect 53800 537684 53806 537696
rect 82906 537684 82912 537696
rect 82964 537684 82970 537736
rect 97074 537684 97080 537736
rect 97132 537724 97138 537736
rect 102134 537724 102140 537736
rect 97132 537696 102140 537724
rect 97132 537684 97138 537696
rect 102134 537684 102140 537696
rect 102192 537684 102198 537736
rect 102226 537684 102232 537736
rect 102284 537724 102290 537736
rect 110598 537724 110604 537736
rect 102284 537696 110604 537724
rect 102284 537684 102290 537696
rect 110598 537684 110604 537696
rect 110656 537684 110662 537736
rect 46658 537616 46664 537668
rect 46716 537656 46722 537668
rect 79686 537656 79692 537668
rect 46716 537628 79692 537656
rect 46716 537616 46722 537628
rect 79686 537616 79692 537628
rect 79744 537616 79750 537668
rect 84102 537616 84108 537668
rect 84160 537656 84166 537668
rect 89990 537656 89996 537668
rect 84160 537628 89996 537656
rect 84160 537616 84166 537628
rect 89990 537616 89996 537628
rect 90048 537616 90054 537668
rect 102870 537616 102876 537668
rect 102928 537656 102934 537668
rect 128538 537656 128544 537668
rect 102928 537628 128544 537656
rect 102928 537616 102934 537628
rect 128538 537616 128544 537628
rect 128596 537616 128602 537668
rect 53190 537548 53196 537600
rect 53248 537588 53254 537600
rect 86126 537588 86132 537600
rect 53248 537560 86132 537588
rect 53248 537548 53254 537560
rect 86126 537548 86132 537560
rect 86184 537548 86190 537600
rect 95786 537548 95792 537600
rect 95844 537588 95850 537600
rect 121638 537588 121644 537600
rect 95844 537560 121644 537588
rect 95844 537548 95850 537560
rect 121638 537548 121644 537560
rect 121696 537548 121702 537600
rect 15838 537480 15844 537532
rect 15896 537520 15902 537532
rect 57514 537520 57520 537532
rect 15896 537492 57520 537520
rect 15896 537480 15902 537492
rect 57514 537480 57520 537492
rect 57572 537520 57578 537532
rect 91278 537520 91284 537532
rect 57572 537492 91284 537520
rect 57572 537480 57578 537492
rect 91278 537480 91284 537492
rect 91336 537480 91342 537532
rect 100294 537480 100300 537532
rect 100352 537520 100358 537532
rect 132678 537520 132684 537532
rect 100352 537492 132684 537520
rect 100352 537480 100358 537492
rect 132678 537480 132684 537492
rect 132736 537480 132742 537532
rect 83458 536800 83464 536852
rect 83516 536840 83522 536852
rect 85482 536840 85488 536852
rect 83516 536812 85488 536840
rect 83516 536800 83522 536812
rect 85482 536800 85488 536812
rect 85540 536800 85546 536852
rect 94498 536800 94504 536852
rect 94556 536840 94562 536852
rect 94556 536812 102088 536840
rect 94556 536800 94562 536812
rect 102060 536772 102088 536812
rect 117406 536772 117412 536784
rect 102060 536744 117412 536772
rect 117406 536732 117412 536744
rect 117464 536732 117470 536784
rect 101950 536664 101956 536716
rect 102008 536704 102014 536716
rect 105538 536704 105544 536716
rect 102008 536676 105544 536704
rect 102008 536664 102014 536676
rect 105538 536664 105544 536676
rect 105596 536664 105602 536716
rect 38470 536052 38476 536104
rect 38528 536092 38534 536104
rect 71314 536092 71320 536104
rect 38528 536064 71320 536092
rect 38528 536052 38534 536064
rect 71314 536052 71320 536064
rect 71372 536052 71378 536104
rect 117406 535440 117412 535492
rect 117464 535480 117470 535492
rect 118694 535480 118700 535492
rect 117464 535452 118700 535480
rect 117464 535440 117470 535452
rect 118694 535440 118700 535452
rect 118752 535440 118758 535492
rect 57790 534964 57796 535016
rect 57848 535004 57854 535016
rect 75178 535004 75184 535016
rect 57848 534976 75184 535004
rect 57848 534964 57854 534976
rect 75178 534964 75184 534976
rect 75236 534964 75242 535016
rect 51994 534896 52000 534948
rect 52052 534936 52058 534948
rect 78398 534936 78404 534948
rect 52052 534908 78404 534936
rect 52052 534896 52058 534908
rect 78398 534896 78404 534908
rect 78456 534896 78462 534948
rect 50890 534828 50896 534880
rect 50948 534868 50954 534880
rect 83550 534868 83556 534880
rect 50948 534840 83556 534868
rect 50948 534828 50954 534840
rect 83550 534828 83556 534840
rect 83608 534828 83614 534880
rect 45278 534760 45284 534812
rect 45336 534800 45342 534812
rect 77754 534800 77760 534812
rect 45336 534772 77760 534800
rect 45336 534760 45342 534772
rect 77754 534760 77760 534772
rect 77812 534760 77818 534812
rect 91002 534760 91008 534812
rect 91060 534800 91066 534812
rect 115934 534800 115940 534812
rect 91060 534772 115940 534800
rect 91060 534760 91066 534772
rect 115934 534760 115940 534772
rect 115992 534760 115998 534812
rect 39942 534692 39948 534744
rect 40000 534732 40006 534744
rect 73246 534732 73252 534744
rect 40000 534704 73252 534732
rect 40000 534692 40006 534704
rect 73246 534692 73252 534704
rect 73304 534692 73310 534744
rect 93854 534692 93860 534744
rect 93912 534732 93918 534744
rect 128354 534732 128360 534744
rect 93912 534704 128360 534732
rect 93912 534692 93918 534704
rect 128354 534692 128360 534704
rect 128412 534692 128418 534744
rect 420914 534692 420920 534744
rect 420972 534732 420978 534744
rect 429194 534732 429200 534744
rect 420972 534704 429200 534732
rect 420972 534692 420978 534704
rect 429194 534692 429200 534704
rect 429252 534692 429258 534744
rect 52362 533332 52368 533384
rect 52420 533372 52426 533384
rect 52420 533344 64874 533372
rect 52420 533332 52426 533344
rect 64846 533304 64874 533344
rect 69290 533332 69296 533384
rect 69348 533372 69354 533384
rect 69750 533372 69756 533384
rect 69348 533344 69756 533372
rect 69348 533332 69354 533344
rect 69750 533332 69756 533344
rect 69808 533332 69814 533384
rect 72418 533304 72424 533316
rect 64846 533276 72424 533304
rect 72418 533264 72424 533276
rect 72476 533264 72482 533316
rect 52086 532176 52092 532228
rect 52144 532216 52150 532228
rect 72602 532216 72608 532228
rect 52144 532188 72608 532216
rect 52144 532176 52150 532188
rect 72602 532176 72608 532188
rect 72660 532176 72666 532228
rect 55122 532108 55128 532160
rect 55180 532148 55186 532160
rect 76466 532148 76472 532160
rect 55180 532120 76472 532148
rect 55180 532108 55186 532120
rect 76466 532108 76472 532120
rect 76524 532108 76530 532160
rect 45370 532040 45376 532092
rect 45428 532080 45434 532092
rect 75086 532080 75092 532092
rect 45428 532052 75092 532080
rect 45428 532040 45434 532052
rect 75086 532040 75092 532052
rect 75144 532040 75150 532092
rect 84838 532040 84844 532092
rect 84896 532080 84902 532092
rect 111978 532080 111984 532092
rect 84896 532052 111984 532080
rect 84896 532040 84902 532052
rect 111978 532040 111984 532052
rect 112036 532040 112042 532092
rect 39666 531972 39672 532024
rect 39724 532012 39730 532024
rect 71866 532012 71872 532024
rect 39724 531984 71872 532012
rect 39724 531972 39730 531984
rect 71866 531972 71872 531984
rect 71924 531972 71930 532024
rect 93762 531972 93768 532024
rect 93820 532012 93826 532024
rect 123018 532012 123024 532024
rect 93820 531984 123024 532012
rect 93820 531972 93826 531984
rect 123018 531972 123024 531984
rect 123076 531972 123082 532024
rect 41046 529252 41052 529304
rect 41104 529292 41110 529304
rect 70394 529292 70400 529304
rect 41104 529264 70400 529292
rect 41104 529252 41110 529264
rect 70394 529252 70400 529264
rect 70452 529252 70458 529304
rect 42518 529184 42524 529236
rect 42576 529224 42582 529236
rect 77110 529224 77116 529236
rect 42576 529196 77116 529224
rect 42576 529184 42582 529196
rect 77110 529184 77116 529196
rect 77168 529184 77174 529236
rect 110690 529184 110696 529236
rect 110748 529224 110754 529236
rect 116670 529224 116676 529236
rect 110748 529196 116676 529224
rect 110748 529184 110754 529196
rect 116670 529184 116676 529196
rect 116728 529184 116734 529236
rect 110690 528612 110696 528624
rect 106246 528584 110696 528612
rect 3142 528504 3148 528556
rect 3200 528544 3206 528556
rect 106246 528544 106274 528584
rect 110690 528572 110696 528584
rect 110748 528572 110754 528624
rect 3200 528516 106274 528544
rect 3200 528504 3206 528516
rect 69198 525716 69204 525768
rect 69256 525756 69262 525768
rect 579798 525756 579804 525768
rect 69256 525728 579804 525756
rect 69256 525716 69262 525728
rect 579798 525716 579804 525728
rect 579856 525716 579862 525768
rect 2774 514768 2780 514820
rect 2832 514808 2838 514820
rect 4798 514808 4804 514820
rect 2832 514780 4804 514808
rect 2832 514768 2838 514780
rect 4798 514768 4804 514780
rect 4856 514768 4862 514820
rect 431218 510620 431224 510672
rect 431276 510660 431282 510672
rect 580166 510660 580172 510672
rect 431276 510632 580172 510660
rect 431276 510620 431282 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 114830 499576 114836 499588
rect 93872 499548 114836 499576
rect 87414 499468 87420 499520
rect 87472 499508 87478 499520
rect 93872 499508 93900 499548
rect 114830 499536 114836 499548
rect 114888 499576 114894 499588
rect 131206 499576 131212 499588
rect 114888 499548 131212 499576
rect 114888 499536 114894 499548
rect 131206 499536 131212 499548
rect 131264 499536 131270 499588
rect 87472 499480 93900 499508
rect 87472 499468 87478 499480
rect 89346 498856 89352 498908
rect 89404 498896 89410 498908
rect 113542 498896 113548 498908
rect 89404 498868 113548 498896
rect 89404 498856 89410 498868
rect 113542 498856 113548 498868
rect 113600 498856 113606 498908
rect 69658 498788 69664 498840
rect 69716 498828 69722 498840
rect 74534 498828 74540 498840
rect 69716 498800 74540 498828
rect 69716 498788 69722 498800
rect 74534 498788 74540 498800
rect 74592 498828 74598 498840
rect 80606 498828 80612 498840
rect 74592 498800 80612 498828
rect 74592 498788 74598 498800
rect 80606 498788 80612 498800
rect 80664 498788 80670 498840
rect 88058 498788 88064 498840
rect 88116 498828 88122 498840
rect 128446 498828 128452 498840
rect 88116 498800 128452 498828
rect 88116 498788 88122 498800
rect 128446 498788 128452 498800
rect 128504 498788 128510 498840
rect 4798 498108 4804 498160
rect 4856 498148 4862 498160
rect 59170 498148 59176 498160
rect 4856 498120 59176 498148
rect 4856 498108 4862 498120
rect 59170 498108 59176 498120
rect 59228 498108 59234 498160
rect 59170 497632 59176 497684
rect 59228 497672 59234 497684
rect 91094 497672 91100 497684
rect 59228 497644 91100 497672
rect 59228 497632 59234 497644
rect 91094 497632 91100 497644
rect 91152 497632 91158 497684
rect 93210 497632 93216 497684
rect 93268 497672 93274 497684
rect 117498 497672 117504 497684
rect 93268 497644 117504 497672
rect 93268 497632 93274 497644
rect 117498 497632 117504 497644
rect 117556 497632 117562 497684
rect 85574 497564 85580 497616
rect 85632 497604 85638 497616
rect 120166 497604 120172 497616
rect 85632 497576 120172 497604
rect 85632 497564 85638 497576
rect 120166 497564 120172 497576
rect 120224 497604 120230 497616
rect 126974 497604 126980 497616
rect 120224 497576 126980 497604
rect 120224 497564 120230 497576
rect 126974 497564 126980 497576
rect 127032 497564 127038 497616
rect 84102 497496 84108 497548
rect 84160 497536 84166 497548
rect 120258 497536 120264 497548
rect 84160 497508 120264 497536
rect 84160 497496 84166 497508
rect 120258 497496 120264 497508
rect 120316 497496 120322 497548
rect 83274 497428 83280 497480
rect 83332 497468 83338 497480
rect 122926 497468 122932 497480
rect 83332 497440 122932 497468
rect 83332 497428 83338 497440
rect 122926 497428 122932 497440
rect 122984 497468 122990 497480
rect 131390 497468 131396 497480
rect 122984 497440 131396 497468
rect 122984 497428 122990 497440
rect 131390 497428 131396 497440
rect 131448 497428 131454 497480
rect 59280 496828 67588 496856
rect 53650 496748 53656 496800
rect 53708 496788 53714 496800
rect 58066 496788 58072 496800
rect 53708 496760 58072 496788
rect 53708 496748 53714 496760
rect 58066 496748 58072 496760
rect 58124 496788 58130 496800
rect 59280 496788 59308 496828
rect 58124 496760 59308 496788
rect 67560 496788 67588 496828
rect 430574 496788 430580 496800
rect 67560 496760 430580 496788
rect 58124 496748 58130 496760
rect 430574 496748 430580 496760
rect 430632 496748 430638 496800
rect 53650 496272 53656 496324
rect 53708 496312 53714 496324
rect 83458 496312 83464 496324
rect 53708 496284 83464 496312
rect 53708 496272 53714 496284
rect 83458 496272 83464 496284
rect 83516 496272 83522 496324
rect 81526 496204 81532 496256
rect 81584 496244 81590 496256
rect 116118 496244 116124 496256
rect 81584 496216 116124 496244
rect 81584 496204 81590 496216
rect 116118 496204 116124 496216
rect 116176 496204 116182 496256
rect 430574 496204 430580 496256
rect 430632 496244 430638 496256
rect 431218 496244 431224 496256
rect 430632 496216 431224 496244
rect 430632 496204 430638 496216
rect 431218 496204 431224 496216
rect 431276 496204 431282 496256
rect 79686 496136 79692 496188
rect 79744 496176 79750 496188
rect 113266 496176 113272 496188
rect 79744 496148 113272 496176
rect 79744 496136 79750 496148
rect 113266 496136 113272 496148
rect 113324 496176 113330 496188
rect 116578 496176 116584 496188
rect 113324 496148 116584 496176
rect 113324 496136 113330 496148
rect 116578 496136 116584 496148
rect 116636 496136 116642 496188
rect 49418 496068 49424 496120
rect 49476 496108 49482 496120
rect 80974 496108 80980 496120
rect 49476 496080 80980 496108
rect 49476 496068 49482 496080
rect 80974 496068 80980 496080
rect 81032 496068 81038 496120
rect 95050 496068 95056 496120
rect 95108 496108 95114 496120
rect 131114 496108 131120 496120
rect 95108 496080 131120 496108
rect 95108 496068 95114 496080
rect 131114 496068 131120 496080
rect 131172 496108 131178 496120
rect 141050 496108 141056 496120
rect 131172 496080 141056 496108
rect 131172 496068 131178 496080
rect 141050 496068 141056 496080
rect 141108 496068 141114 496120
rect 78398 495456 78404 495508
rect 78456 495496 78462 495508
rect 112070 495496 112076 495508
rect 78456 495468 112076 495496
rect 78456 495456 78462 495468
rect 112070 495456 112076 495468
rect 112128 495456 112134 495508
rect 116118 495456 116124 495508
rect 116176 495496 116182 495508
rect 121546 495496 121552 495508
rect 116176 495468 121552 495496
rect 116176 495456 116182 495468
rect 121546 495456 121552 495468
rect 121604 495456 121610 495508
rect 3418 495388 3424 495440
rect 3476 495428 3482 495440
rect 83274 495428 83280 495440
rect 3476 495400 83280 495428
rect 3476 495388 3482 495400
rect 83274 495388 83280 495400
rect 83332 495388 83338 495440
rect 75178 494980 75184 495032
rect 75236 495020 75242 495032
rect 78398 495020 78404 495032
rect 75236 494992 78404 495020
rect 75236 494980 75242 494992
rect 78398 494980 78404 494992
rect 78456 494980 78462 495032
rect 94958 494980 94964 495032
rect 95016 495020 95022 495032
rect 111886 495020 111892 495032
rect 95016 494992 111892 495020
rect 95016 494980 95022 494992
rect 111886 494980 111892 494992
rect 111944 495020 111950 495032
rect 114830 495020 114836 495032
rect 111944 494992 114836 495020
rect 111944 494980 111950 494992
rect 114830 494980 114836 494992
rect 114888 494980 114894 495032
rect 98638 494912 98644 494964
rect 98696 494952 98702 494964
rect 120350 494952 120356 494964
rect 98696 494924 120356 494952
rect 98696 494912 98702 494924
rect 120350 494912 120356 494924
rect 120408 494912 120414 494964
rect 94866 494844 94872 494896
rect 94924 494884 94930 494896
rect 116026 494884 116032 494896
rect 94924 494856 116032 494884
rect 94924 494844 94930 494856
rect 116026 494844 116032 494856
rect 116084 494884 116090 494896
rect 132494 494884 132500 494896
rect 116084 494856 132500 494884
rect 116084 494844 116090 494856
rect 132494 494844 132500 494856
rect 132552 494844 132558 494896
rect 80974 494776 80980 494828
rect 81032 494816 81038 494828
rect 118786 494816 118792 494828
rect 81032 494788 118792 494816
rect 81032 494776 81038 494788
rect 118786 494776 118792 494788
rect 118844 494816 118850 494828
rect 125870 494816 125876 494828
rect 118844 494788 125876 494816
rect 118844 494776 118850 494788
rect 125870 494776 125876 494788
rect 125928 494776 125934 494828
rect 82906 494708 82912 494760
rect 82964 494748 82970 494760
rect 122834 494748 122840 494760
rect 82964 494720 122840 494748
rect 82964 494708 82970 494720
rect 122834 494708 122840 494720
rect 122892 494748 122898 494760
rect 130102 494748 130108 494760
rect 122892 494720 130108 494748
rect 122892 494708 122898 494720
rect 130102 494708 130108 494720
rect 130160 494708 130166 494760
rect 92474 494028 92480 494080
rect 92532 494068 92538 494080
rect 93762 494068 93768 494080
rect 92532 494040 93768 494068
rect 92532 494028 92538 494040
rect 93762 494028 93768 494040
rect 93820 494068 93826 494080
rect 110690 494068 110696 494080
rect 93820 494040 110696 494068
rect 93820 494028 93826 494040
rect 110690 494028 110696 494040
rect 110748 494028 110754 494080
rect 91922 493824 91928 493876
rect 91980 493864 91986 493876
rect 95050 493864 95056 493876
rect 91980 493836 95056 493864
rect 91980 493824 91986 493836
rect 95050 493824 95056 493836
rect 95108 493824 95114 493876
rect 95786 493484 95792 493536
rect 95844 493524 95850 493536
rect 95844 493496 113174 493524
rect 95844 493484 95850 493496
rect 90266 493416 90272 493468
rect 90324 493456 90330 493468
rect 110414 493456 110420 493468
rect 90324 493428 110420 493456
rect 90324 493416 90330 493428
rect 110414 493416 110420 493428
rect 110472 493416 110478 493468
rect 113146 493456 113174 493496
rect 113358 493456 113364 493468
rect 113146 493428 113364 493456
rect 113358 493416 113364 493428
rect 113416 493456 113422 493468
rect 127158 493456 127164 493468
rect 113416 493428 127164 493456
rect 113416 493416 113422 493428
rect 127158 493416 127164 493428
rect 127216 493416 127222 493468
rect 54110 493348 54116 493400
rect 54168 493388 54174 493400
rect 54938 493388 54944 493400
rect 54168 493360 54944 493388
rect 54168 493348 54174 493360
rect 54938 493348 54944 493360
rect 54996 493388 55002 493400
rect 74810 493388 74816 493400
rect 54996 493360 74816 493388
rect 54996 493348 55002 493360
rect 74810 493348 74816 493360
rect 74868 493348 74874 493400
rect 88702 493348 88708 493400
rect 88760 493388 88766 493400
rect 120074 493388 120080 493400
rect 88760 493360 120080 493388
rect 88760 493348 88766 493360
rect 120074 493348 120080 493360
rect 120132 493388 120138 493400
rect 122834 493388 122840 493400
rect 120132 493360 122840 493388
rect 120132 493348 120138 493360
rect 122834 493348 122840 493360
rect 122892 493348 122898 493400
rect 43990 493280 43996 493332
rect 44048 493320 44054 493332
rect 49510 493320 49516 493332
rect 44048 493292 49516 493320
rect 44048 493280 44054 493292
rect 49510 493280 49516 493292
rect 49568 493320 49574 493332
rect 71682 493320 71688 493332
rect 49568 493292 71688 493320
rect 49568 493280 49574 493292
rect 71682 493280 71688 493292
rect 71740 493280 71746 493332
rect 93210 493280 93216 493332
rect 93268 493320 93274 493332
rect 129826 493320 129832 493332
rect 93268 493292 129832 493320
rect 93268 493280 93274 493292
rect 129826 493280 129832 493292
rect 129884 493320 129890 493332
rect 139394 493320 139400 493332
rect 129884 493292 139400 493320
rect 129884 493280 129890 493292
rect 139394 493280 139400 493292
rect 139452 493280 139458 493332
rect 75822 493008 75828 493060
rect 75880 493048 75886 493060
rect 81526 493048 81532 493060
rect 75880 493020 81532 493048
rect 75880 493008 75886 493020
rect 81526 493008 81532 493020
rect 81584 493008 81590 493060
rect 81618 492804 81624 492856
rect 81676 492844 81682 492856
rect 96522 492844 96528 492856
rect 81676 492816 96528 492844
rect 81676 492804 81682 492816
rect 96522 492804 96528 492816
rect 96580 492804 96586 492856
rect 46566 492736 46572 492788
rect 46624 492776 46630 492788
rect 53834 492776 53840 492788
rect 46624 492748 53840 492776
rect 46624 492736 46630 492748
rect 53834 492736 53840 492748
rect 53892 492736 53898 492788
rect 57882 492736 57888 492788
rect 57940 492776 57946 492788
rect 90266 492776 90272 492788
rect 57940 492748 90272 492776
rect 57940 492736 57946 492748
rect 90266 492736 90272 492748
rect 90324 492736 90330 492788
rect 39850 492668 39856 492720
rect 39908 492708 39914 492720
rect 70946 492708 70952 492720
rect 39908 492680 70952 492708
rect 39908 492668 39914 492680
rect 70946 492668 70952 492680
rect 71004 492668 71010 492720
rect 77754 492668 77760 492720
rect 77812 492708 77818 492720
rect 120074 492708 120080 492720
rect 77812 492680 120080 492708
rect 77812 492668 77818 492680
rect 120074 492668 120080 492680
rect 120132 492668 120138 492720
rect 72418 492600 72424 492652
rect 72476 492640 72482 492652
rect 77772 492640 77800 492668
rect 72476 492612 77800 492640
rect 72476 492600 72482 492612
rect 84838 492600 84844 492652
rect 84896 492640 84902 492652
rect 92474 492640 92480 492652
rect 84896 492612 92480 492640
rect 84896 492600 84902 492612
rect 92474 492600 92480 492612
rect 92532 492600 92538 492652
rect 97718 492600 97724 492652
rect 97776 492640 97782 492652
rect 99282 492640 99288 492652
rect 97776 492612 99288 492640
rect 97776 492600 97782 492612
rect 99282 492600 99288 492612
rect 99340 492600 99346 492652
rect 53834 492124 53840 492176
rect 53892 492164 53898 492176
rect 54478 492164 54484 492176
rect 53892 492136 54484 492164
rect 53892 492124 53898 492136
rect 54478 492124 54484 492136
rect 54536 492164 54542 492176
rect 70394 492164 70400 492176
rect 54536 492136 70400 492164
rect 54536 492124 54542 492136
rect 70394 492124 70400 492136
rect 70452 492124 70458 492176
rect 50706 492056 50712 492108
rect 50764 492096 50770 492108
rect 70026 492096 70032 492108
rect 50764 492068 70032 492096
rect 50764 492056 50770 492068
rect 70026 492056 70032 492068
rect 70084 492056 70090 492108
rect 86126 492056 86132 492108
rect 86184 492096 86190 492108
rect 87138 492096 87144 492108
rect 86184 492068 87144 492096
rect 86184 492056 86190 492068
rect 87138 492056 87144 492068
rect 87196 492096 87202 492108
rect 89898 492096 89904 492108
rect 87196 492068 89904 492096
rect 87196 492056 87202 492068
rect 89898 492056 89904 492068
rect 89956 492056 89962 492108
rect 92014 492056 92020 492108
rect 92072 492096 92078 492108
rect 102410 492096 102416 492108
rect 92072 492068 102416 492096
rect 92072 492056 92078 492068
rect 102410 492056 102416 492068
rect 102468 492056 102474 492108
rect 114462 492056 114468 492108
rect 114520 492096 114526 492108
rect 125686 492096 125692 492108
rect 114520 492068 125692 492096
rect 114520 492056 114526 492068
rect 125686 492056 125692 492068
rect 125744 492056 125750 492108
rect 39758 491988 39764 492040
rect 39816 492028 39822 492040
rect 48038 492028 48044 492040
rect 39816 492000 48044 492028
rect 39816 491988 39822 492000
rect 48038 491988 48044 492000
rect 48096 492028 48102 492040
rect 72234 492028 72240 492040
rect 48096 492000 72240 492028
rect 48096 491988 48102 492000
rect 72234 491988 72240 492000
rect 72292 491988 72298 492040
rect 76466 491988 76472 492040
rect 76524 492028 76530 492040
rect 110506 492028 110512 492040
rect 76524 492000 110512 492028
rect 76524 491988 76530 492000
rect 110506 491988 110512 492000
rect 110564 492028 110570 492040
rect 123018 492028 123024 492040
rect 110564 492000 123024 492028
rect 110564 491988 110570 492000
rect 123018 491988 123024 492000
rect 123076 491988 123082 492040
rect 56134 491920 56140 491972
rect 56192 491960 56198 491972
rect 90634 491960 90640 491972
rect 56192 491932 90640 491960
rect 56192 491920 56198 491932
rect 90634 491920 90640 491932
rect 90692 491920 90698 491972
rect 97074 491920 97080 491972
rect 97132 491960 97138 491972
rect 131298 491960 131304 491972
rect 97132 491932 131304 491960
rect 97132 491920 97138 491932
rect 131298 491920 131304 491932
rect 131356 491960 131362 491972
rect 143534 491960 143540 491972
rect 131356 491932 143540 491960
rect 131356 491920 131362 491932
rect 143534 491920 143540 491932
rect 143592 491920 143598 491972
rect 89990 491784 89996 491836
rect 90048 491824 90054 491836
rect 91002 491824 91008 491836
rect 90048 491796 91008 491824
rect 90048 491784 90054 491796
rect 91002 491784 91008 491796
rect 91060 491784 91066 491836
rect 92566 491648 92572 491700
rect 92624 491688 92630 491700
rect 94958 491688 94964 491700
rect 92624 491660 94964 491688
rect 92624 491648 92630 491660
rect 94958 491648 94964 491660
rect 95016 491648 95022 491700
rect 95142 491648 95148 491700
rect 95200 491688 95206 491700
rect 96338 491688 96344 491700
rect 95200 491660 96344 491688
rect 95200 491648 95206 491660
rect 96338 491648 96344 491660
rect 96396 491648 96402 491700
rect 91002 491512 91008 491564
rect 91060 491552 91066 491564
rect 99926 491552 99932 491564
rect 91060 491524 99932 491552
rect 91060 491512 91066 491524
rect 99926 491512 99932 491524
rect 99984 491512 99990 491564
rect 71774 491444 71780 491496
rect 71832 491484 71838 491496
rect 76742 491484 76748 491496
rect 71832 491456 76748 491484
rect 71832 491444 71838 491456
rect 76742 491444 76748 491456
rect 76800 491444 76806 491496
rect 86770 491444 86776 491496
rect 86828 491484 86834 491496
rect 96430 491484 96436 491496
rect 86828 491456 96436 491484
rect 86828 491444 86834 491456
rect 96430 491444 96436 491456
rect 96488 491444 96494 491496
rect 99006 491444 99012 491496
rect 99064 491484 99070 491496
rect 110414 491484 110420 491496
rect 99064 491456 110420 491484
rect 99064 491444 99070 491456
rect 110414 491444 110420 491456
rect 110472 491444 110478 491496
rect 54846 491376 54852 491428
rect 54904 491416 54910 491428
rect 65610 491416 65616 491428
rect 54904 491388 65616 491416
rect 54904 491376 54910 491388
rect 65610 491376 65616 491388
rect 65668 491416 65674 491428
rect 65978 491416 65984 491428
rect 65668 491388 65984 491416
rect 65668 491376 65674 491388
rect 65978 491376 65984 491388
rect 66036 491376 66042 491428
rect 98362 491376 98368 491428
rect 98420 491416 98426 491428
rect 113450 491416 113456 491428
rect 98420 491388 113456 491416
rect 98420 491376 98426 491388
rect 113450 491376 113456 491388
rect 113508 491416 113514 491428
rect 114462 491416 114468 491428
rect 113508 491388 114468 491416
rect 113508 491376 113514 491388
rect 114462 491376 114468 491388
rect 114520 491376 114526 491428
rect 80054 491348 80060 491360
rect 48976 491320 80060 491348
rect 48976 491292 49004 491320
rect 80054 491308 80060 491320
rect 80112 491308 80118 491360
rect 93854 491308 93860 491360
rect 93912 491348 93918 491360
rect 99282 491348 99288 491360
rect 93912 491320 99288 491348
rect 93912 491308 93918 491320
rect 99282 491308 99288 491320
rect 99340 491308 99346 491360
rect 99650 491308 99656 491360
rect 99708 491348 99714 491360
rect 114554 491348 114560 491360
rect 99708 491320 114560 491348
rect 99708 491308 99714 491320
rect 114554 491308 114560 491320
rect 114612 491308 114618 491360
rect 46842 491240 46848 491292
rect 46900 491280 46906 491292
rect 48958 491280 48964 491292
rect 46900 491252 48964 491280
rect 46900 491240 46906 491252
rect 48958 491240 48964 491252
rect 49016 491240 49022 491292
rect 96522 491240 96528 491292
rect 96580 491280 96586 491292
rect 115106 491280 115112 491292
rect 96580 491252 115112 491280
rect 96580 491240 96586 491252
rect 115106 491240 115112 491252
rect 115164 491280 115170 491292
rect 118878 491280 118884 491292
rect 115164 491252 118884 491280
rect 115164 491240 115170 491252
rect 118878 491240 118884 491252
rect 118936 491240 118942 491292
rect 110414 491172 110420 491224
rect 110472 491212 110478 491224
rect 111702 491212 111708 491224
rect 110472 491184 111708 491212
rect 110472 491172 110478 491184
rect 111702 491172 111708 491184
rect 111760 491212 111766 491224
rect 127066 491212 127072 491224
rect 111760 491184 127072 491212
rect 111760 491172 111766 491184
rect 127066 491172 127072 491184
rect 127124 491172 127130 491224
rect 89898 490696 89904 490748
rect 89956 490736 89962 490748
rect 99374 490736 99380 490748
rect 89956 490708 99380 490736
rect 89956 490696 89962 490708
rect 99374 490696 99380 490708
rect 99432 490696 99438 490748
rect 58986 490628 58992 490680
rect 59044 490668 59050 490680
rect 79042 490668 79048 490680
rect 59044 490640 79048 490668
rect 59044 490628 59050 490640
rect 79042 490628 79048 490640
rect 79100 490628 79106 490680
rect 96246 490628 96252 490680
rect 96304 490668 96310 490680
rect 113358 490668 113364 490680
rect 96304 490640 113364 490668
rect 96304 490628 96310 490640
rect 113358 490628 113364 490640
rect 113416 490628 113422 490680
rect 42610 490560 42616 490612
rect 42668 490600 42674 490612
rect 49602 490600 49608 490612
rect 42668 490572 49608 490600
rect 42668 490560 42674 490572
rect 49602 490560 49608 490572
rect 49660 490600 49666 490612
rect 73246 490600 73252 490612
rect 49660 490572 73252 490600
rect 49660 490560 49666 490572
rect 73246 490560 73252 490572
rect 73304 490560 73310 490612
rect 86862 490560 86868 490612
rect 86920 490600 86926 490612
rect 109126 490600 109132 490612
rect 86920 490572 109132 490600
rect 86920 490560 86926 490572
rect 109126 490560 109132 490572
rect 109184 490560 109190 490612
rect 104894 489920 104900 489932
rect 91572 489892 104900 489920
rect 91572 489864 91600 489892
rect 104894 489880 104900 489892
rect 104952 489880 104958 489932
rect 35802 489812 35808 489864
rect 35860 489852 35866 489864
rect 67634 489852 67640 489864
rect 35860 489824 67640 489852
rect 35860 489812 35866 489824
rect 67634 489812 67640 489824
rect 67692 489812 67698 489864
rect 91554 489812 91560 489864
rect 91612 489812 91618 489864
rect 102042 489812 102048 489864
rect 102100 489852 102106 489864
rect 109034 489852 109040 489864
rect 102100 489824 109040 489852
rect 102100 489812 102106 489824
rect 109034 489812 109040 489824
rect 109092 489812 109098 489864
rect 109310 489812 109316 489864
rect 109368 489852 109374 489864
rect 118786 489852 118792 489864
rect 109368 489824 118792 489852
rect 109368 489812 109374 489824
rect 118786 489812 118792 489824
rect 118844 489852 118850 489864
rect 121454 489852 121460 489864
rect 118844 489824 121460 489852
rect 118844 489812 118850 489824
rect 121454 489812 121460 489824
rect 121512 489812 121518 489864
rect 103422 489132 103428 489184
rect 103480 489172 103486 489184
rect 117406 489172 117412 489184
rect 103480 489144 117412 489172
rect 103480 489132 103486 489144
rect 117406 489132 117412 489144
rect 117464 489132 117470 489184
rect 121454 489132 121460 489184
rect 121512 489172 121518 489184
rect 579614 489172 579620 489184
rect 121512 489144 579620 489172
rect 121512 489132 121518 489144
rect 579614 489132 579620 489144
rect 579672 489132 579678 489184
rect 34330 488520 34336 488572
rect 34388 488560 34394 488572
rect 35802 488560 35808 488572
rect 34388 488532 35808 488560
rect 34388 488520 34394 488532
rect 35802 488520 35808 488532
rect 35860 488520 35866 488572
rect 103422 488452 103428 488504
rect 103480 488492 103486 488504
rect 111794 488492 111800 488504
rect 103480 488464 111800 488492
rect 103480 488452 103486 488464
rect 111794 488452 111800 488464
rect 111852 488452 111858 488504
rect 109034 488384 109040 488436
rect 109092 488424 109098 488436
rect 110322 488424 110328 488436
rect 109092 488396 110328 488424
rect 109092 488384 109098 488396
rect 110322 488384 110328 488396
rect 110380 488424 110386 488436
rect 117314 488424 117320 488436
rect 110380 488396 117320 488424
rect 110380 488384 110386 488396
rect 117314 488384 117320 488396
rect 117372 488384 117378 488436
rect 111794 487840 111800 487892
rect 111852 487880 111858 487892
rect 128446 487880 128452 487892
rect 111852 487852 128452 487880
rect 111852 487840 111858 487852
rect 128446 487840 128452 487852
rect 128504 487840 128510 487892
rect 48222 487772 48228 487824
rect 48280 487812 48286 487824
rect 57790 487812 57796 487824
rect 48280 487784 57796 487812
rect 48280 487772 48286 487784
rect 57790 487772 57796 487784
rect 57848 487772 57854 487824
rect 103422 487772 103428 487824
rect 103480 487812 103486 487824
rect 133138 487812 133144 487824
rect 103480 487784 133144 487812
rect 103480 487772 103486 487784
rect 133138 487772 133144 487784
rect 133196 487812 133202 487824
rect 136726 487812 136732 487824
rect 133196 487784 136732 487812
rect 133196 487772 133202 487784
rect 136726 487772 136732 487784
rect 136784 487772 136790 487824
rect 114554 487500 114560 487552
rect 114612 487540 114618 487552
rect 118786 487540 118792 487552
rect 114612 487512 118792 487540
rect 114612 487500 114618 487512
rect 118786 487500 118792 487512
rect 118844 487500 118850 487552
rect 57606 487160 57612 487212
rect 57664 487200 57670 487212
rect 57790 487200 57796 487212
rect 57664 487172 57796 487200
rect 57664 487160 57670 487172
rect 57790 487160 57796 487172
rect 57848 487200 57854 487212
rect 67634 487200 67640 487212
rect 57848 487172 67640 487200
rect 57848 487160 57854 487172
rect 67634 487160 67640 487172
rect 67692 487160 67698 487212
rect 103422 487092 103428 487144
rect 103480 487132 103486 487144
rect 135254 487132 135260 487144
rect 103480 487104 135260 487132
rect 103480 487092 103486 487104
rect 135254 487092 135260 487104
rect 135312 487132 135318 487144
rect 136542 487132 136548 487144
rect 135312 487104 136548 487132
rect 135312 487092 135318 487104
rect 136542 487092 136548 487104
rect 136600 487092 136606 487144
rect 136542 486480 136548 486532
rect 136600 486520 136606 486532
rect 150526 486520 150532 486532
rect 136600 486492 150532 486520
rect 136600 486480 136606 486492
rect 150526 486480 150532 486492
rect 150584 486480 150590 486532
rect 41230 486412 41236 486464
rect 41288 486452 41294 486464
rect 67634 486452 67640 486464
rect 41288 486424 67640 486452
rect 41288 486412 41294 486424
rect 67634 486412 67640 486424
rect 67692 486412 67698 486464
rect 103422 486412 103428 486464
rect 103480 486452 103486 486464
rect 106182 486452 106188 486464
rect 103480 486424 106188 486452
rect 103480 486412 103486 486424
rect 106182 486412 106188 486424
rect 106240 486452 106246 486464
rect 135346 486452 135352 486464
rect 106240 486424 135352 486452
rect 106240 486412 106246 486424
rect 135346 486412 135352 486424
rect 135404 486412 135410 486464
rect 65610 485840 65616 485852
rect 64846 485812 65616 485840
rect 50798 485732 50804 485784
rect 50856 485772 50862 485784
rect 64846 485772 64874 485812
rect 65610 485800 65616 485812
rect 65668 485840 65674 485852
rect 67634 485840 67640 485852
rect 65668 485812 67640 485840
rect 65668 485800 65674 485812
rect 67634 485800 67640 485812
rect 67692 485800 67698 485852
rect 50856 485744 64874 485772
rect 50856 485732 50862 485744
rect 102134 485052 102140 485104
rect 102192 485092 102198 485104
rect 111794 485092 111800 485104
rect 102192 485064 111800 485092
rect 102192 485052 102198 485064
rect 111794 485052 111800 485064
rect 111852 485092 111858 485104
rect 112622 485092 112628 485104
rect 111852 485064 112628 485092
rect 111852 485052 111858 485064
rect 112622 485052 112628 485064
rect 112680 485052 112686 485104
rect 67266 484576 67272 484628
rect 67324 484616 67330 484628
rect 68646 484616 68652 484628
rect 67324 484588 68652 484616
rect 67324 484576 67330 484588
rect 68646 484576 68652 484588
rect 68704 484576 68710 484628
rect 47578 484480 47584 484492
rect 46952 484452 47584 484480
rect 44082 484304 44088 484356
rect 44140 484344 44146 484356
rect 46952 484344 46980 484452
rect 47578 484440 47584 484452
rect 47636 484480 47642 484492
rect 67634 484480 67640 484492
rect 47636 484452 67640 484480
rect 47636 484440 47642 484452
rect 67634 484440 67640 484452
rect 67692 484440 67698 484492
rect 99650 484372 99656 484424
rect 99708 484412 99714 484424
rect 112530 484412 112536 484424
rect 99708 484384 112536 484412
rect 99708 484372 99714 484384
rect 112530 484372 112536 484384
rect 112588 484372 112594 484424
rect 112622 484372 112628 484424
rect 112680 484412 112686 484424
rect 121454 484412 121460 484424
rect 112680 484384 121460 484412
rect 112680 484372 112686 484384
rect 121454 484372 121460 484384
rect 121512 484372 121518 484424
rect 44140 484316 46980 484344
rect 44140 484304 44146 484316
rect 56226 484304 56232 484356
rect 56284 484344 56290 484356
rect 56502 484344 56508 484356
rect 56284 484316 56508 484344
rect 56284 484304 56290 484316
rect 56502 484304 56508 484316
rect 56560 484304 56566 484356
rect 99926 484304 99932 484356
rect 99984 484344 99990 484356
rect 103514 484344 103520 484356
rect 99984 484316 103520 484344
rect 99984 484304 99990 484316
rect 103514 484304 103520 484316
rect 103572 484304 103578 484356
rect 56226 483624 56232 483676
rect 56284 483664 56290 483676
rect 67634 483664 67640 483676
rect 56284 483636 67640 483664
rect 56284 483624 56290 483636
rect 67634 483624 67640 483636
rect 67692 483624 67698 483676
rect 102134 483624 102140 483676
rect 102192 483664 102198 483676
rect 122926 483664 122932 483676
rect 102192 483636 122932 483664
rect 102192 483624 102198 483636
rect 122926 483624 122932 483636
rect 122984 483624 122990 483676
rect 36998 483012 37004 483064
rect 37056 483052 37062 483064
rect 137278 483052 137284 483064
rect 37056 483024 52500 483052
rect 137191 483024 137284 483052
rect 37056 483012 37062 483024
rect 52472 482984 52500 483024
rect 137278 483012 137284 483024
rect 137336 483052 137342 483064
rect 147950 483052 147956 483064
rect 137336 483024 147956 483052
rect 137336 483012 137342 483024
rect 147950 483012 147956 483024
rect 148008 483012 148014 483064
rect 53098 482984 53104 482996
rect 52472 482956 53104 482984
rect 53098 482944 53104 482956
rect 53156 482984 53162 482996
rect 67634 482984 67640 482996
rect 53156 482956 67640 482984
rect 53156 482944 53162 482956
rect 67634 482944 67640 482956
rect 67692 482944 67698 482996
rect 102134 482944 102140 482996
rect 102192 482984 102198 482996
rect 137296 482984 137324 483012
rect 102192 482956 137324 482984
rect 102192 482944 102198 482956
rect 48038 481652 48044 481704
rect 48096 481692 48102 481704
rect 65518 481692 65524 481704
rect 48096 481664 65524 481692
rect 48096 481652 48102 481664
rect 65518 481652 65524 481664
rect 65576 481692 65582 481704
rect 65978 481692 65984 481704
rect 65576 481664 65984 481692
rect 65576 481652 65582 481664
rect 65978 481652 65984 481664
rect 66036 481652 66042 481704
rect 102134 481652 102140 481704
rect 102192 481692 102198 481704
rect 117038 481692 117044 481704
rect 102192 481664 117044 481692
rect 102192 481652 102198 481664
rect 117038 481652 117044 481664
rect 117096 481652 117102 481704
rect 64598 481584 64604 481636
rect 64656 481624 64662 481636
rect 68002 481624 68008 481636
rect 64656 481596 68008 481624
rect 64656 481584 64662 481596
rect 68002 481584 68008 481596
rect 68060 481584 68066 481636
rect 102318 481584 102324 481636
rect 102376 481624 102382 481636
rect 128630 481624 128636 481636
rect 102376 481596 128636 481624
rect 102376 481584 102382 481596
rect 128630 481584 128636 481596
rect 128688 481584 128694 481636
rect 65978 481516 65984 481568
rect 66036 481556 66042 481568
rect 67634 481556 67640 481568
rect 66036 481528 67640 481556
rect 66036 481516 66042 481528
rect 67634 481516 67640 481528
rect 67692 481516 67698 481568
rect 102134 480904 102140 480956
rect 102192 480944 102198 480956
rect 113174 480944 113180 480956
rect 102192 480916 113180 480944
rect 102192 480904 102198 480916
rect 113174 480904 113180 480916
rect 113232 480904 113238 480956
rect 128630 480904 128636 480956
rect 128688 480944 128694 480956
rect 146294 480944 146300 480956
rect 128688 480916 146300 480944
rect 128688 480904 128694 480916
rect 146294 480904 146300 480916
rect 146352 480904 146358 480956
rect 59170 480156 59176 480208
rect 59228 480196 59234 480208
rect 67634 480196 67640 480208
rect 59228 480168 67640 480196
rect 59228 480156 59234 480168
rect 67634 480156 67640 480168
rect 67692 480156 67698 480208
rect 102134 480156 102140 480208
rect 102192 480196 102198 480208
rect 140774 480196 140780 480208
rect 102192 480168 140780 480196
rect 102192 480156 102198 480168
rect 140774 480156 140780 480168
rect 140832 480156 140838 480208
rect 102134 479680 102140 479732
rect 102192 479720 102198 479732
rect 104986 479720 104992 479732
rect 102192 479692 104992 479720
rect 102192 479680 102198 479692
rect 104986 479680 104992 479692
rect 105044 479720 105050 479732
rect 106182 479720 106188 479732
rect 105044 479692 106188 479720
rect 105044 479680 105050 479692
rect 106182 479680 106188 479692
rect 106240 479680 106246 479732
rect 112530 479476 112536 479528
rect 112588 479516 112594 479528
rect 117314 479516 117320 479528
rect 112588 479488 117320 479516
rect 112588 479476 112594 479488
rect 117314 479476 117320 479488
rect 117372 479476 117378 479528
rect 140774 479476 140780 479528
rect 140832 479516 140838 479528
rect 145006 479516 145012 479528
rect 140832 479488 145012 479516
rect 140832 479476 140838 479488
rect 145006 479476 145012 479488
rect 145064 479476 145070 479528
rect 109770 478864 109776 478916
rect 109828 478904 109834 478916
rect 136634 478904 136640 478916
rect 109828 478876 136640 478904
rect 109828 478864 109834 478876
rect 136634 478864 136640 478876
rect 136692 478864 136698 478916
rect 63034 477572 63040 477624
rect 63092 477612 63098 477624
rect 63218 477612 63224 477624
rect 63092 477584 63224 477612
rect 63092 477572 63098 477584
rect 63218 477572 63224 477584
rect 63276 477572 63282 477624
rect 102134 477504 102140 477556
rect 102192 477544 102198 477556
rect 115842 477544 115848 477556
rect 102192 477516 115848 477544
rect 102192 477504 102198 477516
rect 115842 477504 115848 477516
rect 115900 477504 115906 477556
rect 61746 477436 61752 477488
rect 61804 477476 61810 477488
rect 63218 477476 63224 477488
rect 61804 477448 63224 477476
rect 61804 477436 61810 477448
rect 63218 477436 63224 477448
rect 63276 477476 63282 477488
rect 67726 477476 67732 477488
rect 63276 477448 67732 477476
rect 63276 477436 63282 477448
rect 67726 477436 67732 477448
rect 67784 477436 67790 477488
rect 102318 477436 102324 477488
rect 102376 477476 102382 477488
rect 114738 477476 114744 477488
rect 102376 477448 114744 477476
rect 102376 477436 102382 477448
rect 114738 477436 114744 477448
rect 114796 477476 114802 477488
rect 116026 477476 116032 477488
rect 114796 477448 116032 477476
rect 114796 477436 114802 477448
rect 116026 477436 116032 477448
rect 116084 477436 116090 477488
rect 102134 477368 102140 477420
rect 102192 477408 102198 477420
rect 109770 477408 109776 477420
rect 102192 477380 109776 477408
rect 102192 477368 102198 477380
rect 109770 477368 109776 477380
rect 109828 477368 109834 477420
rect 106182 476756 106188 476808
rect 106240 476796 106246 476808
rect 151814 476796 151820 476808
rect 106240 476768 151820 476796
rect 106240 476756 106246 476768
rect 151814 476756 151820 476768
rect 151872 476756 151878 476808
rect 35802 476076 35808 476128
rect 35860 476116 35866 476128
rect 67634 476116 67640 476128
rect 35860 476088 67640 476116
rect 35860 476076 35866 476088
rect 67634 476076 67640 476088
rect 67692 476076 67698 476128
rect 117958 476076 117964 476128
rect 118016 476116 118022 476128
rect 120166 476116 120172 476128
rect 118016 476088 120172 476116
rect 118016 476076 118022 476088
rect 120166 476076 120172 476088
rect 120224 476076 120230 476128
rect 102410 476008 102416 476060
rect 102468 476048 102474 476060
rect 103422 476048 103428 476060
rect 102468 476020 103428 476048
rect 102468 476008 102474 476020
rect 103422 476008 103428 476020
rect 103480 476048 103486 476060
rect 142154 476048 142160 476060
rect 103480 476020 142160 476048
rect 103480 476008 103486 476020
rect 142154 476008 142160 476020
rect 142212 476008 142218 476060
rect 102318 475940 102324 475992
rect 102376 475980 102382 475992
rect 125778 475980 125784 475992
rect 102376 475952 125784 475980
rect 102376 475940 102382 475952
rect 125778 475940 125784 475952
rect 125836 475980 125842 475992
rect 131758 475980 131764 475992
rect 125836 475952 131764 475980
rect 125836 475940 125842 475952
rect 131758 475940 131764 475952
rect 131816 475940 131822 475992
rect 102134 475872 102140 475924
rect 102192 475912 102198 475924
rect 117958 475912 117964 475924
rect 102192 475884 117964 475912
rect 102192 475872 102198 475884
rect 117958 475872 117964 475884
rect 118016 475872 118022 475924
rect 55950 475328 55956 475380
rect 56008 475368 56014 475380
rect 56318 475368 56324 475380
rect 56008 475340 56324 475368
rect 56008 475328 56014 475340
rect 56318 475328 56324 475340
rect 56376 475368 56382 475380
rect 67634 475368 67640 475380
rect 56376 475340 67640 475368
rect 56376 475328 56382 475340
rect 67634 475328 67640 475340
rect 67692 475328 67698 475380
rect 105630 474852 105636 474904
rect 105688 474892 105694 474904
rect 107930 474892 107936 474904
rect 105688 474864 107936 474892
rect 105688 474852 105694 474864
rect 107930 474852 107936 474864
rect 107988 474852 107994 474904
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 25498 474756 25504 474768
rect 3476 474728 25504 474756
rect 3476 474716 3482 474728
rect 25498 474716 25504 474728
rect 25556 474716 25562 474768
rect 67634 474756 67640 474768
rect 64800 474728 67640 474756
rect 34422 474648 34428 474700
rect 34480 474688 34486 474700
rect 64230 474688 64236 474700
rect 34480 474660 64236 474688
rect 34480 474648 34486 474660
rect 64230 474648 64236 474660
rect 64288 474688 64294 474700
rect 64800 474688 64828 474728
rect 67634 474716 67640 474728
rect 67692 474716 67698 474768
rect 64288 474660 64828 474688
rect 64288 474648 64294 474660
rect 102134 474648 102140 474700
rect 102192 474688 102198 474700
rect 142246 474688 142252 474700
rect 102192 474660 142252 474688
rect 102192 474648 102198 474660
rect 142246 474648 142252 474660
rect 142304 474688 142310 474700
rect 150618 474688 150624 474700
rect 142304 474660 150624 474688
rect 142304 474648 142310 474660
rect 150618 474648 150624 474660
rect 150676 474648 150682 474700
rect 66070 473288 66076 473340
rect 66128 473328 66134 473340
rect 67634 473328 67640 473340
rect 66128 473300 67640 473328
rect 66128 473288 66134 473300
rect 67634 473288 67640 473300
rect 67692 473288 67698 473340
rect 102318 473288 102324 473340
rect 102376 473328 102382 473340
rect 106366 473328 106372 473340
rect 102376 473300 106372 473328
rect 102376 473288 102382 473300
rect 106366 473288 106372 473300
rect 106424 473328 106430 473340
rect 107562 473328 107568 473340
rect 106424 473300 107568 473328
rect 106424 473288 106430 473300
rect 107562 473288 107568 473300
rect 107620 473288 107626 473340
rect 99558 472744 99564 472796
rect 99616 472784 99622 472796
rect 110598 472784 110604 472796
rect 99616 472756 110604 472784
rect 99616 472744 99622 472756
rect 110598 472744 110604 472756
rect 110656 472744 110662 472796
rect 107562 472676 107568 472728
rect 107620 472716 107626 472728
rect 118878 472716 118884 472728
rect 107620 472688 118884 472716
rect 107620 472676 107626 472688
rect 118878 472676 118884 472688
rect 118936 472676 118942 472728
rect 48222 472608 48228 472660
rect 48280 472648 48286 472660
rect 66070 472648 66076 472660
rect 48280 472620 66076 472648
rect 48280 472608 48286 472620
rect 66070 472608 66076 472620
rect 66128 472608 66134 472660
rect 102134 472608 102140 472660
rect 102192 472648 102198 472660
rect 133874 472648 133880 472660
rect 102192 472620 133880 472648
rect 102192 472608 102198 472620
rect 133874 472608 133880 472620
rect 133932 472608 133938 472660
rect 102134 471928 102140 471980
rect 102192 471968 102198 471980
rect 124306 471968 124312 471980
rect 102192 471940 124312 471968
rect 102192 471928 102198 471940
rect 124306 471928 124312 471940
rect 124364 471968 124370 471980
rect 129734 471968 129740 471980
rect 124364 471940 129740 471968
rect 124364 471928 124370 471940
rect 129734 471928 129740 471940
rect 129792 471928 129798 471980
rect 64966 471588 64972 471640
rect 65024 471628 65030 471640
rect 67634 471628 67640 471640
rect 65024 471600 67640 471628
rect 65024 471588 65030 471600
rect 67634 471588 67640 471600
rect 67692 471588 67698 471640
rect 118878 471316 118884 471368
rect 118936 471356 118942 471368
rect 146386 471356 146392 471368
rect 118936 471328 146392 471356
rect 118936 471316 118942 471328
rect 146386 471316 146392 471328
rect 146444 471316 146450 471368
rect 50798 471248 50804 471300
rect 50856 471288 50862 471300
rect 63034 471288 63040 471300
rect 50856 471260 63040 471288
rect 50856 471248 50862 471260
rect 63034 471248 63040 471260
rect 63092 471288 63098 471300
rect 67634 471288 67640 471300
rect 63092 471260 67640 471288
rect 63092 471248 63098 471260
rect 67634 471248 67640 471260
rect 67692 471248 67698 471300
rect 102870 471248 102876 471300
rect 102928 471288 102934 471300
rect 139486 471288 139492 471300
rect 102928 471260 139492 471288
rect 102928 471248 102934 471260
rect 139486 471248 139492 471260
rect 139544 471248 139550 471300
rect 59078 470568 59084 470620
rect 59136 470608 59142 470620
rect 64966 470608 64972 470620
rect 59136 470580 64972 470608
rect 59136 470568 59142 470580
rect 64966 470568 64972 470580
rect 65024 470568 65030 470620
rect 102318 470568 102324 470620
rect 102376 470608 102382 470620
rect 107562 470608 107568 470620
rect 102376 470580 107568 470608
rect 102376 470568 102382 470580
rect 107562 470568 107568 470580
rect 107620 470608 107626 470620
rect 112622 470608 112628 470620
rect 107620 470580 112628 470608
rect 107620 470568 107626 470580
rect 112622 470568 112628 470580
rect 112680 470568 112686 470620
rect 139486 470568 139492 470620
rect 139544 470608 139550 470620
rect 142338 470608 142344 470620
rect 139544 470580 142344 470608
rect 139544 470568 139550 470580
rect 142338 470568 142344 470580
rect 142396 470568 142402 470620
rect 146386 470568 146392 470620
rect 146444 470608 146450 470620
rect 579890 470608 579896 470620
rect 146444 470580 579896 470608
rect 146444 470568 146450 470580
rect 579890 470568 579896 470580
rect 579948 470568 579954 470620
rect 102134 470500 102140 470552
rect 102192 470540 102198 470552
rect 130010 470540 130016 470552
rect 102192 470512 130016 470540
rect 102192 470500 102198 470512
rect 130010 470500 130016 470512
rect 130068 470500 130074 470552
rect 130010 469888 130016 469940
rect 130068 469928 130074 469940
rect 151998 469928 152004 469940
rect 130068 469900 152004 469928
rect 130068 469888 130074 469900
rect 151998 469888 152004 469900
rect 152056 469888 152062 469940
rect 103606 469820 103612 469872
rect 103664 469860 103670 469872
rect 138106 469860 138112 469872
rect 103664 469832 138112 469860
rect 103664 469820 103670 469832
rect 138106 469820 138112 469832
rect 138164 469860 138170 469872
rect 142246 469860 142252 469872
rect 138164 469832 142252 469860
rect 138164 469820 138170 469832
rect 142246 469820 142252 469832
rect 142304 469820 142310 469872
rect 64506 469480 64512 469532
rect 64564 469520 64570 469532
rect 66162 469520 66168 469532
rect 64564 469492 66168 469520
rect 64564 469480 64570 469492
rect 66162 469480 66168 469492
rect 66220 469520 66226 469532
rect 67726 469520 67732 469532
rect 66220 469492 67732 469520
rect 66220 469480 66226 469492
rect 67726 469480 67732 469492
rect 67784 469480 67790 469532
rect 43806 469208 43812 469260
rect 43864 469248 43870 469260
rect 66070 469248 66076 469260
rect 43864 469220 66076 469248
rect 43864 469208 43870 469220
rect 66070 469208 66076 469220
rect 66128 469248 66134 469260
rect 67634 469248 67640 469260
rect 66128 469220 67640 469248
rect 66128 469208 66134 469220
rect 67634 469208 67640 469220
rect 67692 469208 67698 469260
rect 64690 469072 64696 469124
rect 64748 469112 64754 469124
rect 66070 469112 66076 469124
rect 64748 469084 66076 469112
rect 64748 469072 64754 469084
rect 66070 469072 66076 469084
rect 66128 469072 66134 469124
rect 66070 468188 66076 468240
rect 66128 468228 66134 468240
rect 67634 468228 67640 468240
rect 66128 468200 67640 468228
rect 66128 468188 66134 468200
rect 67634 468188 67640 468200
rect 67692 468188 67698 468240
rect 60366 467848 60372 467900
rect 60424 467888 60430 467900
rect 63310 467888 63316 467900
rect 60424 467860 63316 467888
rect 60424 467848 60430 467860
rect 63310 467848 63316 467860
rect 63368 467888 63374 467900
rect 67726 467888 67732 467900
rect 63368 467860 67732 467888
rect 63368 467848 63374 467860
rect 67726 467848 67732 467860
rect 67784 467848 67790 467900
rect 61746 466760 61752 466812
rect 61804 466800 61810 466812
rect 63126 466800 63132 466812
rect 61804 466772 63132 466800
rect 61804 466760 61810 466772
rect 63126 466760 63132 466772
rect 63184 466800 63190 466812
rect 67634 466800 67640 466812
rect 63184 466772 67640 466800
rect 63184 466760 63190 466772
rect 67634 466760 67640 466772
rect 67692 466760 67698 466812
rect 102134 466488 102140 466540
rect 102192 466528 102198 466540
rect 115198 466528 115204 466540
rect 102192 466500 115204 466528
rect 102192 466488 102198 466500
rect 115198 466488 115204 466500
rect 115256 466528 115262 466540
rect 115842 466528 115848 466540
rect 115256 466500 115848 466528
rect 115256 466488 115262 466500
rect 115842 466488 115848 466500
rect 115900 466488 115906 466540
rect 103146 466420 103152 466472
rect 103204 466460 103210 466472
rect 103204 466432 118740 466460
rect 103204 466420 103210 466432
rect 102134 466352 102140 466404
rect 102192 466392 102198 466404
rect 118712 466392 118740 466432
rect 119982 466392 119988 466404
rect 102192 466364 103514 466392
rect 118712 466364 119988 466392
rect 102192 466352 102198 466364
rect 103486 466256 103514 466364
rect 119982 466352 119988 466364
rect 120040 466392 120046 466404
rect 136818 466392 136824 466404
rect 120040 466364 136824 466392
rect 120040 466352 120046 466364
rect 136818 466352 136824 466364
rect 136876 466352 136882 466404
rect 115842 466284 115848 466336
rect 115900 466324 115906 466336
rect 124214 466324 124220 466336
rect 115900 466296 124220 466324
rect 115900 466284 115906 466296
rect 124214 466284 124220 466296
rect 124272 466284 124278 466336
rect 114646 466256 114652 466268
rect 103486 466228 114652 466256
rect 114646 466216 114652 466228
rect 114704 466256 114710 466268
rect 121730 466256 121736 466268
rect 114704 466228 121736 466256
rect 114704 466216 114710 466228
rect 121730 466216 121736 466228
rect 121788 466216 121794 466268
rect 102134 465672 102140 465724
rect 102192 465712 102198 465724
rect 103330 465712 103336 465724
rect 102192 465684 103336 465712
rect 102192 465672 102198 465684
rect 103330 465672 103336 465684
rect 103388 465712 103394 465724
rect 107746 465712 107752 465724
rect 103388 465684 107752 465712
rect 103388 465672 103394 465684
rect 107746 465672 107752 465684
rect 107804 465672 107810 465724
rect 65518 465100 65524 465112
rect 64846 465072 65524 465100
rect 57698 464992 57704 465044
rect 57756 465032 57762 465044
rect 64846 465032 64874 465072
rect 65518 465060 65524 465072
rect 65576 465100 65582 465112
rect 67726 465100 67732 465112
rect 65576 465072 67732 465100
rect 65576 465060 65582 465072
rect 67726 465060 67732 465072
rect 67784 465060 67790 465112
rect 127618 465100 127624 465112
rect 127531 465072 127624 465100
rect 127618 465060 127624 465072
rect 127676 465100 127682 465112
rect 138106 465100 138112 465112
rect 127676 465072 138112 465100
rect 127676 465060 127682 465072
rect 138106 465060 138112 465072
rect 138164 465060 138170 465112
rect 57756 465004 64874 465032
rect 57756 464992 57762 465004
rect 102134 464992 102140 465044
rect 102192 465032 102198 465044
rect 127636 465032 127664 465060
rect 102192 465004 127664 465032
rect 102192 464992 102198 465004
rect 101398 464924 101404 464976
rect 101456 464964 101462 464976
rect 102226 464964 102232 464976
rect 101456 464936 102232 464964
rect 101456 464924 101462 464936
rect 102226 464924 102232 464936
rect 102284 464924 102290 464976
rect 108482 464380 108488 464432
rect 108540 464420 108546 464432
rect 111978 464420 111984 464432
rect 108540 464392 111984 464420
rect 108540 464380 108546 464392
rect 111978 464380 111984 464392
rect 112036 464380 112042 464432
rect 427814 464312 427820 464364
rect 427872 464352 427878 464364
rect 497458 464352 497464 464364
rect 427872 464324 497464 464352
rect 427872 464312 427878 464324
rect 497458 464312 497464 464324
rect 497516 464312 497522 464364
rect 102134 464108 102140 464160
rect 102192 464148 102198 464160
rect 105630 464148 105636 464160
rect 102192 464120 105636 464148
rect 102192 464108 102198 464120
rect 105630 464108 105636 464120
rect 105688 464108 105694 464160
rect 60458 463768 60464 463820
rect 60516 463808 60522 463820
rect 64138 463808 64144 463820
rect 60516 463780 64144 463808
rect 60516 463768 60522 463780
rect 64138 463768 64144 463780
rect 64196 463808 64202 463820
rect 67634 463808 67640 463820
rect 64196 463780 67640 463808
rect 64196 463768 64202 463780
rect 67634 463768 67640 463780
rect 67692 463768 67698 463820
rect 67818 463740 67824 463752
rect 53576 463712 67824 463740
rect 52270 463632 52276 463684
rect 52328 463672 52334 463684
rect 53098 463672 53104 463684
rect 52328 463644 53104 463672
rect 52328 463632 52334 463644
rect 53098 463632 53104 463644
rect 53156 463672 53162 463684
rect 53576 463672 53604 463712
rect 67818 463700 67824 463712
rect 67876 463700 67882 463752
rect 124214 463740 124220 463752
rect 120000 463712 124220 463740
rect 53156 463644 53604 463672
rect 53156 463632 53162 463644
rect 60458 463632 60464 463684
rect 60516 463672 60522 463684
rect 61838 463672 61844 463684
rect 60516 463644 61844 463672
rect 60516 463632 60522 463644
rect 61838 463632 61844 463644
rect 61896 463672 61902 463684
rect 67726 463672 67732 463684
rect 61896 463644 67732 463672
rect 61896 463632 61902 463644
rect 67726 463632 67732 463644
rect 67784 463632 67790 463684
rect 102134 463632 102140 463684
rect 102192 463672 102198 463684
rect 119430 463672 119436 463684
rect 102192 463644 119436 463672
rect 102192 463632 102198 463644
rect 119430 463632 119436 463644
rect 119488 463672 119494 463684
rect 120000 463672 120028 463712
rect 124214 463700 124220 463712
rect 124272 463700 124278 463752
rect 119488 463644 120028 463672
rect 119488 463632 119494 463644
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 67634 462380 67640 462392
rect 60752 462352 67640 462380
rect 52270 462272 52276 462324
rect 52328 462312 52334 462324
rect 53190 462312 53196 462324
rect 52328 462284 53196 462312
rect 52328 462272 52334 462284
rect 53190 462272 53196 462284
rect 53248 462272 53254 462324
rect 59170 462272 59176 462324
rect 59228 462312 59234 462324
rect 60752 462312 60780 462352
rect 67634 462340 67640 462352
rect 67692 462340 67698 462392
rect 107562 462340 107568 462392
rect 107620 462380 107626 462392
rect 140958 462380 140964 462392
rect 107620 462352 140964 462380
rect 107620 462340 107626 462352
rect 140958 462340 140964 462352
rect 141016 462340 141022 462392
rect 59228 462284 60780 462312
rect 59228 462272 59234 462284
rect 102226 462272 102232 462324
rect 102284 462312 102290 462324
rect 124398 462312 124404 462324
rect 102284 462284 124404 462312
rect 102284 462272 102290 462284
rect 124398 462272 124404 462284
rect 124456 462312 124462 462324
rect 125962 462312 125968 462324
rect 124456 462284 125968 462312
rect 124456 462272 124462 462284
rect 125962 462272 125968 462284
rect 126020 462272 126026 462324
rect 59262 462204 59268 462256
rect 59320 462244 59326 462256
rect 63218 462244 63224 462256
rect 59320 462216 63224 462244
rect 59320 462204 59326 462216
rect 63218 462204 63224 462216
rect 63276 462204 63282 462256
rect 102134 462204 102140 462256
rect 102192 462244 102198 462256
rect 107562 462244 107568 462256
rect 102192 462216 107568 462244
rect 102192 462204 102198 462216
rect 107562 462204 107568 462216
rect 107620 462204 107626 462256
rect 52178 461592 52184 461644
rect 52236 461632 52242 461644
rect 59170 461632 59176 461644
rect 52236 461604 59176 461632
rect 52236 461592 52242 461604
rect 59170 461592 59176 461604
rect 59228 461592 59234 461644
rect 63218 460912 63224 460964
rect 63276 460952 63282 460964
rect 67634 460952 67640 460964
rect 63276 460924 67640 460952
rect 63276 460912 63282 460924
rect 67634 460912 67640 460924
rect 67692 460912 67698 460964
rect 107010 460952 107016 460964
rect 106246 460924 107016 460952
rect 102134 460844 102140 460896
rect 102192 460884 102198 460896
rect 106246 460884 106274 460924
rect 107010 460912 107016 460924
rect 107068 460952 107074 460964
rect 147858 460952 147864 460964
rect 107068 460924 147864 460952
rect 107068 460912 107074 460924
rect 147858 460912 147864 460924
rect 147916 460912 147922 460964
rect 102192 460856 106274 460884
rect 102192 460844 102198 460856
rect 50982 460232 50988 460284
rect 51040 460272 51046 460284
rect 67634 460272 67640 460284
rect 51040 460244 67640 460272
rect 51040 460232 51046 460244
rect 67634 460232 67640 460244
rect 67692 460232 67698 460284
rect 42702 460164 42708 460216
rect 42760 460204 42766 460216
rect 67726 460204 67732 460216
rect 42760 460176 67732 460204
rect 42760 460164 42766 460176
rect 67726 460164 67732 460176
rect 67784 460164 67790 460216
rect 50706 459552 50712 459604
rect 50764 459592 50770 459604
rect 50982 459592 50988 459604
rect 50764 459564 50988 459592
rect 50764 459552 50770 459564
rect 50982 459552 50988 459564
rect 51040 459552 51046 459604
rect 102226 459552 102232 459604
rect 102284 459592 102290 459604
rect 107470 459592 107476 459604
rect 102284 459564 107476 459592
rect 102284 459552 102290 459564
rect 107470 459552 107476 459564
rect 107528 459592 107534 459604
rect 107528 459564 107608 459592
rect 107528 459552 107534 459564
rect 107580 459524 107608 459564
rect 116670 459552 116676 459604
rect 116728 459592 116734 459604
rect 133966 459592 133972 459604
rect 116728 459564 133972 459592
rect 116728 459552 116734 459564
rect 133966 459552 133972 459564
rect 134024 459552 134030 459604
rect 138014 459524 138020 459536
rect 107580 459496 138020 459524
rect 138014 459484 138020 459496
rect 138072 459484 138078 459536
rect 102134 459416 102140 459468
rect 102192 459456 102198 459468
rect 116670 459456 116676 459468
rect 102192 459428 116676 459456
rect 102192 459416 102198 459428
rect 116670 459416 116676 459428
rect 116728 459416 116734 459468
rect 35158 458872 35164 458924
rect 35216 458912 35222 458924
rect 42702 458912 42708 458924
rect 35216 458884 42708 458912
rect 35216 458872 35222 458884
rect 42702 458872 42708 458884
rect 42760 458872 42766 458924
rect 37090 458804 37096 458856
rect 37148 458844 37154 458856
rect 67450 458844 67456 458856
rect 37148 458816 67456 458844
rect 37148 458804 37154 458816
rect 67450 458804 67456 458816
rect 67508 458844 67514 458856
rect 67634 458844 67640 458856
rect 67508 458816 67640 458844
rect 67508 458804 67514 458816
rect 67634 458804 67640 458816
rect 67692 458804 67698 458856
rect 107562 458804 107568 458856
rect 107620 458844 107626 458856
rect 135438 458844 135444 458856
rect 107620 458816 135444 458844
rect 107620 458804 107626 458816
rect 135438 458804 135444 458816
rect 135496 458804 135502 458856
rect 33778 458300 33784 458312
rect 33336 458272 33784 458300
rect 30282 458124 30288 458176
rect 30340 458164 30346 458176
rect 33336 458164 33364 458272
rect 33778 458260 33784 458272
rect 33836 458300 33842 458312
rect 67634 458300 67640 458312
rect 33836 458272 67640 458300
rect 33836 458260 33842 458272
rect 67634 458260 67640 458272
rect 67692 458260 67698 458312
rect 135438 458192 135444 458244
rect 135496 458232 135502 458244
rect 139486 458232 139492 458244
rect 135496 458204 139492 458232
rect 135496 458192 135502 458204
rect 139486 458192 139492 458204
rect 139544 458192 139550 458244
rect 30340 458136 33364 458164
rect 30340 458124 30346 458136
rect 43714 458124 43720 458176
rect 43772 458164 43778 458176
rect 48130 458164 48136 458176
rect 43772 458136 48136 458164
rect 43772 458124 43778 458136
rect 48130 458124 48136 458136
rect 48188 458164 48194 458176
rect 67726 458164 67732 458176
rect 48188 458136 67732 458164
rect 48188 458124 48194 458136
rect 67726 458124 67732 458136
rect 67784 458124 67790 458176
rect 103238 458124 103244 458176
rect 103296 458164 103302 458176
rect 125594 458164 125600 458176
rect 103296 458136 125600 458164
rect 103296 458124 103302 458136
rect 125594 458124 125600 458136
rect 125652 458124 125658 458176
rect 102134 458056 102140 458108
rect 102192 458096 102198 458108
rect 107562 458096 107568 458108
rect 102192 458068 107568 458096
rect 102192 458056 102198 458068
rect 107562 458056 107568 458068
rect 107620 458056 107626 458108
rect 43898 457444 43904 457496
rect 43956 457484 43962 457496
rect 44082 457484 44088 457496
rect 43956 457456 44088 457484
rect 43956 457444 43962 457456
rect 44082 457444 44088 457456
rect 44140 457484 44146 457496
rect 67634 457484 67640 457496
rect 44140 457456 67640 457484
rect 44140 457444 44146 457456
rect 67634 457444 67640 457456
rect 67692 457444 67698 457496
rect 431954 457444 431960 457496
rect 432012 457484 432018 457496
rect 579614 457484 579620 457496
rect 432012 457456 579620 457484
rect 432012 457444 432018 457456
rect 579614 457444 579620 457456
rect 579672 457444 579678 457496
rect 106182 456764 106188 456816
rect 106240 456804 106246 456816
rect 151906 456804 151912 456816
rect 106240 456776 151912 456804
rect 106240 456764 106246 456776
rect 151906 456764 151912 456776
rect 151964 456764 151970 456816
rect 42426 456696 42432 456748
rect 42484 456736 42490 456748
rect 44082 456736 44088 456748
rect 42484 456708 44088 456736
rect 42484 456696 42490 456708
rect 44082 456696 44088 456708
rect 44140 456696 44146 456748
rect 102134 456696 102140 456748
rect 102192 456736 102198 456748
rect 139578 456736 139584 456748
rect 102192 456708 139584 456736
rect 102192 456696 102198 456708
rect 139578 456696 139584 456708
rect 139636 456736 139642 456748
rect 140314 456736 140320 456748
rect 139636 456708 140320 456736
rect 139636 456696 139642 456708
rect 140314 456696 140320 456708
rect 140372 456696 140378 456748
rect 102226 456628 102232 456680
rect 102284 456668 102290 456680
rect 105538 456668 105544 456680
rect 102284 456640 105544 456668
rect 102284 456628 102290 456640
rect 105538 456628 105544 456640
rect 105596 456668 105602 456680
rect 106182 456668 106188 456680
rect 105596 456640 106188 456668
rect 105596 456628 105602 456640
rect 106182 456628 106188 456640
rect 106240 456628 106246 456680
rect 35710 456016 35716 456068
rect 35768 456056 35774 456068
rect 67634 456056 67640 456068
rect 35768 456028 67640 456056
rect 35768 456016 35774 456028
rect 67634 456016 67640 456028
rect 67692 456016 67698 456068
rect 140314 456016 140320 456068
rect 140372 456056 140378 456068
rect 149146 456056 149152 456068
rect 140372 456028 149152 456056
rect 140372 456016 140378 456028
rect 149146 456016 149152 456028
rect 149204 456016 149210 456068
rect 105538 455948 105544 456000
rect 105596 455988 105602 456000
rect 109126 455988 109132 456000
rect 105596 455960 109132 455988
rect 105596 455948 105602 455960
rect 109126 455948 109132 455960
rect 109184 455948 109190 456000
rect 56502 455812 56508 455864
rect 56560 455852 56566 455864
rect 57974 455852 57980 455864
rect 56560 455824 57980 455852
rect 56560 455812 56566 455824
rect 57974 455812 57980 455824
rect 58032 455812 58038 455864
rect 132586 455444 132592 455456
rect 103486 455416 132592 455444
rect 35710 455336 35716 455388
rect 35768 455376 35774 455388
rect 36630 455376 36636 455388
rect 35768 455348 36636 455376
rect 35768 455336 35774 455348
rect 36630 455336 36636 455348
rect 36688 455336 36694 455388
rect 57974 455336 57980 455388
rect 58032 455376 58038 455388
rect 67634 455376 67640 455388
rect 58032 455348 67640 455376
rect 58032 455336 58038 455348
rect 67634 455336 67640 455348
rect 67692 455336 67698 455388
rect 102134 455336 102140 455388
rect 102192 455376 102198 455388
rect 103486 455376 103514 455416
rect 132586 455404 132592 455416
rect 132644 455404 132650 455456
rect 102192 455348 103514 455376
rect 102192 455336 102198 455348
rect 107654 455336 107660 455388
rect 107712 455376 107718 455388
rect 108298 455376 108304 455388
rect 107712 455348 108304 455376
rect 107712 455336 107718 455348
rect 108298 455336 108304 455348
rect 108356 455336 108362 455388
rect 102134 454792 102140 454844
rect 102192 454832 102198 454844
rect 107654 454832 107660 454844
rect 102192 454804 107660 454832
rect 102192 454792 102198 454804
rect 107654 454792 107660 454804
rect 107712 454792 107718 454844
rect 100662 454724 100668 454776
rect 100720 454764 100726 454776
rect 113174 454764 113180 454776
rect 100720 454736 113180 454764
rect 100720 454724 100726 454736
rect 113174 454724 113180 454736
rect 113232 454724 113238 454776
rect 106182 454656 106188 454708
rect 106240 454696 106246 454708
rect 134242 454696 134248 454708
rect 106240 454668 134248 454696
rect 106240 454656 106246 454668
rect 134242 454656 134248 454668
rect 134300 454696 134306 454708
rect 143718 454696 143724 454708
rect 134300 454668 143724 454696
rect 134300 454656 134306 454668
rect 143718 454656 143724 454668
rect 143776 454656 143782 454708
rect 46842 453976 46848 454028
rect 46900 454016 46906 454028
rect 54846 454016 54852 454028
rect 46900 453988 54852 454016
rect 46900 453976 46906 453988
rect 54846 453976 54852 453988
rect 54904 454016 54910 454028
rect 67634 454016 67640 454028
rect 54904 453988 67640 454016
rect 54904 453976 54910 453988
rect 67634 453976 67640 453988
rect 67692 453976 67698 454028
rect 54478 453296 54484 453348
rect 54536 453336 54542 453348
rect 55030 453336 55036 453348
rect 54536 453308 55036 453336
rect 54536 453296 54542 453308
rect 55030 453296 55036 453308
rect 55088 453336 55094 453348
rect 67634 453336 67640 453348
rect 55088 453308 67640 453336
rect 55088 453296 55094 453308
rect 67634 453296 67640 453308
rect 67692 453296 67698 453348
rect 102870 453296 102876 453348
rect 102928 453336 102934 453348
rect 125594 453336 125600 453348
rect 102928 453308 125600 453336
rect 102928 453296 102934 453308
rect 125594 453296 125600 453308
rect 125652 453296 125658 453348
rect 102134 453228 102140 453280
rect 102192 453268 102198 453280
rect 106182 453268 106188 453280
rect 102192 453240 106188 453268
rect 102192 453228 102198 453240
rect 106182 453228 106188 453240
rect 106240 453228 106246 453280
rect 102134 452548 102140 452600
rect 102192 452588 102198 452600
rect 116210 452588 116216 452600
rect 102192 452560 116216 452588
rect 102192 452548 102198 452560
rect 116210 452548 116216 452560
rect 116268 452588 116274 452600
rect 124858 452588 124864 452600
rect 116268 452560 124864 452588
rect 116268 452548 116274 452560
rect 124858 452548 124864 452560
rect 124916 452548 124922 452600
rect 103606 451868 103612 451920
rect 103664 451908 103670 451920
rect 134150 451908 134156 451920
rect 103664 451880 134156 451908
rect 103664 451868 103670 451880
rect 134150 451868 134156 451880
rect 134208 451908 134214 451920
rect 147766 451908 147772 451920
rect 134208 451880 147772 451908
rect 134208 451868 134214 451880
rect 147766 451868 147772 451880
rect 147824 451868 147830 451920
rect 103698 451664 103704 451716
rect 103756 451704 103762 451716
rect 107838 451704 107844 451716
rect 103756 451676 107844 451704
rect 103756 451664 103762 451676
rect 107838 451664 107844 451676
rect 107896 451664 107902 451716
rect 69198 451296 69204 451308
rect 62776 451268 69204 451296
rect 62776 451240 62804 451268
rect 69198 451256 69204 451268
rect 69256 451256 69262 451308
rect 46750 451188 46756 451240
rect 46808 451228 46814 451240
rect 62758 451228 62764 451240
rect 46808 451200 62764 451228
rect 46808 451188 46814 451200
rect 62758 451188 62764 451200
rect 62816 451188 62822 451240
rect 61378 449936 61384 449948
rect 60752 449908 61384 449936
rect 41138 449828 41144 449880
rect 41196 449868 41202 449880
rect 60752 449868 60780 449908
rect 61378 449896 61384 449908
rect 61436 449936 61442 449948
rect 67634 449936 67640 449948
rect 61436 449908 67640 449936
rect 61436 449896 61442 449908
rect 67634 449896 67640 449908
rect 67692 449896 67698 449948
rect 106918 449896 106924 449948
rect 106976 449936 106982 449948
rect 140774 449936 140780 449948
rect 106976 449908 140780 449936
rect 106976 449896 106982 449908
rect 140774 449896 140780 449908
rect 140832 449896 140838 449948
rect 41196 449840 60780 449868
rect 41196 449828 41202 449840
rect 102134 449828 102140 449880
rect 102192 449868 102198 449880
rect 106936 449868 106964 449896
rect 102192 449840 106964 449868
rect 102192 449828 102198 449840
rect 56410 449148 56416 449200
rect 56468 449188 56474 449200
rect 67634 449188 67640 449200
rect 56468 449160 67640 449188
rect 56468 449148 56474 449160
rect 67634 449148 67640 449160
rect 67692 449148 67698 449200
rect 106182 449148 106188 449200
rect 106240 449188 106246 449200
rect 142430 449188 142436 449200
rect 106240 449160 142436 449188
rect 106240 449148 106246 449160
rect 142430 449148 142436 449160
rect 142488 449188 142494 449200
rect 143810 449188 143816 449200
rect 142488 449160 143816 449188
rect 142488 449148 142494 449160
rect 143810 449148 143816 449160
rect 143868 449148 143874 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 50338 448576 50344 448588
rect 3200 448548 50344 448576
rect 3200 448536 3206 448548
rect 50338 448536 50344 448548
rect 50396 448536 50402 448588
rect 55858 448536 55864 448588
rect 55916 448576 55922 448588
rect 56410 448576 56416 448588
rect 55916 448548 56416 448576
rect 55916 448536 55922 448548
rect 56410 448536 56416 448548
rect 56468 448536 56474 448588
rect 102226 448468 102232 448520
rect 102284 448508 102290 448520
rect 107470 448508 107476 448520
rect 102284 448480 107476 448508
rect 102284 448468 102290 448480
rect 107470 448468 107476 448480
rect 107528 448468 107534 448520
rect 102134 448400 102140 448452
rect 102192 448440 102198 448452
rect 106182 448440 106188 448452
rect 102192 448412 106188 448440
rect 102192 448400 102198 448412
rect 106182 448400 106188 448412
rect 106240 448400 106246 448452
rect 107470 448060 107476 448112
rect 107528 448100 107534 448112
rect 113450 448100 113456 448112
rect 107528 448072 113456 448100
rect 107528 448060 107534 448072
rect 113450 448060 113456 448072
rect 113508 448060 113514 448112
rect 61654 447176 61660 447228
rect 61712 447216 61718 447228
rect 66254 447216 66260 447228
rect 61712 447188 66260 447216
rect 61712 447176 61718 447188
rect 66254 447176 66260 447188
rect 66312 447216 66318 447228
rect 67634 447216 67640 447228
rect 66312 447188 67640 447216
rect 66312 447176 66318 447188
rect 67634 447176 67640 447188
rect 67692 447176 67698 447228
rect 64782 447108 64788 447160
rect 64840 447148 64846 447160
rect 66162 447148 66168 447160
rect 64840 447120 66168 447148
rect 64840 447108 64846 447120
rect 66162 447108 66168 447120
rect 66220 447148 66226 447160
rect 67726 447148 67732 447160
rect 66220 447120 67732 447148
rect 66220 447108 66226 447120
rect 67726 447108 67732 447120
rect 67784 447108 67790 447160
rect 33042 446360 33048 446412
rect 33100 446400 33106 446412
rect 67634 446400 67640 446412
rect 33100 446372 67640 446400
rect 33100 446360 33106 446372
rect 67634 446360 67640 446372
rect 67692 446360 67698 446412
rect 104158 445816 104164 445868
rect 104216 445856 104222 445868
rect 108390 445856 108396 445868
rect 104216 445828 108396 445856
rect 104216 445816 104222 445828
rect 108390 445816 108396 445828
rect 108448 445816 108454 445868
rect 60550 445748 60556 445800
rect 60608 445788 60614 445800
rect 64598 445788 64604 445800
rect 60608 445760 64604 445788
rect 60608 445748 60614 445760
rect 64598 445748 64604 445760
rect 64656 445788 64662 445800
rect 67726 445788 67732 445800
rect 64656 445760 67732 445788
rect 64656 445748 64662 445760
rect 67726 445748 67732 445760
rect 67784 445748 67790 445800
rect 101950 445748 101956 445800
rect 102008 445788 102014 445800
rect 138198 445788 138204 445800
rect 102008 445760 138204 445788
rect 102008 445748 102014 445760
rect 138198 445748 138204 445760
rect 138256 445748 138262 445800
rect 103146 445068 103152 445120
rect 103204 445108 103210 445120
rect 104158 445108 104164 445120
rect 103204 445080 104164 445108
rect 103204 445068 103210 445080
rect 104158 445068 104164 445080
rect 104216 445068 104222 445120
rect 102594 445000 102600 445052
rect 102652 445040 102658 445052
rect 128538 445040 128544 445052
rect 102652 445012 128544 445040
rect 102652 445000 102658 445012
rect 128538 445000 128544 445012
rect 128596 445040 128602 445052
rect 142154 445040 142160 445052
rect 128596 445012 142160 445040
rect 128596 445000 128602 445012
rect 142154 445000 142160 445012
rect 142212 445000 142218 445052
rect 99466 444388 99472 444440
rect 99524 444428 99530 444440
rect 100754 444428 100760 444440
rect 99524 444400 100760 444428
rect 99524 444388 99530 444400
rect 100754 444388 100760 444400
rect 100812 444388 100818 444440
rect 45462 443640 45468 443692
rect 45520 443680 45526 443692
rect 67634 443680 67640 443692
rect 45520 443652 67640 443680
rect 45520 443640 45526 443652
rect 67634 443640 67640 443652
rect 67692 443640 67698 443692
rect 61930 442892 61936 442944
rect 61988 442932 61994 442944
rect 63402 442932 63408 442944
rect 61988 442904 63408 442932
rect 61988 442892 61994 442904
rect 63402 442892 63408 442904
rect 63460 442932 63466 442944
rect 67634 442932 67640 442944
rect 63460 442904 67640 442932
rect 63460 442892 63466 442904
rect 67634 442892 67640 442904
rect 67692 442892 67698 442944
rect 38562 442212 38568 442264
rect 38620 442252 38626 442264
rect 67634 442252 67640 442264
rect 38620 442224 67640 442252
rect 38620 442212 38626 442224
rect 67634 442212 67640 442224
rect 67692 442212 67698 442264
rect 102686 441668 102692 441720
rect 102744 441708 102750 441720
rect 112530 441708 112536 441720
rect 102744 441680 112536 441708
rect 102744 441668 102750 441680
rect 112530 441668 112536 441680
rect 112588 441668 112594 441720
rect 103146 441600 103152 441652
rect 103204 441640 103210 441652
rect 132862 441640 132868 441652
rect 103204 441612 132868 441640
rect 103204 441600 103210 441612
rect 132862 441600 132868 441612
rect 132920 441600 132926 441652
rect 60642 441532 60648 441584
rect 60700 441572 60706 441584
rect 67634 441572 67640 441584
rect 60700 441544 67640 441572
rect 60700 441532 60706 441544
rect 67634 441532 67640 441544
rect 67692 441532 67698 441584
rect 62022 440988 62028 441040
rect 62080 441028 62086 441040
rect 67634 441028 67640 441040
rect 62080 441000 67640 441028
rect 62080 440988 62086 441000
rect 67634 440988 67640 441000
rect 67692 440988 67698 441040
rect 52086 440920 52092 440972
rect 52144 440960 52150 440972
rect 112070 440960 112076 440972
rect 52144 440932 69796 440960
rect 52144 440920 52150 440932
rect 45278 440852 45284 440904
rect 45336 440892 45342 440904
rect 45336 440864 64874 440892
rect 45336 440852 45342 440864
rect 64846 440688 64874 440864
rect 69768 440756 69796 440932
rect 92400 440932 112076 440960
rect 69768 440728 72372 440756
rect 72344 440700 72372 440728
rect 92400 440700 92428 440932
rect 112070 440920 112076 440932
rect 112128 440920 112134 440972
rect 117498 440892 117504 440904
rect 99346 440864 117504 440892
rect 72142 440688 72148 440700
rect 64846 440660 72148 440688
rect 72142 440648 72148 440660
rect 72200 440648 72206 440700
rect 72326 440648 72332 440700
rect 72384 440648 72390 440700
rect 92382 440648 92388 440700
rect 92440 440648 92446 440700
rect 94130 440648 94136 440700
rect 94188 440688 94194 440700
rect 99346 440688 99374 440864
rect 117498 440852 117504 440864
rect 117556 440852 117562 440904
rect 94188 440660 99374 440688
rect 94188 440648 94194 440660
rect 103146 440308 103152 440360
rect 103204 440348 103210 440360
rect 127066 440348 127072 440360
rect 103204 440320 127072 440348
rect 103204 440308 103210 440320
rect 127066 440308 127072 440320
rect 127124 440348 127130 440360
rect 132678 440348 132684 440360
rect 127124 440320 132684 440348
rect 127124 440308 127130 440320
rect 132678 440308 132684 440320
rect 132736 440308 132742 440360
rect 102134 440240 102140 440292
rect 102192 440280 102198 440292
rect 133874 440280 133880 440292
rect 102192 440252 133880 440280
rect 102192 440240 102198 440252
rect 133874 440240 133880 440252
rect 133932 440240 133938 440292
rect 67266 439560 67272 439612
rect 67324 439600 67330 439612
rect 75178 439600 75184 439612
rect 67324 439572 75184 439600
rect 67324 439560 67330 439572
rect 75178 439560 75184 439572
rect 75236 439560 75242 439612
rect 89806 439560 89812 439612
rect 89864 439600 89870 439612
rect 113542 439600 113548 439612
rect 89864 439572 113548 439600
rect 89864 439560 89870 439572
rect 113542 439560 113548 439572
rect 113600 439560 113606 439612
rect 53650 439492 53656 439544
rect 53708 439532 53714 439544
rect 83458 439532 83464 439544
rect 53708 439504 83464 439532
rect 53708 439492 53714 439504
rect 83458 439492 83464 439504
rect 83516 439532 83522 439544
rect 85758 439532 85764 439544
rect 83516 439504 85764 439532
rect 83516 439492 83522 439504
rect 85758 439492 85764 439504
rect 85816 439492 85822 439544
rect 96522 439492 96528 439544
rect 96580 439532 96586 439544
rect 120258 439532 120264 439544
rect 96580 439504 120264 439532
rect 96580 439492 96586 439504
rect 120258 439492 120264 439504
rect 120316 439492 120322 439544
rect 56134 439016 56140 439068
rect 56192 439056 56198 439068
rect 59262 439056 59268 439068
rect 56192 439028 59268 439056
rect 56192 439016 56198 439028
rect 59262 439016 59268 439028
rect 59320 439056 59326 439068
rect 90910 439056 90916 439068
rect 59320 439028 90916 439056
rect 59320 439016 59326 439028
rect 90910 439016 90916 439028
rect 90968 439016 90974 439068
rect 88702 438948 88708 439000
rect 88760 438988 88766 439000
rect 123478 438988 123484 439000
rect 88760 438960 123484 438988
rect 88760 438948 88766 438960
rect 123478 438948 123484 438960
rect 123536 438988 123542 439000
rect 123754 438988 123760 439000
rect 123536 438960 123760 438988
rect 123536 438948 123542 438960
rect 123754 438948 123760 438960
rect 123812 438948 123818 439000
rect 25498 438880 25504 438932
rect 25556 438920 25562 438932
rect 96430 438920 96436 438932
rect 25556 438892 96436 438920
rect 25556 438880 25562 438892
rect 96430 438880 96436 438892
rect 96488 438880 96494 438932
rect 122926 438920 122932 438932
rect 122806 438892 122932 438920
rect 4798 438812 4804 438864
rect 4856 438852 4862 438864
rect 50890 438852 50896 438864
rect 4856 438824 50896 438852
rect 4856 438812 4862 438824
rect 50890 438812 50896 438824
rect 50948 438812 50954 438864
rect 89990 438812 89996 438864
rect 90048 438852 90054 438864
rect 95878 438852 95884 438864
rect 90048 438824 95884 438852
rect 90048 438812 90054 438824
rect 95878 438812 95884 438824
rect 95936 438852 95942 438864
rect 96522 438852 96528 438864
rect 95936 438824 96528 438852
rect 95936 438812 95942 438824
rect 96522 438812 96528 438824
rect 96580 438812 96586 438864
rect 99650 438812 99656 438864
rect 99708 438852 99714 438864
rect 122806 438852 122834 438892
rect 122926 438880 122932 438892
rect 122984 438920 122990 438932
rect 129918 438920 129924 438932
rect 122984 438892 129924 438920
rect 122984 438880 122990 438892
rect 129918 438880 129924 438892
rect 129976 438880 129982 438932
rect 99708 438824 122834 438852
rect 99708 438812 99714 438824
rect 46658 438744 46664 438796
rect 46716 438784 46722 438796
rect 78766 438784 78772 438796
rect 46716 438756 78772 438784
rect 46716 438744 46722 438756
rect 78766 438744 78772 438756
rect 78824 438744 78830 438796
rect 96430 438744 96436 438796
rect 96488 438784 96494 438796
rect 121638 438784 121644 438796
rect 96488 438756 121644 438784
rect 96488 438744 96494 438756
rect 121638 438744 121644 438756
rect 121696 438744 121702 438796
rect 52178 438676 52184 438728
rect 52236 438716 52242 438728
rect 53742 438716 53748 438728
rect 52236 438688 53748 438716
rect 52236 438676 52242 438688
rect 53742 438676 53748 438688
rect 53800 438716 53806 438728
rect 82906 438716 82912 438728
rect 53800 438688 82912 438716
rect 53800 438676 53806 438688
rect 82906 438676 82912 438688
rect 82964 438676 82970 438728
rect 99006 438676 99012 438728
rect 99064 438716 99070 438728
rect 120350 438716 120356 438728
rect 99064 438688 120356 438716
rect 99064 438676 99070 438688
rect 120350 438676 120356 438688
rect 120408 438716 120414 438728
rect 120902 438716 120908 438728
rect 120408 438688 120908 438716
rect 120408 438676 120414 438688
rect 120902 438676 120908 438688
rect 120960 438676 120966 438728
rect 87598 438608 87604 438660
rect 87656 438648 87662 438660
rect 105538 438648 105544 438660
rect 87656 438620 105544 438648
rect 87656 438608 87662 438620
rect 105538 438608 105544 438620
rect 105596 438608 105602 438660
rect 97074 438540 97080 438592
rect 97132 438580 97138 438592
rect 113358 438580 113364 438592
rect 97132 438552 113364 438580
rect 97132 438540 97138 438552
rect 113358 438540 113364 438552
rect 113416 438580 113422 438592
rect 114462 438580 114468 438592
rect 113416 438552 114468 438580
rect 113416 438540 113422 438552
rect 114462 438540 114468 438552
rect 114520 438540 114526 438592
rect 50338 438472 50344 438524
rect 50396 438512 50402 438524
rect 99466 438512 99472 438524
rect 50396 438484 99472 438512
rect 50396 438472 50402 438484
rect 99466 438472 99472 438484
rect 99524 438472 99530 438524
rect 53098 438268 53104 438320
rect 53156 438308 53162 438320
rect 73890 438308 73896 438320
rect 53156 438280 73896 438308
rect 53156 438268 53162 438280
rect 73890 438268 73896 438280
rect 73948 438268 73954 438320
rect 88058 438268 88064 438320
rect 88116 438308 88122 438320
rect 88978 438308 88984 438320
rect 88116 438280 88984 438308
rect 88116 438268 88122 438280
rect 88978 438268 88984 438280
rect 89036 438268 89042 438320
rect 121638 438268 121644 438320
rect 121696 438308 121702 438320
rect 125778 438308 125784 438320
rect 121696 438280 125784 438308
rect 121696 438268 121702 438280
rect 125778 438268 125784 438280
rect 125836 438268 125842 438320
rect 44266 438200 44272 438252
rect 44324 438240 44330 438252
rect 71314 438240 71320 438252
rect 44324 438212 71320 438240
rect 44324 438200 44330 438212
rect 71314 438200 71320 438212
rect 71372 438200 71378 438252
rect 83550 438240 83556 438252
rect 74506 438212 83556 438240
rect 50890 438132 50896 438184
rect 50948 438172 50954 438184
rect 52086 438172 52092 438184
rect 50948 438144 52092 438172
rect 50948 438132 50954 438144
rect 52086 438132 52092 438144
rect 52144 438172 52150 438184
rect 74506 438172 74534 438212
rect 83550 438200 83556 438212
rect 83608 438200 83614 438252
rect 92566 438200 92572 438252
rect 92624 438240 92630 438252
rect 97902 438240 97908 438252
rect 92624 438212 97908 438240
rect 92624 438200 92630 438212
rect 97902 438200 97908 438212
rect 97960 438240 97966 438252
rect 101398 438240 101404 438252
rect 97960 438212 101404 438240
rect 97960 438200 97966 438212
rect 101398 438200 101404 438212
rect 101456 438200 101462 438252
rect 120902 438200 120908 438252
rect 120960 438240 120966 438252
rect 129918 438240 129924 438252
rect 120960 438212 129924 438240
rect 120960 438200 120966 438212
rect 129918 438200 129924 438212
rect 129976 438200 129982 438252
rect 52144 438144 74534 438172
rect 52144 438132 52150 438144
rect 75454 438132 75460 438184
rect 75512 438172 75518 438184
rect 82262 438172 82268 438184
rect 75512 438144 82268 438172
rect 75512 438132 75518 438144
rect 82262 438132 82268 438144
rect 82320 438132 82326 438184
rect 84838 438132 84844 438184
rect 84896 438172 84902 438184
rect 97718 438172 97724 438184
rect 84896 438144 97724 438172
rect 84896 438132 84902 438144
rect 97718 438132 97724 438144
rect 97776 438132 97782 438184
rect 114462 438132 114468 438184
rect 114520 438172 114526 438184
rect 135254 438172 135260 438184
rect 114520 438144 135260 438172
rect 114520 438132 114526 438144
rect 135254 438132 135260 438144
rect 135312 438132 135318 438184
rect 78766 437860 78772 437912
rect 78824 437900 78830 437912
rect 79686 437900 79692 437912
rect 78824 437872 79692 437900
rect 78824 437860 78830 437872
rect 79686 437860 79692 437872
rect 79744 437860 79750 437912
rect 81618 437452 81624 437504
rect 81676 437492 81682 437504
rect 82814 437492 82820 437504
rect 81676 437464 82820 437492
rect 81676 437452 81682 437464
rect 82814 437452 82820 437464
rect 82872 437452 82878 437504
rect 38470 437384 38476 437436
rect 38528 437424 38534 437436
rect 44266 437424 44272 437436
rect 38528 437396 44272 437424
rect 38528 437384 38534 437396
rect 44266 437384 44272 437396
rect 44324 437424 44330 437436
rect 44818 437424 44824 437436
rect 44324 437396 44824 437424
rect 44324 437384 44330 437396
rect 44818 437384 44824 437396
rect 44876 437384 44882 437436
rect 52270 437384 52276 437436
rect 52328 437424 52334 437436
rect 86218 437424 86224 437436
rect 52328 437396 86224 437424
rect 52328 437384 52334 437396
rect 86218 437384 86224 437396
rect 86276 437424 86282 437436
rect 86770 437424 86776 437436
rect 86276 437396 86776 437424
rect 86276 437384 86282 437396
rect 86770 437384 86776 437396
rect 86828 437384 86834 437436
rect 94498 437384 94504 437436
rect 94556 437424 94562 437436
rect 128354 437424 128360 437436
rect 94556 437396 128360 437424
rect 94556 437384 94562 437396
rect 128354 437384 128360 437396
rect 128412 437384 128418 437436
rect 49418 437316 49424 437368
rect 49476 437356 49482 437368
rect 81618 437356 81624 437368
rect 49476 437328 81624 437356
rect 49476 437316 49482 437328
rect 81618 437316 81624 437328
rect 81676 437316 81682 437368
rect 95142 437316 95148 437368
rect 95200 437356 95206 437368
rect 118694 437356 118700 437368
rect 95200 437328 118700 437356
rect 95200 437316 95206 437328
rect 118694 437316 118700 437328
rect 118752 437316 118758 437368
rect 39666 437248 39672 437300
rect 39724 437288 39730 437300
rect 71958 437288 71964 437300
rect 39724 437260 71964 437288
rect 39724 437248 39730 437260
rect 71958 437248 71964 437260
rect 72016 437248 72022 437300
rect 72142 437248 72148 437300
rect 72200 437288 72206 437300
rect 77294 437288 77300 437300
rect 72200 437260 77300 437288
rect 72200 437248 72206 437260
rect 77294 437248 77300 437260
rect 77352 437288 77358 437300
rect 77754 437288 77760 437300
rect 77352 437260 77760 437288
rect 77352 437248 77358 437260
rect 77754 437248 77760 437260
rect 77812 437248 77818 437300
rect 41322 437180 41328 437232
rect 41380 437220 41386 437232
rect 53098 437220 53104 437232
rect 41380 437192 53104 437220
rect 41380 437180 41386 437192
rect 53098 437180 53104 437192
rect 53156 437180 53162 437232
rect 58986 437180 58992 437232
rect 59044 437220 59050 437232
rect 78858 437220 78864 437232
rect 59044 437192 78864 437220
rect 59044 437180 59050 437192
rect 78858 437180 78864 437192
rect 78916 437220 78922 437232
rect 79042 437220 79048 437232
rect 78916 437192 79048 437220
rect 78916 437180 78922 437192
rect 79042 437180 79048 437192
rect 79100 437180 79106 437232
rect 65610 436704 65616 436756
rect 65668 436744 65674 436756
rect 76558 436744 76564 436756
rect 65668 436716 76564 436744
rect 65668 436704 65674 436716
rect 76558 436704 76564 436716
rect 76616 436704 76622 436756
rect 97718 436704 97724 436756
rect 97776 436744 97782 436756
rect 107378 436744 107384 436756
rect 97776 436716 107384 436744
rect 97776 436704 97782 436716
rect 107378 436704 107384 436716
rect 107436 436744 107442 436756
rect 108482 436744 108488 436756
rect 107436 436716 108488 436744
rect 107436 436704 107442 436716
rect 108482 436704 108488 436716
rect 108540 436704 108546 436756
rect 57514 436024 57520 436076
rect 57572 436064 57578 436076
rect 91738 436064 91744 436076
rect 57572 436036 91744 436064
rect 57572 436024 57578 436036
rect 91738 436024 91744 436036
rect 91796 436024 91802 436076
rect 45370 435956 45376 436008
rect 45428 435996 45434 436008
rect 74626 435996 74632 436008
rect 45428 435968 74632 435996
rect 45428 435956 45434 435968
rect 74626 435956 74632 435968
rect 74684 435996 74690 436008
rect 75822 435996 75828 436008
rect 74684 435968 75828 435996
rect 74684 435956 74690 435968
rect 75822 435956 75828 435968
rect 75880 435956 75886 436008
rect 42518 435412 42524 435464
rect 42576 435452 42582 435464
rect 44082 435452 44088 435464
rect 42576 435424 44088 435452
rect 42576 435412 42582 435424
rect 44082 435412 44088 435424
rect 44140 435452 44146 435464
rect 77110 435452 77116 435464
rect 44140 435424 77116 435452
rect 44140 435412 44146 435424
rect 77110 435412 77116 435424
rect 77168 435412 77174 435464
rect 40678 435344 40684 435396
rect 40736 435384 40742 435396
rect 73246 435384 73252 435396
rect 40736 435356 73252 435384
rect 40736 435344 40742 435356
rect 73246 435344 73252 435356
rect 73304 435344 73310 435396
rect 39942 434664 39948 434716
rect 40000 434704 40006 434716
rect 40678 434704 40684 434716
rect 40000 434676 40684 434704
rect 40000 434664 40006 434676
rect 40678 434664 40684 434676
rect 40736 434664 40742 434716
rect 51994 434664 52000 434716
rect 52052 434704 52058 434716
rect 69014 434704 69020 434716
rect 52052 434676 69020 434704
rect 52052 434664 52058 434676
rect 69014 434664 69020 434676
rect 69072 434664 69078 434716
rect 78582 434664 78588 434716
rect 78640 434704 78646 434716
rect 82906 434704 82912 434716
rect 78640 434676 82912 434704
rect 78640 434664 78646 434676
rect 82906 434664 82912 434676
rect 82964 434664 82970 434716
rect 38470 433236 38476 433288
rect 38528 433276 38534 433288
rect 41046 433276 41052 433288
rect 38528 433248 41052 433276
rect 38528 433236 38534 433248
rect 41046 433236 41052 433248
rect 41104 433276 41110 433288
rect 70670 433276 70676 433288
rect 41104 433248 70676 433276
rect 41104 433236 41110 433248
rect 70670 433236 70676 433248
rect 70728 433236 70734 433288
rect 55122 433168 55128 433220
rect 55180 433208 55186 433220
rect 76466 433208 76472 433220
rect 55180 433180 76472 433208
rect 55180 433168 55186 433180
rect 76466 433168 76472 433180
rect 76524 433168 76530 433220
rect 82906 431876 82912 431928
rect 82964 431916 82970 431928
rect 579798 431916 579804 431928
rect 82964 431888 579804 431916
rect 82964 431876 82970 431888
rect 579798 431876 579804 431888
rect 579856 431876 579862 431928
rect 101490 431808 101496 431860
rect 101548 431848 101554 431860
rect 140866 431848 140872 431860
rect 101548 431820 140872 431848
rect 101548 431808 101554 431820
rect 140866 431808 140872 431820
rect 140924 431808 140930 431860
rect 140866 431196 140872 431248
rect 140924 431236 140930 431248
rect 150710 431236 150716 431248
rect 140924 431208 150716 431236
rect 140924 431196 140930 431208
rect 150710 431196 150716 431208
rect 150768 431196 150774 431248
rect 3418 429836 3424 429888
rect 3476 429876 3482 429888
rect 101490 429876 101496 429888
rect 3476 429848 101496 429876
rect 3476 429836 3482 429848
rect 101490 429836 101496 429848
rect 101548 429836 101554 429888
rect 69198 428408 69204 428460
rect 69256 428448 69262 428460
rect 579614 428448 579620 428460
rect 69256 428420 579620 428448
rect 69256 428408 69262 428420
rect 579614 428408 579620 428420
rect 579672 428408 579678 428460
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 3568 422300 115934 422328
rect 3568 422288 3574 422300
rect 115906 422260 115934 422300
rect 118786 422260 118792 422272
rect 115906 422232 118792 422260
rect 118786 422220 118792 422232
rect 118844 422220 118850 422272
rect 118786 420928 118792 420980
rect 118844 420968 118850 420980
rect 119338 420968 119344 420980
rect 118844 420940 119344 420968
rect 118844 420928 118850 420940
rect 119338 420928 119344 420940
rect 119396 420928 119402 420980
rect 525058 418752 525064 418804
rect 525116 418792 525122 418804
rect 579614 418792 579620 418804
rect 525116 418764 579620 418792
rect 525116 418752 525122 418764
rect 579614 418752 579620 418764
rect 579672 418792 579678 418804
rect 579982 418792 579988 418804
rect 579672 418764 579988 418792
rect 579672 418752 579678 418764
rect 579982 418752 579988 418764
rect 580040 418752 580046 418804
rect 87690 404336 87696 404388
rect 87748 404376 87754 404388
rect 579614 404376 579620 404388
rect 87748 404348 579620 404376
rect 87748 404336 87754 404348
rect 579614 404336 579620 404348
rect 579672 404336 579678 404388
rect 104250 403656 104256 403708
rect 104308 403696 104314 403708
rect 128630 403696 128636 403708
rect 104308 403668 128636 403696
rect 104308 403656 104314 403668
rect 128630 403656 128636 403668
rect 128688 403656 128694 403708
rect 96614 403588 96620 403640
rect 96672 403628 96678 403640
rect 127250 403628 127256 403640
rect 96672 403600 127256 403628
rect 96672 403588 96678 403600
rect 127250 403588 127256 403600
rect 127308 403588 127314 403640
rect 61838 402976 61844 403028
rect 61896 403016 61902 403028
rect 289078 403016 289084 403028
rect 61896 402988 289084 403016
rect 61896 402976 61902 402988
rect 289078 402976 289084 402988
rect 289136 402976 289142 403028
rect 93762 402228 93768 402280
rect 93820 402268 93826 402280
rect 130010 402268 130016 402280
rect 93820 402240 130016 402268
rect 93820 402228 93826 402240
rect 130010 402228 130016 402240
rect 130068 402228 130074 402280
rect 70394 401616 70400 401668
rect 70452 401656 70458 401668
rect 71038 401656 71044 401668
rect 70452 401628 71044 401656
rect 70452 401616 70458 401628
rect 71038 401616 71044 401628
rect 71096 401656 71102 401668
rect 358814 401656 358820 401668
rect 71096 401628 358820 401656
rect 71096 401616 71102 401628
rect 358814 401616 358820 401628
rect 358872 401616 358878 401668
rect 104158 401004 104164 401056
rect 104216 401044 104222 401056
rect 132770 401044 132776 401056
rect 104216 401016 132776 401044
rect 104216 401004 104222 401016
rect 132770 401004 132776 401016
rect 132828 401004 132834 401056
rect 86218 400936 86224 400988
rect 86276 400976 86282 400988
rect 123110 400976 123116 400988
rect 86276 400948 123116 400976
rect 86276 400936 86282 400948
rect 123110 400936 123116 400948
rect 123168 400936 123174 400988
rect 93670 400868 93676 400920
rect 93728 400908 93734 400920
rect 131298 400908 131304 400920
rect 93728 400880 131304 400908
rect 93728 400868 93734 400880
rect 131298 400868 131304 400880
rect 131356 400868 131362 400920
rect 69106 400228 69112 400240
rect 62132 400200 69112 400228
rect 50798 400120 50804 400172
rect 50856 400160 50862 400172
rect 62132 400160 62160 400200
rect 69106 400188 69112 400200
rect 69164 400228 69170 400240
rect 357434 400228 357440 400240
rect 69164 400200 357440 400228
rect 69164 400188 69170 400200
rect 357434 400188 357440 400200
rect 357492 400188 357498 400240
rect 50856 400132 62160 400160
rect 50856 400120 50862 400132
rect 107562 399508 107568 399560
rect 107620 399548 107626 399560
rect 117498 399548 117504 399560
rect 107620 399520 117504 399548
rect 107620 399508 107626 399520
rect 117498 399508 117504 399520
rect 117556 399508 117562 399560
rect 91738 399440 91744 399492
rect 91796 399480 91802 399492
rect 124306 399480 124312 399492
rect 91796 399452 124312 399480
rect 91796 399440 91802 399452
rect 124306 399440 124312 399452
rect 124364 399440 124370 399492
rect 94130 398896 94136 398948
rect 94188 398936 94194 398948
rect 115106 398936 115112 398948
rect 94188 398908 115112 398936
rect 94188 398896 94194 398908
rect 115106 398896 115112 398908
rect 115164 398936 115170 398948
rect 115164 398908 122834 398936
rect 115164 398896 115170 398908
rect 50982 398828 50988 398880
rect 51040 398868 51046 398880
rect 107010 398868 107016 398880
rect 51040 398840 107016 398868
rect 51040 398828 51046 398840
rect 107010 398828 107016 398840
rect 107068 398868 107074 398880
rect 114830 398868 114836 398880
rect 107068 398840 114836 398868
rect 107068 398828 107074 398840
rect 114830 398828 114836 398840
rect 114888 398828 114894 398880
rect 122806 398868 122834 398908
rect 160738 398868 160744 398880
rect 122806 398840 160744 398868
rect 160738 398828 160744 398840
rect 160796 398828 160802 398880
rect 108390 398216 108396 398268
rect 108448 398256 108454 398268
rect 136818 398256 136824 398268
rect 108448 398228 136824 398256
rect 108448 398216 108454 398228
rect 136818 398216 136824 398228
rect 136876 398216 136882 398268
rect 56226 398148 56232 398200
rect 56284 398188 56290 398200
rect 71038 398188 71044 398200
rect 56284 398160 71044 398188
rect 56284 398148 56290 398160
rect 71038 398148 71044 398160
rect 71096 398148 71102 398200
rect 108298 398148 108304 398200
rect 108356 398188 108362 398200
rect 140866 398188 140872 398200
rect 108356 398160 140872 398188
rect 108356 398148 108362 398160
rect 140866 398148 140872 398160
rect 140924 398148 140930 398200
rect 3142 398080 3148 398132
rect 3200 398120 3206 398132
rect 116026 398120 116032 398132
rect 3200 398092 116032 398120
rect 3200 398080 3206 398092
rect 116026 398080 116032 398092
rect 116084 398080 116090 398132
rect 98638 397536 98644 397588
rect 98696 397576 98702 397588
rect 188338 397576 188344 397588
rect 98696 397548 188344 397576
rect 98696 397536 98702 397548
rect 188338 397536 188344 397548
rect 188396 397536 188402 397588
rect 67358 397468 67364 397520
rect 67416 397508 67422 397520
rect 202138 397508 202144 397520
rect 67416 397480 202144 397508
rect 67416 397468 67422 397480
rect 202138 397468 202144 397480
rect 202196 397468 202202 397520
rect 95878 396856 95884 396908
rect 95936 396896 95942 396908
rect 120718 396896 120724 396908
rect 95936 396868 120724 396896
rect 95936 396856 95942 396868
rect 120718 396856 120724 396868
rect 120776 396856 120782 396908
rect 69658 396788 69664 396840
rect 69716 396828 69722 396840
rect 94498 396828 94504 396840
rect 69716 396800 94504 396828
rect 69716 396788 69722 396800
rect 94498 396788 94504 396800
rect 94556 396788 94562 396840
rect 101122 396788 101128 396840
rect 101180 396828 101186 396840
rect 131206 396828 131212 396840
rect 101180 396800 131212 396828
rect 101180 396788 101186 396800
rect 131206 396788 131212 396800
rect 131264 396828 131270 396840
rect 131264 396800 132494 396828
rect 131264 396788 131270 396800
rect 46750 396720 46756 396772
rect 46808 396760 46814 396772
rect 77294 396760 77300 396772
rect 46808 396732 77300 396760
rect 46808 396720 46814 396732
rect 77294 396720 77300 396732
rect 77352 396720 77358 396772
rect 95142 396720 95148 396772
rect 95200 396760 95206 396772
rect 125686 396760 125692 396772
rect 95200 396732 125692 396760
rect 95200 396720 95206 396732
rect 125686 396720 125692 396732
rect 125744 396720 125750 396772
rect 132466 396760 132494 396800
rect 178678 396760 178684 396772
rect 132466 396732 178684 396760
rect 178678 396720 178684 396732
rect 178736 396720 178742 396772
rect 72418 396040 72424 396092
rect 72476 396080 72482 396092
rect 146938 396080 146944 396092
rect 72476 396052 146944 396080
rect 72476 396040 72482 396052
rect 146938 396040 146944 396052
rect 146996 396040 147002 396092
rect 116578 395972 116584 396024
rect 116636 396012 116642 396024
rect 120258 396012 120264 396024
rect 116636 395984 120264 396012
rect 116636 395972 116642 395984
rect 120258 395972 120264 395984
rect 120316 395972 120322 396024
rect 46566 395360 46572 395412
rect 46624 395400 46630 395412
rect 81802 395400 81808 395412
rect 46624 395372 81808 395400
rect 46624 395360 46630 395372
rect 81802 395360 81808 395372
rect 81860 395360 81866 395412
rect 110598 395360 110604 395412
rect 110656 395400 110662 395412
rect 127158 395400 127164 395412
rect 110656 395372 127164 395400
rect 110656 395360 110662 395372
rect 127158 395360 127164 395372
rect 127216 395360 127222 395412
rect 42610 395292 42616 395344
rect 42668 395332 42674 395344
rect 84838 395332 84844 395344
rect 42668 395304 84844 395332
rect 42668 395292 42674 395304
rect 84838 395292 84844 395304
rect 84896 395292 84902 395344
rect 88334 395292 88340 395344
rect 88392 395332 88398 395344
rect 123018 395332 123024 395344
rect 88392 395304 123024 395332
rect 88392 395292 88398 395304
rect 123018 395292 123024 395304
rect 123076 395332 123082 395344
rect 170398 395332 170404 395344
rect 123076 395304 170404 395332
rect 123076 395292 123082 395304
rect 170398 395292 170404 395304
rect 170456 395292 170462 395344
rect 39574 394816 39580 394868
rect 39632 394856 39638 394868
rect 110598 394856 110604 394868
rect 39632 394828 110604 394856
rect 39632 394816 39638 394828
rect 110598 394816 110604 394828
rect 110656 394816 110662 394868
rect 81802 394748 81808 394800
rect 81860 394788 81866 394800
rect 154574 394788 154580 394800
rect 81860 394760 154580 394788
rect 81860 394748 81866 394760
rect 154574 394748 154580 394760
rect 154632 394748 154638 394800
rect 84838 394680 84844 394732
rect 84896 394720 84902 394732
rect 85114 394720 85120 394732
rect 84896 394692 85120 394720
rect 84896 394680 84902 394692
rect 85114 394680 85120 394692
rect 85172 394720 85178 394732
rect 195238 394720 195244 394732
rect 85172 394692 195244 394720
rect 85172 394680 85178 394692
rect 195238 394680 195244 394692
rect 195296 394680 195302 394732
rect 77846 394136 77852 394188
rect 77904 394176 77910 394188
rect 87690 394176 87696 394188
rect 77904 394148 87696 394176
rect 77904 394136 77910 394148
rect 87690 394136 87696 394148
rect 87748 394136 87754 394188
rect 105630 394136 105636 394188
rect 105688 394176 105694 394188
rect 117590 394176 117596 394188
rect 105688 394148 117596 394176
rect 105688 394136 105694 394148
rect 117590 394136 117596 394148
rect 117648 394136 117654 394188
rect 57698 394068 57704 394120
rect 57756 394108 57762 394120
rect 83458 394108 83464 394120
rect 57756 394080 83464 394108
rect 57756 394068 57762 394080
rect 83458 394068 83464 394080
rect 83516 394068 83522 394120
rect 103330 394068 103336 394120
rect 103388 394108 103394 394120
rect 116118 394108 116124 394120
rect 103388 394080 116124 394108
rect 103388 394068 103394 394080
rect 116118 394068 116124 394080
rect 116176 394068 116182 394120
rect 47946 394000 47952 394052
rect 48004 394040 48010 394052
rect 78766 394040 78772 394052
rect 48004 394012 78772 394040
rect 48004 394000 48010 394012
rect 78766 394000 78772 394012
rect 78824 394000 78830 394052
rect 99282 394000 99288 394052
rect 99340 394040 99346 394052
rect 135438 394040 135444 394052
rect 99340 394012 135444 394040
rect 99340 394000 99346 394012
rect 135438 394000 135444 394012
rect 135496 394000 135502 394052
rect 39850 393932 39856 393984
rect 39908 393972 39914 393984
rect 82998 393972 83004 393984
rect 39908 393944 83004 393972
rect 39908 393932 39914 393944
rect 82998 393932 83004 393944
rect 83056 393932 83062 393984
rect 98546 393932 98552 393984
rect 98604 393972 98610 393984
rect 126974 393972 126980 393984
rect 98604 393944 126980 393972
rect 98604 393932 98610 393944
rect 126974 393932 126980 393944
rect 127032 393972 127038 393984
rect 196618 393972 196624 393984
rect 127032 393944 196624 393972
rect 127032 393932 127038 393944
rect 196618 393932 196624 393944
rect 196676 393932 196682 393984
rect 82998 393388 83004 393440
rect 83056 393428 83062 393440
rect 150434 393428 150440 393440
rect 83056 393400 150440 393428
rect 83056 393388 83062 393400
rect 150434 393388 150440 393400
rect 150492 393388 150498 393440
rect 147674 393360 147680 393372
rect 64892 393332 147680 393360
rect 53650 393252 53656 393304
rect 53708 393292 53714 393304
rect 64892 393292 64920 393332
rect 147674 393320 147680 393332
rect 147732 393320 147738 393372
rect 53708 393264 64920 393292
rect 53708 393252 53714 393264
rect 60642 392640 60648 392692
rect 60700 392680 60706 392692
rect 89806 392680 89812 392692
rect 60700 392652 89812 392680
rect 60700 392640 60706 392652
rect 89806 392640 89812 392652
rect 89864 392640 89870 392692
rect 97442 392640 97448 392692
rect 97500 392680 97506 392692
rect 131390 392680 131396 392692
rect 97500 392652 131396 392680
rect 97500 392640 97506 392652
rect 131390 392640 131396 392652
rect 131448 392680 131454 392692
rect 139578 392680 139584 392692
rect 131448 392652 139584 392680
rect 131448 392640 131454 392652
rect 139578 392640 139584 392652
rect 139636 392640 139642 392692
rect 43990 392572 43996 392624
rect 44048 392612 44054 392624
rect 82906 392612 82912 392624
rect 44048 392584 82912 392612
rect 44048 392572 44054 392584
rect 82906 392572 82912 392584
rect 82964 392572 82970 392624
rect 88242 392572 88248 392624
rect 88300 392612 88306 392624
rect 121546 392612 121552 392624
rect 88300 392584 121552 392612
rect 88300 392572 88306 392584
rect 121546 392572 121552 392584
rect 121604 392612 121610 392624
rect 186958 392612 186964 392624
rect 121604 392584 186964 392612
rect 121604 392572 121610 392584
rect 186958 392572 186964 392584
rect 187016 392572 187022 392624
rect 91554 392096 91560 392148
rect 91612 392136 91618 392148
rect 92382 392136 92388 392148
rect 91612 392108 92388 392136
rect 91612 392096 91618 392108
rect 92382 392096 92388 392108
rect 92440 392136 92446 392148
rect 121546 392136 121552 392148
rect 92440 392108 121552 392136
rect 92440 392096 92446 392108
rect 121546 392096 121552 392108
rect 121604 392096 121610 392148
rect 82906 392028 82912 392080
rect 82964 392068 82970 392080
rect 83642 392068 83648 392080
rect 82964 392040 83648 392068
rect 82964 392028 82970 392040
rect 83642 392028 83648 392040
rect 83700 392068 83706 392080
rect 138014 392068 138020 392080
rect 83700 392040 138020 392068
rect 83700 392028 83706 392040
rect 138014 392028 138020 392040
rect 138072 392028 138078 392080
rect 51718 391960 51724 392012
rect 51776 392000 51782 392012
rect 51776 391972 115888 392000
rect 51776 391960 51782 391972
rect 115860 391932 115888 391972
rect 121638 391932 121644 391944
rect 115860 391904 121644 391932
rect 121638 391892 121644 391904
rect 121696 391892 121702 391944
rect 109402 391620 109408 391672
rect 109460 391660 109466 391672
rect 110690 391660 110696 391672
rect 109460 391632 110696 391660
rect 109460 391620 109466 391632
rect 110690 391620 110696 391632
rect 110748 391620 110754 391672
rect 39758 391280 39764 391332
rect 39816 391320 39822 391332
rect 52454 391320 52460 391332
rect 39816 391292 52460 391320
rect 39816 391280 39822 391292
rect 52454 391280 52460 391292
rect 52512 391280 52518 391332
rect 57606 391280 57612 391332
rect 57664 391320 57670 391332
rect 78214 391320 78220 391332
rect 57664 391292 78220 391320
rect 57664 391280 57670 391292
rect 78214 391280 78220 391292
rect 78272 391280 78278 391332
rect 112530 391280 112536 391332
rect 112588 391320 112594 391332
rect 131206 391320 131212 391332
rect 112588 391292 131212 391320
rect 112588 391280 112594 391292
rect 131206 391280 131212 391292
rect 131264 391280 131270 391332
rect 47578 391212 47584 391264
rect 47636 391252 47642 391264
rect 75546 391252 75552 391264
rect 47636 391224 75552 391252
rect 47636 391212 47642 391224
rect 75546 391212 75552 391224
rect 75604 391212 75610 391264
rect 110690 391212 110696 391264
rect 110748 391252 110754 391264
rect 228358 391252 228364 391264
rect 110748 391224 228364 391252
rect 110748 391212 110754 391224
rect 228358 391212 228364 391224
rect 228416 391212 228422 391264
rect 52454 390736 52460 390788
rect 52512 390776 52518 390788
rect 53190 390776 53196 390788
rect 52512 390748 53196 390776
rect 52512 390736 52518 390748
rect 53190 390736 53196 390748
rect 53248 390776 53254 390788
rect 84470 390776 84476 390788
rect 53248 390748 84476 390776
rect 53248 390736 53254 390748
rect 84470 390736 84476 390748
rect 84528 390736 84534 390788
rect 111702 390736 111708 390788
rect 111760 390776 111766 390788
rect 114922 390776 114928 390788
rect 111760 390748 114928 390776
rect 111760 390736 111766 390748
rect 114922 390736 114928 390748
rect 114980 390736 114986 390788
rect 34330 390668 34336 390720
rect 34388 390708 34394 390720
rect 36538 390708 36544 390720
rect 34388 390680 36544 390708
rect 34388 390668 34394 390680
rect 36538 390668 36544 390680
rect 36596 390708 36602 390720
rect 80054 390708 80060 390720
rect 36596 390680 80060 390708
rect 36596 390668 36602 390680
rect 80054 390668 80060 390680
rect 80112 390668 80118 390720
rect 94038 390668 94044 390720
rect 94096 390708 94102 390720
rect 123478 390708 123484 390720
rect 94096 390680 123484 390708
rect 94096 390668 94102 390680
rect 123478 390668 123484 390680
rect 123536 390708 123542 390720
rect 125870 390708 125876 390720
rect 123536 390680 125876 390708
rect 123536 390668 123542 390680
rect 125870 390668 125876 390680
rect 125928 390668 125934 390720
rect 78214 390600 78220 390652
rect 78272 390640 78278 390652
rect 126974 390640 126980 390652
rect 78272 390612 126980 390640
rect 78272 390600 78278 390612
rect 126974 390600 126980 390612
rect 127032 390600 127038 390652
rect 75546 390532 75552 390584
rect 75604 390572 75610 390584
rect 137278 390572 137284 390584
rect 75604 390544 137284 390572
rect 75604 390532 75610 390544
rect 137278 390532 137284 390544
rect 137336 390532 137342 390584
rect 107470 390464 107476 390516
rect 107528 390504 107534 390516
rect 114278 390504 114284 390516
rect 107528 390476 114284 390504
rect 107528 390464 107534 390476
rect 114278 390464 114284 390476
rect 114336 390464 114342 390516
rect 103238 389852 103244 389904
rect 103296 389892 103302 389904
rect 115290 389892 115296 389904
rect 103296 389864 115296 389892
rect 103296 389852 103302 389864
rect 115290 389852 115296 389864
rect 115348 389852 115354 389904
rect 130378 389852 130384 389904
rect 130436 389892 130442 389904
rect 139394 389892 139400 389904
rect 130436 389864 139400 389892
rect 130436 389852 130442 389864
rect 139394 389852 139400 389864
rect 139452 389852 139458 389904
rect 49510 389784 49516 389836
rect 49568 389824 49574 389836
rect 82814 389824 82820 389836
rect 49568 389796 82820 389824
rect 49568 389784 49574 389796
rect 82814 389784 82820 389796
rect 82872 389784 82878 389836
rect 96522 389784 96528 389836
rect 96580 389824 96586 389836
rect 130102 389824 130108 389836
rect 96580 389796 130108 389824
rect 96580 389784 96586 389796
rect 130102 389784 130108 389796
rect 130160 389824 130166 389836
rect 142430 389824 142436 389836
rect 130160 389796 142436 389824
rect 130160 389784 130166 389796
rect 142430 389784 142436 389796
rect 142488 389784 142494 389836
rect 57790 389308 57796 389360
rect 57848 389348 57854 389360
rect 104526 389348 104532 389360
rect 57848 389320 104532 389348
rect 57848 389308 57854 389320
rect 104526 389308 104532 389320
rect 104584 389308 104590 389360
rect 114278 389308 114284 389360
rect 114336 389348 114342 389360
rect 118786 389348 118792 389360
rect 114336 389320 118792 389348
rect 114336 389308 114342 389320
rect 118786 389308 118792 389320
rect 118844 389308 118850 389360
rect 119338 389308 119344 389360
rect 119396 389348 119402 389360
rect 128538 389348 128544 389360
rect 119396 389320 128544 389348
rect 119396 389308 119402 389320
rect 128538 389308 128544 389320
rect 128596 389308 128602 389360
rect 57238 389240 57244 389292
rect 57296 389280 57302 389292
rect 57606 389280 57612 389292
rect 57296 389252 57612 389280
rect 57296 389240 57302 389252
rect 57606 389240 57612 389252
rect 57664 389280 57670 389292
rect 79318 389280 79324 389292
rect 57664 389252 79324 389280
rect 57664 389240 57670 389252
rect 79318 389240 79324 389252
rect 79376 389240 79382 389292
rect 101030 389240 101036 389292
rect 101088 389280 101094 389292
rect 102042 389280 102048 389292
rect 101088 389252 102048 389280
rect 101088 389240 101094 389252
rect 102042 389240 102048 389252
rect 102100 389280 102106 389292
rect 128354 389280 128360 389292
rect 102100 389252 128360 389280
rect 102100 389240 102106 389252
rect 128354 389240 128360 389252
rect 128412 389240 128418 389292
rect 102594 389172 102600 389224
rect 102652 389212 102658 389224
rect 136910 389212 136916 389224
rect 102652 389184 136916 389212
rect 102652 389172 102658 389184
rect 136910 389172 136916 389184
rect 136968 389212 136974 389224
rect 198090 389212 198096 389224
rect 136968 389184 198096 389212
rect 136968 389172 136974 389184
rect 198090 389172 198096 389184
rect 198148 389172 198154 389224
rect 37090 389104 37096 389156
rect 37148 389144 37154 389156
rect 37148 389116 64874 389144
rect 37148 389104 37154 389116
rect 64846 389076 64874 389116
rect 71038 389104 71044 389156
rect 71096 389144 71102 389156
rect 74810 389144 74816 389156
rect 71096 389116 74816 389144
rect 71096 389104 71102 389116
rect 74810 389104 74816 389116
rect 74868 389104 74874 389156
rect 115750 389104 115756 389156
rect 115808 389144 115814 389156
rect 119338 389144 119344 389156
rect 115808 389116 119344 389144
rect 115808 389104 115814 389116
rect 119338 389104 119344 389116
rect 119396 389104 119402 389156
rect 72418 389076 72424 389088
rect 64846 389048 72424 389076
rect 72418 389036 72424 389048
rect 72476 389036 72482 389088
rect 98454 388628 98460 388680
rect 98512 388668 98518 388680
rect 109402 388668 109408 388680
rect 98512 388640 109408 388668
rect 98512 388628 98518 388640
rect 109402 388628 109408 388640
rect 109460 388628 109466 388680
rect 97902 388560 97908 388612
rect 97960 388600 97966 388612
rect 111794 388600 111800 388612
rect 97960 388572 111800 388600
rect 97960 388560 97966 388572
rect 111794 388560 111800 388572
rect 111852 388560 111858 388612
rect 91002 388492 91008 388544
rect 91060 388532 91066 388544
rect 120074 388532 120080 388544
rect 91060 388504 120080 388532
rect 91060 388492 91066 388504
rect 120074 388492 120080 388504
rect 120132 388532 120138 388544
rect 122006 388532 122012 388544
rect 120132 388504 122012 388532
rect 120132 388492 120138 388504
rect 122006 388492 122012 388504
rect 122064 388492 122070 388544
rect 4798 388424 4804 388476
rect 4856 388464 4862 388476
rect 37090 388464 37096 388476
rect 4856 388436 37096 388464
rect 4856 388424 4862 388436
rect 37090 388424 37096 388436
rect 37148 388424 37154 388476
rect 41138 388424 41144 388476
rect 41196 388464 41202 388476
rect 48038 388464 48044 388476
rect 41196 388436 48044 388464
rect 41196 388424 41202 388436
rect 48038 388424 48044 388436
rect 48096 388464 48102 388476
rect 71774 388464 71780 388476
rect 48096 388436 71780 388464
rect 48096 388424 48102 388436
rect 71774 388424 71780 388436
rect 71832 388424 71838 388476
rect 86402 388424 86408 388476
rect 86460 388464 86466 388476
rect 98638 388464 98644 388476
rect 86460 388436 98644 388464
rect 86460 388424 86466 388436
rect 98638 388424 98644 388436
rect 98696 388424 98702 388476
rect 106918 388424 106924 388476
rect 106976 388464 106982 388476
rect 141050 388464 141056 388476
rect 106976 388436 141056 388464
rect 106976 388424 106982 388436
rect 141050 388424 141056 388436
rect 141108 388464 141114 388476
rect 204898 388464 204904 388476
rect 141108 388436 204904 388464
rect 141108 388424 141114 388436
rect 204898 388424 204904 388436
rect 204956 388424 204962 388476
rect 74902 388084 74908 388136
rect 74960 388124 74966 388136
rect 184198 388124 184204 388136
rect 74960 388096 184204 388124
rect 74960 388084 74966 388096
rect 184198 388084 184204 388096
rect 184256 388084 184262 388136
rect 112162 388016 112168 388068
rect 112220 388056 112226 388068
rect 112438 388056 112444 388068
rect 112220 388028 112444 388056
rect 112220 388016 112226 388028
rect 112438 388016 112444 388028
rect 112496 388056 112502 388068
rect 119338 388056 119344 388068
rect 112496 388028 119344 388056
rect 112496 388016 112502 388028
rect 119338 388016 119344 388028
rect 119396 388016 119402 388068
rect 58526 387948 58532 388000
rect 58584 387988 58590 388000
rect 87046 387988 87052 388000
rect 58584 387960 87052 387988
rect 58584 387948 58590 387960
rect 87046 387948 87052 387960
rect 87104 387948 87110 388000
rect 48958 387880 48964 387932
rect 49016 387920 49022 387932
rect 52362 387920 52368 387932
rect 49016 387892 52368 387920
rect 49016 387880 49022 387892
rect 52362 387880 52368 387892
rect 52420 387920 52426 387932
rect 92934 387920 92940 387932
rect 52420 387892 92940 387920
rect 52420 387880 52426 387892
rect 92934 387880 92940 387892
rect 92992 387880 92998 387932
rect 109586 387880 109592 387932
rect 109644 387920 109650 387932
rect 110322 387920 110328 387932
rect 109644 387892 110328 387920
rect 109644 387880 109650 387892
rect 110322 387880 110328 387892
rect 110380 387920 110386 387932
rect 200758 387920 200764 387932
rect 110380 387892 200764 387920
rect 110380 387880 110386 387892
rect 200758 387880 200764 387892
rect 200816 387880 200822 387932
rect 54938 387812 54944 387864
rect 54996 387852 55002 387864
rect 55122 387852 55128 387864
rect 54996 387824 55128 387852
rect 54996 387812 55002 387824
rect 55122 387812 55128 387824
rect 55180 387852 55186 387864
rect 69750 387852 69756 387864
rect 55180 387824 69756 387852
rect 55180 387812 55186 387824
rect 69750 387812 69756 387824
rect 69808 387812 69814 387864
rect 92842 387812 92848 387864
rect 92900 387852 92906 387864
rect 92900 387824 93854 387852
rect 92900 387812 92906 387824
rect 93826 387784 93854 387824
rect 108942 387812 108948 387864
rect 109000 387852 109006 387864
rect 115842 387852 115848 387864
rect 109000 387824 115848 387852
rect 109000 387812 109006 387824
rect 115842 387812 115848 387824
rect 115900 387812 115906 387864
rect 120258 387784 120264 387796
rect 93826 387756 120264 387784
rect 120258 387744 120264 387756
rect 120316 387744 120322 387796
rect 56410 387200 56416 387252
rect 56468 387240 56474 387252
rect 71958 387240 71964 387252
rect 56468 387212 71964 387240
rect 56468 387200 56474 387212
rect 71958 387200 71964 387212
rect 72016 387200 72022 387252
rect 70118 387132 70124 387184
rect 70176 387172 70182 387184
rect 87598 387172 87604 387184
rect 70176 387144 87604 387172
rect 70176 387132 70182 387144
rect 87598 387132 87604 387144
rect 87656 387132 87662 387184
rect 107378 387132 107384 387184
rect 107436 387172 107442 387184
rect 124398 387172 124404 387184
rect 107436 387144 124404 387172
rect 107436 387132 107442 387144
rect 124398 387132 124404 387144
rect 124456 387132 124462 387184
rect 48038 387064 48044 387116
rect 48096 387104 48102 387116
rect 74626 387104 74632 387116
rect 48096 387076 74632 387104
rect 48096 387064 48102 387076
rect 74626 387064 74632 387076
rect 74684 387064 74690 387116
rect 88978 387064 88984 387116
rect 89036 387104 89042 387116
rect 118694 387104 118700 387116
rect 89036 387076 118700 387104
rect 89036 387064 89042 387076
rect 118694 387064 118700 387076
rect 118752 387064 118758 387116
rect 50890 386520 50896 386572
rect 50948 386560 50954 386572
rect 80606 386560 80612 386572
rect 50948 386532 80612 386560
rect 50948 386520 50954 386532
rect 80606 386520 80612 386532
rect 80664 386520 80670 386572
rect 103882 386520 103888 386572
rect 103940 386560 103946 386572
rect 122098 386560 122104 386572
rect 103940 386532 122104 386560
rect 103940 386520 103946 386532
rect 122098 386520 122104 386532
rect 122156 386520 122162 386572
rect 39758 386452 39764 386504
rect 39816 386492 39822 386504
rect 103790 386492 103796 386504
rect 39816 386464 103796 386492
rect 39816 386452 39822 386464
rect 103790 386452 103796 386464
rect 103848 386492 103854 386504
rect 103974 386492 103980 386504
rect 103848 386464 103980 386492
rect 103848 386452 103854 386464
rect 103974 386452 103980 386464
rect 104032 386452 104038 386504
rect 110322 386452 110328 386504
rect 110380 386492 110386 386504
rect 132494 386492 132500 386504
rect 110380 386464 132500 386492
rect 110380 386452 110386 386464
rect 132494 386452 132500 386464
rect 132552 386452 132558 386504
rect 74810 386384 74816 386436
rect 74868 386424 74874 386436
rect 286318 386424 286324 386436
rect 74868 386396 286324 386424
rect 74868 386384 74874 386396
rect 286318 386384 286324 386396
rect 286376 386384 286382 386436
rect 104894 386316 104900 386368
rect 104952 386356 104958 386368
rect 105906 386356 105912 386368
rect 104952 386328 105912 386356
rect 104952 386316 104958 386328
rect 105906 386316 105912 386328
rect 105964 386316 105970 386368
rect 41230 385772 41236 385824
rect 41288 385812 41294 385824
rect 50798 385812 50804 385824
rect 41288 385784 50804 385812
rect 41288 385772 41294 385784
rect 50798 385772 50804 385784
rect 50856 385772 50862 385824
rect 46658 385704 46664 385756
rect 46716 385744 46722 385756
rect 78858 385744 78864 385756
rect 46716 385716 78864 385744
rect 46716 385704 46722 385716
rect 78858 385704 78864 385716
rect 78916 385704 78922 385756
rect 112714 385704 112720 385756
rect 112772 385744 112778 385756
rect 117406 385744 117412 385756
rect 112772 385716 117412 385744
rect 112772 385704 112778 385716
rect 117406 385704 117412 385716
rect 117464 385704 117470 385756
rect 43990 385636 43996 385688
rect 44048 385676 44054 385688
rect 100662 385676 100668 385688
rect 44048 385648 100668 385676
rect 44048 385636 44054 385648
rect 100662 385636 100668 385648
rect 100720 385676 100726 385688
rect 120258 385676 120264 385688
rect 100720 385648 120264 385676
rect 100720 385636 100726 385648
rect 120258 385636 120264 385648
rect 120316 385636 120322 385688
rect 77478 385336 77484 385348
rect 64846 385308 77484 385336
rect 50798 385024 50804 385076
rect 50856 385064 50862 385076
rect 64846 385064 64874 385308
rect 77478 385296 77484 385308
rect 77536 385296 77542 385348
rect 90266 385296 90272 385348
rect 90324 385336 90330 385348
rect 90324 385308 93854 385336
rect 90324 385296 90330 385308
rect 50856 385036 64874 385064
rect 93826 385064 93854 385308
rect 100018 385296 100024 385348
rect 100076 385336 100082 385348
rect 100076 385308 103514 385336
rect 100076 385296 100082 385308
rect 103486 385132 103514 385308
rect 106274 385296 106280 385348
rect 106332 385336 106338 385348
rect 106332 385308 113174 385336
rect 106332 385296 106338 385308
rect 113146 385200 113174 385308
rect 120074 385200 120080 385212
rect 113146 385172 120080 385200
rect 120074 385160 120080 385172
rect 120132 385160 120138 385212
rect 287698 385132 287704 385144
rect 103486 385104 287704 385132
rect 287698 385092 287704 385104
rect 287756 385092 287762 385144
rect 308398 385064 308404 385076
rect 93826 385036 308404 385064
rect 50856 385024 50862 385036
rect 308398 385024 308404 385036
rect 308456 385024 308462 385076
rect 115934 384956 115940 385008
rect 115992 384996 115998 385008
rect 128446 384996 128452 385008
rect 115992 384968 128452 384996
rect 115992 384956 115998 384968
rect 128446 384956 128452 384968
rect 128504 384956 128510 385008
rect 63126 383732 63132 383784
rect 63184 383772 63190 383784
rect 65886 383772 65892 383784
rect 63184 383744 65892 383772
rect 63184 383732 63190 383744
rect 65886 383732 65892 383744
rect 65944 383732 65950 383784
rect 34422 383664 34428 383716
rect 34480 383704 34486 383716
rect 68738 383704 68744 383716
rect 34480 383676 68744 383704
rect 34480 383664 34486 383676
rect 68738 383664 68744 383676
rect 68796 383664 68802 383716
rect 118510 383664 118516 383716
rect 118568 383704 118574 383716
rect 360838 383704 360844 383716
rect 118568 383676 360844 383704
rect 118568 383664 118574 383676
rect 360838 383664 360844 383676
rect 360896 383664 360902 383716
rect 118602 383596 118608 383648
rect 118660 383636 118666 383648
rect 136726 383636 136732 383648
rect 118660 383608 136732 383636
rect 118660 383596 118666 383608
rect 136726 383596 136732 383608
rect 136784 383596 136790 383648
rect 136726 382916 136732 382968
rect 136784 382956 136790 382968
rect 145098 382956 145104 382968
rect 136784 382928 145104 382956
rect 136784 382916 136790 382928
rect 145098 382916 145104 382928
rect 145156 382916 145162 382968
rect 41322 382236 41328 382288
rect 41380 382276 41386 382288
rect 67634 382276 67640 382288
rect 41380 382248 67640 382276
rect 41380 382236 41386 382248
rect 67634 382236 67640 382248
rect 67692 382236 67698 382288
rect 118602 381488 118608 381540
rect 118660 381528 118666 381540
rect 135346 381528 135352 381540
rect 118660 381500 135352 381528
rect 118660 381488 118666 381500
rect 135346 381488 135352 381500
rect 135404 381488 135410 381540
rect 49602 380808 49608 380860
rect 49660 380848 49666 380860
rect 67634 380848 67640 380860
rect 49660 380820 67640 380848
rect 49660 380808 49666 380820
rect 67634 380808 67640 380820
rect 67692 380808 67698 380860
rect 118602 380808 118608 380860
rect 118660 380848 118666 380860
rect 121454 380848 121460 380860
rect 118660 380820 121460 380848
rect 118660 380808 118666 380820
rect 121454 380808 121460 380820
rect 121512 380848 121518 380860
rect 122190 380848 122196 380860
rect 121512 380820 122196 380848
rect 121512 380808 121518 380820
rect 122190 380808 122196 380820
rect 122248 380808 122254 380860
rect 48130 380264 48136 380316
rect 48188 380304 48194 380316
rect 49602 380304 49608 380316
rect 48188 380276 49608 380304
rect 48188 380264 48194 380276
rect 49602 380264 49608 380276
rect 49660 380264 49666 380316
rect 118326 380128 118332 380180
rect 118384 380168 118390 380180
rect 295978 380168 295984 380180
rect 118384 380140 295984 380168
rect 118384 380128 118390 380140
rect 295978 380128 295984 380140
rect 296036 380128 296042 380180
rect 64230 379516 64236 379568
rect 64288 379556 64294 379568
rect 65978 379556 65984 379568
rect 64288 379528 65984 379556
rect 64288 379516 64294 379528
rect 65978 379516 65984 379528
rect 66036 379556 66042 379568
rect 67634 379556 67640 379568
rect 66036 379528 67640 379556
rect 66036 379516 66042 379528
rect 67634 379516 67640 379528
rect 67692 379516 67698 379568
rect 118602 378836 118608 378888
rect 118660 378876 118666 378888
rect 122834 378876 122840 378888
rect 118660 378848 122840 378876
rect 118660 378836 118666 378848
rect 122834 378836 122840 378848
rect 122892 378876 122898 378888
rect 123018 378876 123024 378888
rect 122892 378848 123024 378876
rect 122892 378836 122898 378848
rect 123018 378836 123024 378848
rect 123076 378836 123082 378888
rect 119338 378768 119344 378820
rect 119396 378808 119402 378820
rect 276658 378808 276664 378820
rect 119396 378780 276664 378808
rect 119396 378768 119402 378780
rect 276658 378768 276664 378780
rect 276716 378768 276722 378820
rect 519538 378768 519544 378820
rect 519596 378808 519602 378820
rect 579614 378808 579620 378820
rect 519596 378780 579620 378808
rect 519596 378768 519602 378780
rect 579614 378768 579620 378780
rect 579672 378768 579678 378820
rect 118602 378156 118608 378208
rect 118660 378196 118666 378208
rect 122190 378196 122196 378208
rect 118660 378168 122196 378196
rect 118660 378156 118666 378168
rect 122190 378156 122196 378168
rect 122248 378196 122254 378208
rect 122248 378168 122834 378196
rect 122248 378156 122254 378168
rect 122806 378128 122834 378168
rect 147950 378128 147956 378140
rect 122806 378100 147956 378128
rect 147950 378088 147956 378100
rect 148008 378088 148014 378140
rect 48222 377408 48228 377460
rect 48280 377448 48286 377460
rect 67634 377448 67640 377460
rect 48280 377420 67640 377448
rect 48280 377408 48286 377420
rect 67634 377408 67640 377420
rect 67692 377408 67698 377460
rect 147950 377408 147956 377460
rect 148008 377448 148014 377460
rect 441614 377448 441620 377460
rect 148008 377420 441620 377448
rect 148008 377408 148014 377420
rect 441614 377408 441620 377420
rect 441672 377408 441678 377460
rect 118418 376728 118424 376780
rect 118476 376768 118482 376780
rect 143626 376768 143632 376780
rect 118476 376740 143632 376768
rect 118476 376728 118482 376740
rect 143626 376728 143632 376740
rect 143684 376728 143690 376780
rect 118602 376660 118608 376712
rect 118660 376700 118666 376712
rect 146294 376700 146300 376712
rect 118660 376672 146300 376700
rect 118660 376660 118666 376672
rect 146294 376660 146300 376672
rect 146352 376700 146358 376712
rect 149054 376700 149060 376712
rect 146352 376672 149060 376700
rect 146352 376660 146358 376672
rect 149054 376660 149060 376672
rect 149112 376660 149118 376712
rect 117774 376252 117780 376304
rect 117832 376292 117838 376304
rect 120258 376292 120264 376304
rect 117832 376264 120264 376292
rect 117832 376252 117838 376264
rect 120258 376252 120264 376264
rect 120316 376252 120322 376304
rect 42610 375368 42616 375420
rect 42668 375408 42674 375420
rect 48222 375408 48228 375420
rect 42668 375380 48228 375408
rect 42668 375368 42674 375380
rect 48222 375368 48228 375380
rect 48280 375368 48286 375420
rect 43806 375300 43812 375352
rect 43864 375340 43870 375352
rect 69106 375340 69112 375352
rect 43864 375312 69112 375340
rect 43864 375300 43870 375312
rect 69106 375300 69112 375312
rect 69164 375300 69170 375352
rect 118602 375300 118608 375352
rect 118660 375340 118666 375352
rect 145006 375340 145012 375352
rect 118660 375312 145012 375340
rect 118660 375300 118666 375312
rect 145006 375300 145012 375312
rect 145064 375340 145070 375352
rect 146202 375340 146208 375352
rect 145064 375312 146208 375340
rect 145064 375300 145070 375312
rect 146202 375300 146208 375312
rect 146260 375300 146266 375352
rect 64506 374620 64512 374672
rect 64564 374660 64570 374672
rect 64782 374660 64788 374672
rect 64564 374632 64788 374660
rect 64564 374620 64570 374632
rect 64782 374620 64788 374632
rect 64840 374660 64846 374672
rect 67634 374660 67640 374672
rect 64840 374632 67640 374660
rect 64840 374620 64846 374632
rect 67634 374620 67640 374632
rect 67692 374620 67698 374672
rect 60366 373940 60372 373992
rect 60424 373980 60430 373992
rect 65886 373980 65892 373992
rect 60424 373952 65892 373980
rect 60424 373940 60430 373952
rect 65886 373940 65892 373952
rect 65944 373940 65950 373992
rect 118602 373940 118608 373992
rect 118660 373980 118666 373992
rect 151814 373980 151820 373992
rect 118660 373952 151820 373980
rect 118660 373940 118666 373952
rect 151814 373940 151820 373952
rect 151872 373940 151878 373992
rect 3234 372512 3240 372564
rect 3292 372552 3298 372564
rect 51718 372552 51724 372564
rect 3292 372524 51724 372552
rect 3292 372512 3298 372524
rect 51718 372512 51724 372524
rect 51776 372512 51782 372564
rect 61838 372512 61844 372564
rect 61896 372552 61902 372564
rect 67634 372552 67640 372564
rect 61896 372524 67640 372552
rect 61896 372512 61902 372524
rect 67634 372512 67640 372524
rect 67692 372512 67698 372564
rect 66070 371900 66076 371952
rect 66128 371940 66134 371952
rect 67726 371940 67732 371952
rect 66128 371912 67732 371940
rect 66128 371900 66134 371912
rect 67726 371900 67732 371912
rect 67784 371900 67790 371952
rect 60550 371832 60556 371884
rect 60608 371872 60614 371884
rect 69658 371872 69664 371884
rect 60608 371844 69664 371872
rect 60608 371832 60614 371844
rect 69658 371832 69664 371844
rect 69716 371832 69722 371884
rect 117866 370472 117872 370524
rect 117924 370512 117930 370524
rect 136726 370512 136732 370524
rect 117924 370484 136732 370512
rect 117924 370472 117930 370484
rect 136726 370472 136732 370484
rect 136784 370472 136790 370524
rect 65518 370132 65524 370184
rect 65576 370172 65582 370184
rect 68370 370172 68376 370184
rect 65576 370144 68376 370172
rect 65576 370132 65582 370144
rect 68370 370132 68376 370144
rect 68428 370132 68434 370184
rect 116026 369860 116032 369912
rect 116084 369900 116090 369912
rect 116210 369900 116216 369912
rect 116084 369872 116216 369900
rect 116084 369860 116090 369872
rect 116210 369860 116216 369872
rect 116268 369860 116274 369912
rect 118050 369860 118056 369912
rect 118108 369900 118114 369912
rect 151814 369900 151820 369912
rect 118108 369872 151820 369900
rect 118108 369860 118114 369872
rect 151814 369860 151820 369872
rect 151872 369860 151878 369912
rect 53650 369792 53656 369844
rect 53708 369832 53714 369844
rect 67634 369832 67640 369844
rect 53708 369804 67640 369832
rect 53708 369792 53714 369804
rect 67634 369792 67640 369804
rect 67692 369792 67698 369844
rect 117314 369112 117320 369164
rect 117372 369152 117378 369164
rect 120166 369152 120172 369164
rect 117372 369124 120172 369152
rect 117372 369112 117378 369124
rect 120166 369112 120172 369124
rect 120224 369152 120230 369164
rect 131114 369152 131120 369164
rect 120224 369124 131120 369152
rect 120224 369112 120230 369124
rect 131114 369112 131120 369124
rect 131172 369112 131178 369164
rect 117406 368568 117412 368620
rect 117464 368608 117470 368620
rect 117682 368608 117688 368620
rect 117464 368580 117688 368608
rect 117464 368568 117470 368580
rect 117682 368568 117688 368580
rect 117740 368568 117746 368620
rect 131390 368500 131396 368552
rect 131448 368540 131454 368552
rect 131758 368540 131764 368552
rect 131448 368512 131764 368540
rect 131448 368500 131454 368512
rect 131758 368500 131764 368512
rect 131816 368540 131822 368552
rect 146294 368540 146300 368552
rect 131816 368512 146300 368540
rect 131816 368500 131822 368512
rect 146294 368500 146300 368512
rect 146352 368500 146358 368552
rect 117406 368432 117412 368484
rect 117464 368472 117470 368484
rect 150618 368472 150624 368484
rect 117464 368444 150624 368472
rect 117464 368432 117470 368444
rect 150618 368432 150624 368444
rect 150676 368472 150682 368484
rect 151170 368472 151176 368484
rect 150676 368444 151176 368472
rect 150676 368432 150682 368444
rect 151170 368432 151176 368444
rect 151228 368432 151234 368484
rect 117314 368364 117320 368416
rect 117372 368404 117378 368416
rect 131390 368404 131396 368416
rect 117372 368376 131396 368404
rect 117372 368364 117378 368376
rect 131390 368364 131396 368376
rect 131448 368364 131454 368416
rect 60366 367752 60372 367804
rect 60424 367792 60430 367804
rect 69750 367792 69756 367804
rect 60424 367764 69756 367792
rect 60424 367752 60430 367764
rect 69750 367752 69756 367764
rect 69808 367752 69814 367804
rect 151170 367684 151176 367736
rect 151228 367724 151234 367736
rect 152090 367724 152096 367736
rect 151228 367696 152096 367724
rect 151228 367684 151234 367696
rect 152090 367684 152096 367696
rect 152148 367684 152154 367736
rect 60458 367004 60464 367056
rect 60516 367044 60522 367056
rect 68002 367044 68008 367056
rect 60516 367016 68008 367044
rect 60516 367004 60522 367016
rect 68002 367004 68008 367016
rect 68060 367004 68066 367056
rect 117314 367004 117320 367056
rect 117372 367044 117378 367056
rect 134058 367044 134064 367056
rect 117372 367016 134064 367044
rect 117372 367004 117378 367016
rect 134058 367004 134064 367016
rect 134116 367044 134122 367056
rect 136634 367044 136640 367056
rect 134116 367016 136640 367044
rect 134116 367004 134122 367016
rect 136634 367004 136640 367016
rect 136692 367004 136698 367056
rect 59170 366324 59176 366376
rect 59228 366364 59234 366376
rect 67634 366364 67640 366376
rect 59228 366336 67640 366364
rect 59228 366324 59234 366336
rect 67634 366324 67640 366336
rect 67692 366324 67698 366376
rect 136726 366324 136732 366376
rect 136784 366364 136790 366376
rect 579614 366364 579620 366376
rect 136784 366336 579620 366364
rect 136784 366324 136790 366336
rect 579614 366324 579620 366336
rect 579672 366324 579678 366376
rect 63218 365644 63224 365696
rect 63276 365684 63282 365696
rect 64690 365684 64696 365696
rect 63276 365656 64696 365684
rect 63276 365644 63282 365656
rect 64690 365644 64696 365656
rect 64748 365644 64754 365696
rect 119062 365644 119068 365696
rect 119120 365684 119126 365696
rect 129734 365684 129740 365696
rect 119120 365656 129740 365684
rect 119120 365644 119126 365656
rect 129734 365644 129740 365656
rect 129792 365644 129798 365696
rect 34330 365576 34336 365628
rect 34388 365616 34394 365628
rect 35158 365616 35164 365628
rect 34388 365588 35164 365616
rect 34388 365576 34394 365588
rect 35158 365576 35164 365588
rect 35216 365576 35222 365628
rect 119890 365032 119896 365084
rect 119948 365072 119954 365084
rect 146386 365072 146392 365084
rect 119948 365044 146392 365072
rect 119948 365032 119954 365044
rect 146386 365032 146392 365044
rect 146444 365032 146450 365084
rect 122098 364964 122104 365016
rect 122156 365004 122162 365016
rect 305638 365004 305644 365016
rect 122156 364976 305644 365004
rect 122156 364964 122162 364976
rect 305638 364964 305644 364976
rect 305696 364964 305702 365016
rect 117314 364828 117320 364880
rect 117372 364868 117378 364880
rect 119890 364868 119896 364880
rect 117372 364840 119896 364868
rect 117372 364828 117378 364840
rect 119890 364828 119896 364840
rect 119948 364828 119954 364880
rect 64690 364352 64696 364404
rect 64748 364392 64754 364404
rect 67634 364392 67640 364404
rect 64748 364364 67640 364392
rect 64748 364352 64754 364364
rect 67634 364352 67640 364364
rect 67692 364352 67698 364404
rect 50706 364284 50712 364336
rect 50764 364324 50770 364336
rect 67726 364324 67732 364336
rect 50764 364296 67732 364324
rect 50764 364284 50770 364296
rect 67726 364284 67732 364296
rect 67784 364284 67790 364336
rect 34330 363604 34336 363656
rect 34388 363644 34394 363656
rect 67634 363644 67640 363656
rect 34388 363616 67640 363644
rect 34388 363604 34394 363616
rect 67634 363604 67640 363616
rect 67692 363604 67698 363656
rect 117682 363604 117688 363656
rect 117740 363644 117746 363656
rect 307018 363644 307024 363656
rect 117740 363616 307024 363644
rect 117740 363604 117746 363616
rect 307018 363604 307024 363616
rect 307076 363604 307082 363656
rect 48222 362992 48228 363044
rect 48280 363032 48286 363044
rect 50706 363032 50712 363044
rect 48280 363004 50712 363032
rect 48280 362992 48286 363004
rect 50706 362992 50712 363004
rect 50764 362992 50770 363044
rect 42426 362924 42432 362976
rect 42484 362964 42490 362976
rect 59078 362964 59084 362976
rect 42484 362936 59084 362964
rect 42484 362924 42490 362936
rect 59078 362924 59084 362936
rect 59136 362924 59142 362976
rect 117314 362856 117320 362908
rect 117372 362896 117378 362908
rect 151998 362896 152004 362908
rect 117372 362868 152004 362896
rect 117372 362856 117378 362868
rect 151998 362856 152004 362868
rect 152056 362896 152062 362908
rect 153102 362896 153108 362908
rect 152056 362868 153108 362896
rect 152056 362856 152062 362868
rect 153102 362856 153108 362868
rect 153160 362856 153166 362908
rect 35710 362176 35716 362228
rect 35768 362216 35774 362228
rect 42426 362216 42432 362228
rect 35768 362188 42432 362216
rect 35768 362176 35774 362188
rect 42426 362176 42432 362188
rect 42484 362176 42490 362228
rect 117314 362176 117320 362228
rect 117372 362216 117378 362228
rect 121362 362216 121368 362228
rect 117372 362188 121368 362216
rect 117372 362176 117378 362188
rect 121362 362176 121368 362188
rect 121420 362216 121426 362228
rect 142338 362216 142344 362228
rect 121420 362188 142344 362216
rect 121420 362176 121426 362188
rect 142338 362176 142344 362188
rect 142396 362176 142402 362228
rect 153102 362176 153108 362228
rect 153160 362216 153166 362228
rect 191098 362216 191104 362228
rect 153160 362188 191104 362216
rect 153160 362176 153166 362188
rect 191098 362176 191104 362188
rect 191156 362176 191162 362228
rect 59078 361496 59084 361548
rect 59136 361536 59142 361548
rect 67634 361536 67640 361548
rect 59136 361508 67640 361536
rect 59136 361496 59142 361508
rect 67634 361496 67640 361508
rect 67692 361496 67698 361548
rect 141786 361496 141792 361548
rect 141844 361536 141850 361548
rect 142246 361536 142252 361548
rect 141844 361508 142252 361536
rect 141844 361496 141850 361508
rect 142246 361496 142252 361508
rect 142304 361496 142310 361548
rect 118878 360272 118884 360324
rect 118936 360312 118942 360324
rect 119982 360312 119988 360324
rect 118936 360284 119988 360312
rect 118936 360272 118942 360284
rect 119982 360272 119988 360284
rect 120040 360312 120046 360324
rect 134058 360312 134064 360324
rect 120040 360284 134064 360312
rect 120040 360272 120046 360284
rect 134058 360272 134064 360284
rect 134116 360272 134122 360324
rect 117314 360204 117320 360256
rect 117372 360244 117378 360256
rect 141418 360244 141424 360256
rect 117372 360216 141424 360244
rect 117372 360204 117378 360216
rect 141418 360204 141424 360216
rect 141476 360244 141482 360256
rect 141786 360244 141792 360256
rect 141476 360216 141792 360244
rect 141476 360204 141482 360216
rect 141786 360204 141792 360216
rect 141844 360204 141850 360256
rect 43714 359456 43720 359508
rect 43772 359496 43778 359508
rect 59078 359496 59084 359508
rect 43772 359468 59084 359496
rect 43772 359456 43778 359468
rect 59078 359456 59084 359468
rect 59136 359456 59142 359508
rect 59078 358776 59084 358828
rect 59136 358816 59142 358828
rect 67634 358816 67640 358828
rect 59136 358788 67640 358816
rect 59136 358776 59142 358788
rect 67634 358776 67640 358788
rect 67692 358776 67698 358828
rect 117866 358776 117872 358828
rect 117924 358816 117930 358828
rect 206278 358816 206284 358828
rect 117924 358788 206284 358816
rect 117924 358776 117930 358788
rect 206278 358776 206284 358788
rect 206336 358776 206342 358828
rect 36630 358028 36636 358080
rect 36688 358068 36694 358080
rect 53834 358068 53840 358080
rect 36688 358040 53840 358068
rect 36688 358028 36694 358040
rect 53834 358028 53840 358040
rect 53892 358028 53898 358080
rect 56502 358028 56508 358080
rect 56560 358068 56566 358080
rect 67634 358068 67640 358080
rect 56560 358040 67640 358068
rect 56560 358028 56566 358040
rect 67634 358028 67640 358040
rect 67692 358028 67698 358080
rect 118602 358028 118608 358080
rect 118660 358068 118666 358080
rect 121638 358068 121644 358080
rect 118660 358040 121644 358068
rect 118660 358028 118666 358040
rect 121638 358028 121644 358040
rect 121696 358068 121702 358080
rect 143534 358068 143540 358080
rect 121696 358040 143540 358068
rect 121696 358028 121702 358040
rect 143534 358028 143540 358040
rect 143592 358028 143598 358080
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 43438 357456 43444 357468
rect 3200 357428 43444 357456
rect 3200 357416 3206 357428
rect 43438 357416 43444 357428
rect 43496 357416 43502 357468
rect 53834 357416 53840 357468
rect 53892 357456 53898 357468
rect 54938 357456 54944 357468
rect 53892 357428 54944 357456
rect 53892 357416 53898 357428
rect 54938 357416 54944 357428
rect 54996 357456 55002 357468
rect 67726 357456 67732 357468
rect 54996 357428 67732 357456
rect 54996 357416 55002 357428
rect 67726 357416 67732 357428
rect 67784 357416 67790 357468
rect 131390 356668 131396 356720
rect 131448 356708 131454 356720
rect 138106 356708 138112 356720
rect 131448 356680 138112 356708
rect 131448 356668 131454 356680
rect 138106 356668 138112 356680
rect 138164 356668 138170 356720
rect 118602 356124 118608 356176
rect 118660 356164 118666 356176
rect 131390 356164 131396 356176
rect 118660 356136 131396 356164
rect 118660 356124 118666 356136
rect 131390 356124 131396 356136
rect 131448 356164 131454 356176
rect 131758 356164 131764 356176
rect 131448 356136 131764 356164
rect 131448 356124 131454 356136
rect 131758 356124 131764 356136
rect 131816 356124 131822 356176
rect 52270 356056 52276 356108
rect 52328 356096 52334 356108
rect 52328 356068 54524 356096
rect 52328 356056 52334 356068
rect 54496 356040 54524 356068
rect 59998 356056 60004 356108
rect 60056 356096 60062 356108
rect 60056 356068 65564 356096
rect 60056 356056 60062 356068
rect 54478 355988 54484 356040
rect 54536 356028 54542 356040
rect 65536 356028 65564 356068
rect 118142 356056 118148 356108
rect 118200 356096 118206 356108
rect 308490 356096 308496 356108
rect 118200 356068 308496 356096
rect 118200 356056 118206 356068
rect 308490 356056 308496 356068
rect 308548 356056 308554 356108
rect 67634 356028 67640 356040
rect 54536 356000 64874 356028
rect 65536 356000 67640 356028
rect 54536 355988 54542 356000
rect 46842 355920 46848 355972
rect 46900 355960 46906 355972
rect 59998 355960 60004 355972
rect 46900 355932 60004 355960
rect 46900 355920 46906 355932
rect 59998 355920 60004 355932
rect 60056 355920 60062 355972
rect 64846 355960 64874 356000
rect 67634 355988 67640 356000
rect 67692 355988 67698 356040
rect 67726 355960 67732 355972
rect 64846 355932 67732 355960
rect 67726 355920 67732 355932
rect 67784 355920 67790 355972
rect 118602 355308 118608 355360
rect 118660 355348 118666 355360
rect 280798 355348 280804 355360
rect 118660 355320 280804 355348
rect 118660 355308 118666 355320
rect 280798 355308 280804 355320
rect 280856 355308 280862 355360
rect 118510 354628 118516 354680
rect 118568 354668 118574 354680
rect 140958 354668 140964 354680
rect 118568 354640 140964 354668
rect 118568 354628 118574 354640
rect 140958 354628 140964 354640
rect 141016 354628 141022 354680
rect 118602 354016 118608 354068
rect 118660 354056 118666 354068
rect 124214 354056 124220 354068
rect 118660 354028 124220 354056
rect 118660 354016 118666 354028
rect 124214 354016 124220 354028
rect 124272 354016 124278 354068
rect 119338 353948 119344 354000
rect 119396 353988 119402 354000
rect 580350 353988 580356 354000
rect 119396 353960 580356 353988
rect 119396 353948 119402 353960
rect 580350 353948 580356 353960
rect 580408 353948 580414 354000
rect 62758 353268 62764 353320
rect 62816 353308 62822 353320
rect 67358 353308 67364 353320
rect 62816 353280 67364 353308
rect 62816 353268 62822 353280
rect 67358 353268 67364 353280
rect 67416 353308 67422 353320
rect 67634 353308 67640 353320
rect 67416 353280 67640 353308
rect 67416 353268 67422 353280
rect 67634 353268 67640 353280
rect 67692 353268 67698 353320
rect 124214 353268 124220 353320
rect 124272 353308 124278 353320
rect 125594 353308 125600 353320
rect 124272 353280 125600 353308
rect 124272 353268 124278 353280
rect 125594 353268 125600 353280
rect 125652 353268 125658 353320
rect 140958 353268 140964 353320
rect 141016 353308 141022 353320
rect 142246 353308 142252 353320
rect 141016 353280 142252 353308
rect 141016 353268 141022 353280
rect 142246 353268 142252 353280
rect 142304 353268 142310 353320
rect 61378 352588 61384 352640
rect 61436 352628 61442 352640
rect 67634 352628 67640 352640
rect 61436 352600 67640 352628
rect 61436 352588 61442 352600
rect 67634 352588 67640 352600
rect 67692 352588 67698 352640
rect 42794 352520 42800 352572
rect 42852 352560 42858 352572
rect 43898 352560 43904 352572
rect 42852 352532 43904 352560
rect 42852 352520 42858 352532
rect 43898 352520 43904 352532
rect 43956 352560 43962 352572
rect 68922 352560 68928 352572
rect 43956 352532 68928 352560
rect 43956 352520 43962 352532
rect 68922 352520 68928 352532
rect 68980 352520 68986 352572
rect 118602 352520 118608 352572
rect 118660 352560 118666 352572
rect 124214 352560 124220 352572
rect 118660 352532 124220 352560
rect 118660 352520 118666 352532
rect 124214 352520 124220 352532
rect 124272 352560 124278 352572
rect 125962 352560 125968 352572
rect 124272 352532 125968 352560
rect 124272 352520 124278 352532
rect 125962 352520 125968 352532
rect 126020 352520 126026 352572
rect 504358 352520 504364 352572
rect 504416 352560 504422 352572
rect 579614 352560 579620 352572
rect 504416 352532 579620 352560
rect 504416 352520 504422 352532
rect 579614 352520 579620 352532
rect 579672 352520 579678 352572
rect 7558 351908 7564 351960
rect 7616 351948 7622 351960
rect 42794 351948 42800 351960
rect 7616 351920 42800 351948
rect 7616 351908 7622 351920
rect 42794 351908 42800 351920
rect 42852 351908 42858 351960
rect 61378 351908 61384 351960
rect 61436 351948 61442 351960
rect 61838 351948 61844 351960
rect 61436 351920 61844 351948
rect 61436 351908 61442 351920
rect 61838 351908 61844 351920
rect 61896 351908 61902 351960
rect 118050 351840 118056 351892
rect 118108 351880 118114 351892
rect 147858 351880 147864 351892
rect 118108 351852 147864 351880
rect 118108 351840 118114 351852
rect 147858 351840 147864 351852
rect 147916 351840 147922 351892
rect 118602 351228 118608 351280
rect 118660 351268 118666 351280
rect 158714 351268 158720 351280
rect 118660 351240 158720 351268
rect 118660 351228 118666 351240
rect 158714 351228 158720 351240
rect 158772 351228 158778 351280
rect 63310 351160 63316 351212
rect 63368 351200 63374 351212
rect 67910 351200 67916 351212
rect 63368 351172 67916 351200
rect 63368 351160 63374 351172
rect 67910 351160 67916 351172
rect 67968 351160 67974 351212
rect 147858 351160 147864 351212
rect 147916 351200 147922 351212
rect 213178 351200 213184 351212
rect 147916 351172 213184 351200
rect 147916 351160 147922 351172
rect 213178 351160 213184 351172
rect 213236 351160 213242 351212
rect 46842 350548 46848 350600
rect 46900 350588 46906 350600
rect 46900 350560 55214 350588
rect 46900 350548 46906 350560
rect 55186 350520 55214 350560
rect 55858 350520 55864 350532
rect 55186 350492 55864 350520
rect 55858 350480 55864 350492
rect 55916 350520 55922 350532
rect 67634 350520 67640 350532
rect 55916 350492 67640 350520
rect 55916 350480 55922 350492
rect 67634 350480 67640 350492
rect 67692 350480 67698 350532
rect 118602 349800 118608 349852
rect 118660 349840 118666 349852
rect 133966 349840 133972 349852
rect 118660 349812 133972 349840
rect 118660 349800 118666 349812
rect 133966 349800 133972 349812
rect 134024 349800 134030 349852
rect 66162 349732 66168 349784
rect 66220 349772 66226 349784
rect 68370 349772 68376 349784
rect 66220 349744 68376 349772
rect 66220 349732 66226 349744
rect 68370 349732 68376 349744
rect 68428 349732 68434 349784
rect 63310 349120 63316 349172
rect 63368 349160 63374 349172
rect 66254 349160 66260 349172
rect 63368 349132 66260 349160
rect 63368 349120 63374 349132
rect 66254 349120 66260 349132
rect 66312 349160 66318 349172
rect 66312 349132 67128 349160
rect 66312 349120 66318 349132
rect 67100 349092 67128 349132
rect 67634 349092 67640 349104
rect 67100 349064 67640 349092
rect 67634 349052 67640 349064
rect 67692 349052 67698 349104
rect 118602 349052 118608 349104
rect 118660 349092 118666 349104
rect 139486 349092 139492 349104
rect 118660 349064 139492 349092
rect 118660 349052 118666 349064
rect 139486 349052 139492 349064
rect 139544 349092 139550 349104
rect 139762 349092 139768 349104
rect 139544 349064 139768 349092
rect 139544 349052 139550 349064
rect 139762 349052 139768 349064
rect 139820 349052 139826 349104
rect 139762 348372 139768 348424
rect 139820 348412 139826 348424
rect 180058 348412 180064 348424
rect 139820 348384 180064 348412
rect 139820 348372 139826 348384
rect 180058 348372 180064 348384
rect 180116 348372 180122 348424
rect 57882 347760 57888 347812
rect 57940 347800 57946 347812
rect 57940 347772 64874 347800
rect 57940 347760 57946 347772
rect 64846 347732 64874 347772
rect 117866 347760 117872 347812
rect 117924 347800 117930 347812
rect 297358 347800 297364 347812
rect 117924 347772 297364 347800
rect 117924 347760 117930 347772
rect 297358 347760 297364 347772
rect 297416 347760 297422 347812
rect 67726 347732 67732 347744
rect 64846 347704 67732 347732
rect 67726 347692 67732 347704
rect 67784 347692 67790 347744
rect 117406 347692 117412 347744
rect 117464 347732 117470 347744
rect 149146 347732 149152 347744
rect 117464 347704 149152 347732
rect 117464 347692 117470 347704
rect 149146 347692 149152 347704
rect 149204 347732 149210 347744
rect 149698 347732 149704 347744
rect 149204 347704 149704 347732
rect 149204 347692 149210 347704
rect 149698 347692 149704 347704
rect 149756 347692 149762 347744
rect 149698 347080 149704 347132
rect 149756 347120 149762 347132
rect 215938 347120 215944 347132
rect 149756 347092 215944 347120
rect 149756 347080 149762 347092
rect 215938 347080 215944 347092
rect 215996 347080 216002 347132
rect 64598 347012 64604 347064
rect 64656 347052 64662 347064
rect 67634 347052 67640 347064
rect 64656 347024 67640 347052
rect 64656 347012 64662 347024
rect 67634 347012 67640 347024
rect 67692 347012 67698 347064
rect 158714 347012 158720 347064
rect 158772 347052 158778 347064
rect 347038 347052 347044 347064
rect 158772 347024 347044 347052
rect 158772 347012 158778 347024
rect 347038 347012 347044 347024
rect 347096 347012 347102 347064
rect 43438 346332 43444 346384
rect 43496 346372 43502 346384
rect 68186 346372 68192 346384
rect 43496 346344 68192 346372
rect 43496 346332 43502 346344
rect 68186 346332 68192 346344
rect 68244 346332 68250 346384
rect 118602 346332 118608 346384
rect 118660 346372 118666 346384
rect 132586 346372 132592 346384
rect 118660 346344 132592 346372
rect 118660 346332 118666 346344
rect 132586 346332 132592 346344
rect 132644 346372 132650 346384
rect 133782 346372 133788 346384
rect 132644 346344 133788 346372
rect 132644 346332 132650 346344
rect 133782 346332 133788 346344
rect 133840 346332 133846 346384
rect 2774 346264 2780 346316
rect 2832 346304 2838 346316
rect 4798 346304 4804 346316
rect 2832 346276 4804 346304
rect 2832 346264 2838 346276
rect 4798 346264 4804 346276
rect 4856 346264 4862 346316
rect 151906 345760 151912 345772
rect 122806 345732 151912 345760
rect 118510 345652 118516 345704
rect 118568 345692 118574 345704
rect 122098 345692 122104 345704
rect 118568 345664 122104 345692
rect 118568 345652 118574 345664
rect 122098 345652 122104 345664
rect 122156 345692 122162 345704
rect 122806 345692 122834 345732
rect 151906 345720 151912 345732
rect 151964 345720 151970 345772
rect 122156 345664 122834 345692
rect 122156 345652 122162 345664
rect 133782 345652 133788 345704
rect 133840 345692 133846 345704
rect 209038 345692 209044 345704
rect 133840 345664 209044 345692
rect 133840 345652 133846 345664
rect 209038 345652 209044 345664
rect 209096 345652 209102 345704
rect 53650 345040 53656 345092
rect 53708 345080 53714 345092
rect 68646 345080 68652 345092
rect 53708 345052 68652 345080
rect 53708 345040 53714 345052
rect 68646 345040 68652 345052
rect 68704 345040 68710 345092
rect 118602 344972 118608 345024
rect 118660 345012 118666 345024
rect 140866 345012 140872 345024
rect 118660 344984 140872 345012
rect 118660 344972 118666 344984
rect 140866 344972 140872 344984
rect 140924 344972 140930 345024
rect 45462 344292 45468 344344
rect 45520 344332 45526 344344
rect 49418 344332 49424 344344
rect 45520 344304 49424 344332
rect 45520 344292 45526 344304
rect 49418 344292 49424 344304
rect 49476 344292 49482 344344
rect 140866 344292 140872 344344
rect 140924 344332 140930 344344
rect 305730 344332 305736 344344
rect 140924 344304 305736 344332
rect 140924 344292 140930 344304
rect 305730 344292 305736 344304
rect 305788 344292 305794 344344
rect 49418 343612 49424 343664
rect 49476 343652 49482 343664
rect 67634 343652 67640 343664
rect 49476 343624 67640 343652
rect 49476 343612 49482 343624
rect 67634 343612 67640 343624
rect 67692 343612 67698 343664
rect 117774 343544 117780 343596
rect 117832 343584 117838 343596
rect 143718 343584 143724 343596
rect 117832 343556 143724 343584
rect 117832 343544 117838 343556
rect 143718 343544 143724 343556
rect 143776 343584 143782 343596
rect 144822 343584 144828 343596
rect 143776 343556 144828 343584
rect 143776 343544 143782 343556
rect 144822 343544 144828 343556
rect 144880 343544 144886 343596
rect 118602 342864 118608 342916
rect 118660 342904 118666 342916
rect 126146 342904 126152 342916
rect 118660 342876 126152 342904
rect 118660 342864 118666 342876
rect 126146 342864 126152 342876
rect 126204 342864 126210 342916
rect 144822 342864 144828 342916
rect 144880 342904 144886 342916
rect 278038 342904 278044 342916
rect 144880 342876 278044 342904
rect 144880 342864 144886 342876
rect 278038 342864 278044 342876
rect 278096 342864 278102 342916
rect 126146 342320 126152 342372
rect 126204 342360 126210 342372
rect 128446 342360 128452 342372
rect 126204 342332 128452 342360
rect 126204 342320 126210 342332
rect 128446 342320 128452 342332
rect 128504 342320 128510 342372
rect 61930 342252 61936 342304
rect 61988 342292 61994 342304
rect 67266 342292 67272 342304
rect 61988 342264 67272 342292
rect 61988 342252 61994 342264
rect 67266 342252 67272 342264
rect 67324 342292 67330 342304
rect 67634 342292 67640 342304
rect 67324 342264 67640 342292
rect 67324 342252 67330 342264
rect 67634 342252 67640 342264
rect 67692 342252 67698 342304
rect 140866 342292 140872 342304
rect 125520 342264 140872 342292
rect 118602 342184 118608 342236
rect 118660 342224 118666 342236
rect 124858 342224 124864 342236
rect 118660 342196 124864 342224
rect 118660 342184 118666 342196
rect 124858 342184 124864 342196
rect 124916 342224 124922 342236
rect 125520 342224 125548 342264
rect 140866 342252 140872 342264
rect 140924 342252 140930 342304
rect 124916 342196 125548 342224
rect 124916 342184 124922 342196
rect 115750 341572 115756 341624
rect 115808 341612 115814 341624
rect 128630 341612 128636 341624
rect 115808 341584 128636 341612
rect 115808 341572 115814 341584
rect 128630 341572 128636 341584
rect 128688 341572 128694 341624
rect 38562 341504 38568 341556
rect 38620 341544 38626 341556
rect 68646 341544 68652 341556
rect 38620 341516 68652 341544
rect 38620 341504 38626 341516
rect 68646 341504 68652 341516
rect 68704 341504 68710 341556
rect 124858 341504 124864 341556
rect 124916 341544 124922 341556
rect 133966 341544 133972 341556
rect 124916 341516 133972 341544
rect 124916 341504 124922 341516
rect 133966 341504 133972 341516
rect 134024 341544 134030 341556
rect 485038 341544 485044 341556
rect 134024 341516 485044 341544
rect 134024 341504 134030 341516
rect 485038 341504 485044 341516
rect 485096 341504 485102 341556
rect 117498 340212 117504 340264
rect 117556 340252 117562 340264
rect 150710 340252 150716 340264
rect 117556 340224 150716 340252
rect 117556 340212 117562 340224
rect 150710 340212 150716 340224
rect 150768 340212 150774 340264
rect 62022 340144 62028 340196
rect 62080 340184 62086 340196
rect 67910 340184 67916 340196
rect 62080 340156 67916 340184
rect 62080 340144 62086 340156
rect 67910 340144 67916 340156
rect 67968 340144 67974 340196
rect 118418 340144 118424 340196
rect 118476 340184 118482 340196
rect 147766 340184 147772 340196
rect 118476 340156 147772 340184
rect 118476 340144 118482 340156
rect 147766 340144 147772 340156
rect 147824 340184 147830 340196
rect 377398 340184 377404 340196
rect 147824 340156 377404 340184
rect 147824 340144 147830 340156
rect 377398 340144 377404 340156
rect 377456 340144 377462 340196
rect 70394 339940 70400 339992
rect 70452 339980 70458 339992
rect 71038 339980 71044 339992
rect 70452 339952 71044 339980
rect 70452 339940 70458 339952
rect 71038 339940 71044 339952
rect 71096 339940 71102 339992
rect 56410 339532 56416 339584
rect 56468 339572 56474 339584
rect 73246 339572 73252 339584
rect 56468 339544 73252 339572
rect 56468 339532 56474 339544
rect 73246 339532 73252 339544
rect 73304 339532 73310 339584
rect 107930 339532 107936 339584
rect 107988 339572 107994 339584
rect 131206 339572 131212 339584
rect 107988 339544 131212 339572
rect 107988 339532 107994 339544
rect 131206 339532 131212 339544
rect 131264 339532 131270 339584
rect 47946 339464 47952 339516
rect 48004 339504 48010 339516
rect 81618 339504 81624 339516
rect 48004 339476 81624 339504
rect 48004 339464 48010 339476
rect 81618 339464 81624 339476
rect 81676 339464 81682 339516
rect 113266 339464 113272 339516
rect 113324 339504 113330 339516
rect 113818 339504 113824 339516
rect 113324 339476 113824 339504
rect 113324 339464 113330 339476
rect 113818 339464 113824 339476
rect 113876 339504 113882 339516
rect 143810 339504 143816 339516
rect 113876 339476 143816 339504
rect 113876 339464 113882 339476
rect 143810 339464 143816 339476
rect 143868 339464 143874 339516
rect 52086 339396 52092 339448
rect 52144 339436 52150 339448
rect 86218 339436 86224 339448
rect 52144 339408 86224 339436
rect 52144 339396 52150 339408
rect 86218 339396 86224 339408
rect 86276 339396 86282 339448
rect 107378 339396 107384 339448
rect 107436 339436 107442 339448
rect 107562 339436 107568 339448
rect 107436 339408 107568 339436
rect 107436 339396 107442 339408
rect 107562 339396 107568 339408
rect 107620 339436 107626 339448
rect 132862 339436 132868 339448
rect 107620 339408 132868 339436
rect 107620 339396 107626 339408
rect 132862 339396 132868 339408
rect 132920 339396 132926 339448
rect 40678 339328 40684 339380
rect 40736 339368 40742 339380
rect 73890 339368 73896 339380
rect 40736 339340 73896 339368
rect 40736 339328 40742 339340
rect 73890 339328 73896 339340
rect 73948 339328 73954 339380
rect 53742 339260 53748 339312
rect 53800 339300 53806 339312
rect 86770 339300 86776 339312
rect 53800 339272 86776 339300
rect 53800 339260 53806 339272
rect 86770 339260 86776 339272
rect 86828 339260 86834 339312
rect 60366 339192 60372 339244
rect 60424 339232 60430 339244
rect 89990 339232 89996 339244
rect 60424 339204 89996 339232
rect 60424 339192 60430 339204
rect 89990 339192 89996 339204
rect 90048 339232 90054 339244
rect 90358 339232 90364 339244
rect 90048 339204 90364 339232
rect 90048 339192 90054 339204
rect 90358 339192 90364 339204
rect 90416 339192 90422 339244
rect 113082 338920 113088 338972
rect 113140 338960 113146 338972
rect 118786 338960 118792 338972
rect 113140 338932 118792 338960
rect 113140 338920 113146 338932
rect 118786 338920 118792 338932
rect 118844 338920 118850 338972
rect 70302 338852 70308 338904
rect 70360 338892 70366 338904
rect 98638 338892 98644 338904
rect 70360 338864 98644 338892
rect 70360 338852 70366 338864
rect 98638 338852 98644 338864
rect 98696 338852 98702 338904
rect 112438 338852 112444 338904
rect 112496 338892 112502 338904
rect 122190 338892 122196 338904
rect 112496 338864 122196 338892
rect 112496 338852 112502 338864
rect 122190 338852 122196 338864
rect 122248 338852 122254 338904
rect 70486 338784 70492 338836
rect 70544 338824 70550 338836
rect 309778 338824 309784 338836
rect 70544 338796 309784 338824
rect 70544 338784 70550 338796
rect 309778 338784 309784 338796
rect 309836 338784 309842 338836
rect 97902 338716 97908 338768
rect 97960 338756 97966 338768
rect 124398 338756 124404 338768
rect 97960 338728 124404 338756
rect 97960 338716 97966 338728
rect 124398 338716 124404 338728
rect 124456 338756 124462 338768
rect 506474 338756 506480 338768
rect 124456 338728 506480 338756
rect 124456 338716 124462 338728
rect 506474 338716 506480 338728
rect 506532 338756 506538 338768
rect 580258 338756 580264 338768
rect 506532 338728 580264 338756
rect 506532 338716 506538 338728
rect 580258 338716 580264 338728
rect 580316 338716 580322 338768
rect 70670 338144 70676 338156
rect 69952 338116 70676 338144
rect 38470 338036 38476 338088
rect 38528 338076 38534 338088
rect 69952 338076 69980 338116
rect 70670 338104 70676 338116
rect 70728 338104 70734 338156
rect 38528 338048 69980 338076
rect 38528 338036 38534 338048
rect 70026 338036 70032 338088
rect 70084 338076 70090 338088
rect 71774 338076 71780 338088
rect 70084 338048 71780 338076
rect 70084 338036 70090 338048
rect 71774 338036 71780 338048
rect 71832 338036 71838 338088
rect 87414 338036 87420 338088
rect 87472 338076 87478 338088
rect 96706 338076 96712 338088
rect 87472 338048 96712 338076
rect 87472 338036 87478 338048
rect 96706 338036 96712 338048
rect 96764 338076 96770 338088
rect 97902 338076 97908 338088
rect 96764 338048 97908 338076
rect 96764 338036 96770 338048
rect 97902 338036 97908 338048
rect 97960 338036 97966 338088
rect 102134 338036 102140 338088
rect 102192 338076 102198 338088
rect 109954 338076 109960 338088
rect 102192 338048 109960 338076
rect 102192 338036 102198 338048
rect 109954 338036 109960 338048
rect 110012 338036 110018 338088
rect 112530 338036 112536 338088
rect 112588 338076 112594 338088
rect 138106 338076 138112 338088
rect 112588 338048 138112 338076
rect 112588 338036 112594 338048
rect 138106 338036 138112 338048
rect 138164 338036 138170 338088
rect 48038 337968 48044 338020
rect 48096 338008 48102 338020
rect 76466 338008 76472 338020
rect 48096 337980 76472 338008
rect 48096 337968 48102 337980
rect 76466 337968 76472 337980
rect 76524 337968 76530 338020
rect 86770 337968 86776 338020
rect 86828 338008 86834 338020
rect 87598 338008 87604 338020
rect 86828 337980 87604 338008
rect 86828 337968 86834 337980
rect 87598 337968 87604 337980
rect 87656 337968 87662 338020
rect 115106 337968 115112 338020
rect 115164 338008 115170 338020
rect 140774 338008 140780 338020
rect 115164 337980 140780 338008
rect 115164 337968 115170 337980
rect 140774 337968 140780 337980
rect 140832 337968 140838 338020
rect 44818 337900 44824 337952
rect 44876 337940 44882 337952
rect 71314 337940 71320 337952
rect 44876 337912 71320 337940
rect 44876 337900 44882 337912
rect 71314 337900 71320 337912
rect 71372 337900 71378 337952
rect 100294 337900 100300 337952
rect 100352 337940 100358 337952
rect 125778 337940 125784 337952
rect 100352 337912 125784 337940
rect 100352 337900 100358 337912
rect 125778 337900 125784 337912
rect 125836 337940 125842 337952
rect 126882 337940 126888 337952
rect 125836 337912 126888 337940
rect 125836 337900 125842 337912
rect 126882 337900 126888 337912
rect 126940 337900 126946 337952
rect 53098 337832 53104 337884
rect 53156 337872 53162 337884
rect 74534 337872 74540 337884
rect 53156 337844 74540 337872
rect 53156 337832 53162 337844
rect 74534 337832 74540 337844
rect 74592 337872 74598 337884
rect 75178 337872 75184 337884
rect 74592 337844 75184 337872
rect 74592 337832 74598 337844
rect 75178 337832 75184 337844
rect 75236 337832 75242 337884
rect 95786 337832 95792 337884
rect 95844 337872 95850 337884
rect 120166 337872 120172 337884
rect 95844 337844 120172 337872
rect 95844 337832 95850 337844
rect 120166 337832 120172 337844
rect 120224 337832 120230 337884
rect 76558 337696 76564 337748
rect 76616 337736 76622 337748
rect 78398 337736 78404 337748
rect 76616 337708 78404 337736
rect 76616 337696 76622 337708
rect 78398 337696 78404 337708
rect 78456 337696 78462 337748
rect 91278 337696 91284 337748
rect 91336 337736 91342 337748
rect 93670 337736 93676 337748
rect 91336 337708 93676 337736
rect 91336 337696 91342 337708
rect 93670 337696 93676 337708
rect 93728 337696 93734 337748
rect 73246 337560 73252 337612
rect 73304 337600 73310 337612
rect 91002 337600 91008 337612
rect 73304 337572 91008 337600
rect 73304 337560 73310 337572
rect 91002 337560 91008 337572
rect 91060 337560 91066 337612
rect 70670 337492 70676 337544
rect 70728 337532 70734 337544
rect 93302 337532 93308 337544
rect 70728 337504 93308 337532
rect 70728 337492 70734 337504
rect 93302 337492 93308 337504
rect 93360 337492 93366 337544
rect 126882 337492 126888 337544
rect 126940 337532 126946 337544
rect 140774 337532 140780 337544
rect 126940 337504 140780 337532
rect 126940 337492 126946 337504
rect 140774 337492 140780 337504
rect 140832 337492 140838 337544
rect 58986 337424 58992 337476
rect 59044 337464 59050 337476
rect 84194 337464 84200 337476
rect 59044 337436 84200 337464
rect 59044 337424 59050 337436
rect 84194 337424 84200 337436
rect 84252 337424 84258 337476
rect 99650 337424 99656 337476
rect 99708 337464 99714 337476
rect 102042 337464 102048 337476
rect 99708 337436 102048 337464
rect 99708 337424 99714 337436
rect 102042 337424 102048 337436
rect 102100 337464 102106 337476
rect 125686 337464 125692 337476
rect 102100 337436 125692 337464
rect 102100 337424 102106 337436
rect 125686 337424 125692 337436
rect 125744 337424 125750 337476
rect 138106 337424 138112 337476
rect 138164 337464 138170 337476
rect 177298 337464 177304 337476
rect 138164 337436 177304 337464
rect 138164 337424 138170 337436
rect 177298 337424 177304 337436
rect 177356 337424 177362 337476
rect 81618 337356 81624 337408
rect 81676 337396 81682 337408
rect 211798 337396 211804 337408
rect 81676 337368 211804 337396
rect 81676 337356 81682 337368
rect 211798 337356 211804 337368
rect 211856 337356 211862 337408
rect 97074 337016 97080 337068
rect 97132 337056 97138 337068
rect 100018 337056 100024 337068
rect 97132 337028 100024 337056
rect 97132 337016 97138 337028
rect 100018 337016 100024 337028
rect 100076 337016 100082 337068
rect 71314 336880 71320 336932
rect 71372 336920 71378 336932
rect 76650 336920 76656 336932
rect 71372 336892 76656 336920
rect 71372 336880 71378 336892
rect 76650 336880 76656 336892
rect 76708 336880 76714 336932
rect 120166 336744 120172 336796
rect 120224 336784 120230 336796
rect 320818 336784 320824 336796
rect 120224 336756 320824 336784
rect 120224 336744 120230 336756
rect 320818 336744 320824 336756
rect 320876 336744 320882 336796
rect 49510 336676 49516 336728
rect 49568 336716 49574 336728
rect 49568 336688 79272 336716
rect 49568 336676 49574 336688
rect 52178 336608 52184 336660
rect 52236 336648 52242 336660
rect 53742 336648 53748 336660
rect 52236 336620 53748 336648
rect 52236 336608 52242 336620
rect 53742 336608 53748 336620
rect 53800 336608 53806 336660
rect 79134 336648 79140 336660
rect 53944 336620 79140 336648
rect 39666 336540 39672 336592
rect 39724 336580 39730 336592
rect 39724 336552 45554 336580
rect 39724 336540 39730 336552
rect 45526 336444 45554 336552
rect 46750 336472 46756 336524
rect 46808 336512 46814 336524
rect 53944 336512 53972 336620
rect 79134 336608 79140 336620
rect 79192 336608 79198 336660
rect 79244 336648 79272 336688
rect 79318 336676 79324 336728
rect 79376 336716 79382 336728
rect 79686 336716 79692 336728
rect 79376 336688 79692 336716
rect 79376 336676 79382 336688
rect 79686 336676 79692 336688
rect 79744 336676 79750 336728
rect 106090 336676 106096 336728
rect 106148 336716 106154 336728
rect 127066 336716 127072 336728
rect 106148 336688 127072 336716
rect 106148 336676 106154 336688
rect 127066 336676 127072 336688
rect 127124 336676 127130 336728
rect 83458 336648 83464 336660
rect 79244 336620 83464 336648
rect 83458 336608 83464 336620
rect 83516 336608 83522 336660
rect 104158 336608 104164 336660
rect 104216 336648 104222 336660
rect 104802 336648 104808 336660
rect 104216 336620 104808 336648
rect 104216 336608 104222 336620
rect 104802 336608 104808 336620
rect 104860 336648 104866 336660
rect 122926 336648 122932 336660
rect 104860 336620 122932 336648
rect 104860 336608 104866 336620
rect 122926 336608 122932 336620
rect 122984 336608 122990 336660
rect 71958 336580 71964 336592
rect 46808 336484 53972 336512
rect 55186 336552 71964 336580
rect 46808 336472 46814 336484
rect 55186 336444 55214 336552
rect 71958 336540 71964 336552
rect 72016 336540 72022 336592
rect 57698 336472 57704 336524
rect 57756 336512 57762 336524
rect 88978 336512 88984 336524
rect 57756 336484 88984 336512
rect 57756 336472 57762 336484
rect 88978 336472 88984 336484
rect 89036 336472 89042 336524
rect 45526 336416 55214 336444
rect 56318 336404 56324 336456
rect 56376 336444 56382 336456
rect 79318 336444 79324 336456
rect 56376 336416 79324 336444
rect 56376 336404 56382 336416
rect 79318 336404 79324 336416
rect 79376 336404 79382 336456
rect 53742 335996 53748 336048
rect 53800 336036 53806 336048
rect 84838 336036 84844 336048
rect 53800 336008 84844 336036
rect 53800 335996 53806 336008
rect 84838 335996 84844 336008
rect 84896 335996 84902 336048
rect 60550 335248 60556 335300
rect 60608 335288 60614 335300
rect 98362 335288 98368 335300
rect 60608 335260 98368 335288
rect 60608 335248 60614 335260
rect 98362 335248 98368 335260
rect 98420 335248 98426 335300
rect 103514 335248 103520 335300
rect 103572 335288 103578 335300
rect 129918 335288 129924 335300
rect 103572 335260 129924 335288
rect 103572 335248 103578 335260
rect 129918 335248 129924 335260
rect 129976 335248 129982 335300
rect 42702 335180 42708 335232
rect 42760 335220 42766 335232
rect 75822 335220 75828 335232
rect 42760 335192 75828 335220
rect 42760 335180 42766 335192
rect 75822 335180 75828 335192
rect 75880 335180 75886 335232
rect 93670 335180 93676 335232
rect 93728 335220 93734 335232
rect 118694 335220 118700 335232
rect 93728 335192 118700 335220
rect 93728 335180 93734 335192
rect 118694 335180 118700 335192
rect 118752 335180 118758 335232
rect 44082 335112 44088 335164
rect 44140 335152 44146 335164
rect 76558 335152 76564 335164
rect 44140 335124 76564 335152
rect 44140 335112 44146 335124
rect 76558 335112 76564 335124
rect 76616 335112 76622 335164
rect 59262 334704 59268 334756
rect 59320 334744 59326 334756
rect 62022 334744 62028 334756
rect 59320 334716 62028 334744
rect 59320 334704 59326 334716
rect 62022 334704 62028 334716
rect 62080 334744 62086 334756
rect 94498 334744 94504 334756
rect 62080 334716 94504 334744
rect 62080 334704 62086 334716
rect 94498 334704 94504 334716
rect 94556 334704 94562 334756
rect 59170 334636 59176 334688
rect 59228 334676 59234 334688
rect 134610 334676 134616 334688
rect 59228 334648 134616 334676
rect 59228 334636 59234 334648
rect 134610 334636 134616 334648
rect 134668 334636 134674 334688
rect 71774 334568 71780 334620
rect 71832 334608 71838 334620
rect 291838 334608 291844 334620
rect 71832 334580 291844 334608
rect 71832 334568 71838 334580
rect 291838 334568 291844 334580
rect 291896 334568 291902 334620
rect 75270 334092 75276 334144
rect 75328 334132 75334 334144
rect 75822 334132 75828 334144
rect 75328 334104 75828 334132
rect 75328 334092 75334 334104
rect 75822 334092 75828 334104
rect 75880 334092 75886 334144
rect 56410 333956 56416 334008
rect 56468 333996 56474 334008
rect 60550 333996 60556 334008
rect 56468 333968 60556 333996
rect 56468 333956 56474 333968
rect 60550 333956 60556 333968
rect 60608 333956 60614 334008
rect 129734 333956 129740 334008
rect 129792 333996 129798 334008
rect 129918 333996 129924 334008
rect 129792 333968 129924 333996
rect 129792 333956 129798 333968
rect 129918 333956 129924 333968
rect 129976 333956 129982 334008
rect 46658 333888 46664 333940
rect 46716 333928 46722 333940
rect 80698 333928 80704 333940
rect 46716 333900 80704 333928
rect 46716 333888 46722 333900
rect 80698 333888 80704 333900
rect 80756 333888 80762 333940
rect 95050 333888 95056 333940
rect 95108 333928 95114 333940
rect 124306 333928 124312 333940
rect 95108 333900 124312 333928
rect 95108 333888 95114 333900
rect 124306 333888 124312 333900
rect 124364 333888 124370 333940
rect 60642 333820 60648 333872
rect 60700 333860 60706 333872
rect 92566 333860 92572 333872
rect 60700 333832 92572 333860
rect 60700 333820 60706 333832
rect 92566 333820 92572 333832
rect 92624 333820 92630 333872
rect 61838 333276 61844 333328
rect 61896 333316 61902 333328
rect 162118 333316 162124 333328
rect 61896 333288 162124 333316
rect 61896 333276 61902 333288
rect 162118 333276 162124 333288
rect 162176 333276 162182 333328
rect 71958 333208 71964 333260
rect 72016 333248 72022 333260
rect 309134 333248 309140 333260
rect 72016 333220 309140 333248
rect 72016 333208 72022 333220
rect 309134 333208 309140 333220
rect 309192 333208 309198 333260
rect 92566 332596 92572 332648
rect 92624 332636 92630 332648
rect 93118 332636 93124 332648
rect 92624 332608 93124 332636
rect 92624 332596 92630 332608
rect 93118 332596 93124 332608
rect 93176 332596 93182 332648
rect 113910 332528 113916 332580
rect 113968 332568 113974 332580
rect 144914 332568 144920 332580
rect 113968 332540 144920 332568
rect 113968 332528 113974 332540
rect 144914 332528 144920 332540
rect 144972 332568 144978 332580
rect 146202 332568 146208 332580
rect 144972 332540 146208 332568
rect 144972 332528 144978 332540
rect 146202 332528 146208 332540
rect 146260 332528 146266 332580
rect 113174 332052 113180 332104
rect 113232 332092 113238 332104
rect 113910 332092 113916 332104
rect 113232 332064 113916 332092
rect 113232 332052 113238 332064
rect 113910 332052 113916 332064
rect 113968 332052 113974 332104
rect 55030 331984 55036 332036
rect 55088 332024 55094 332036
rect 82262 332024 82268 332036
rect 55088 331996 82268 332024
rect 55088 331984 55094 331996
rect 82262 331984 82268 331996
rect 82320 331984 82326 332036
rect 95142 331984 95148 332036
rect 95200 332024 95206 332036
rect 113266 332024 113272 332036
rect 95200 331996 113272 332024
rect 95200 331984 95206 331996
rect 113266 331984 113272 331996
rect 113324 331984 113330 332036
rect 76466 331916 76472 331968
rect 76524 331956 76530 331968
rect 116578 331956 116584 331968
rect 76524 331928 116584 331956
rect 76524 331916 76530 331928
rect 116578 331916 116584 331928
rect 116636 331916 116642 331968
rect 54938 331848 54944 331900
rect 54996 331888 55002 331900
rect 117958 331888 117964 331900
rect 54996 331860 117964 331888
rect 54996 331848 55002 331860
rect 117958 331848 117964 331860
rect 118016 331848 118022 331900
rect 146202 331848 146208 331900
rect 146260 331888 146266 331900
rect 499574 331888 499580 331900
rect 146260 331860 499580 331888
rect 146260 331848 146266 331860
rect 499574 331848 499580 331860
rect 499632 331848 499638 331900
rect 67358 330488 67364 330540
rect 67416 330528 67422 330540
rect 77294 330528 77300 330540
rect 67416 330500 77300 330528
rect 67416 330488 67422 330500
rect 77294 330488 77300 330500
rect 77352 330488 77358 330540
rect 120166 329808 120172 329860
rect 120224 329848 120230 329860
rect 120718 329848 120724 329860
rect 120224 329820 120724 329848
rect 120224 329808 120230 329820
rect 120718 329808 120724 329820
rect 120776 329848 120782 329860
rect 125778 329848 125784 329860
rect 120776 329820 125784 329848
rect 120776 329808 120782 329820
rect 125778 329808 125784 329820
rect 125836 329808 125842 329860
rect 100938 329740 100944 329792
rect 100996 329780 101002 329792
rect 135254 329780 135260 329792
rect 100996 329752 135260 329780
rect 100996 329740 101002 329752
rect 135254 329740 135260 329752
rect 135312 329780 135318 329792
rect 136542 329780 136548 329792
rect 135312 329752 136548 329780
rect 135312 329740 135318 329752
rect 136542 329740 136548 329752
rect 136600 329740 136606 329792
rect 93210 329672 93216 329724
rect 93268 329712 93274 329724
rect 120166 329712 120172 329724
rect 93268 329684 120172 329712
rect 93268 329672 93274 329684
rect 120166 329672 120172 329684
rect 120224 329672 120230 329724
rect 93762 329060 93768 329112
rect 93820 329100 93826 329112
rect 115106 329100 115112 329112
rect 93820 329072 115112 329100
rect 93820 329060 93826 329072
rect 115106 329060 115112 329072
rect 115164 329060 115170 329112
rect 136542 329060 136548 329112
rect 136600 329100 136606 329112
rect 282178 329100 282184 329112
rect 136600 329072 282184 329100
rect 136600 329060 136606 329072
rect 282178 329060 282184 329072
rect 282236 329060 282242 329112
rect 89346 328380 89352 328432
rect 89404 328420 89410 328432
rect 123110 328420 123116 328432
rect 89404 328392 123116 328420
rect 89404 328380 89410 328392
rect 123110 328380 123116 328392
rect 123168 328420 123174 328432
rect 124122 328420 124128 328432
rect 123168 328392 124128 328420
rect 123168 328380 123174 328392
rect 124122 328380 124128 328392
rect 124180 328380 124186 328432
rect 97718 328312 97724 328364
rect 97776 328352 97782 328364
rect 130010 328352 130016 328364
rect 97776 328324 130016 328352
rect 97776 328312 97782 328324
rect 130010 328312 130016 328324
rect 130068 328352 130074 328364
rect 130378 328352 130384 328364
rect 130068 328324 130384 328352
rect 130068 328312 130074 328324
rect 130378 328312 130384 328324
rect 130436 328312 130442 328364
rect 124122 327768 124128 327820
rect 124180 327808 124186 327820
rect 242158 327808 242164 327820
rect 124180 327780 242164 327808
rect 124180 327768 124186 327780
rect 242158 327768 242164 327780
rect 242216 327768 242222 327820
rect 130378 327700 130384 327752
rect 130436 327740 130442 327752
rect 284938 327740 284944 327752
rect 130436 327712 284944 327740
rect 130436 327700 130442 327712
rect 284938 327700 284944 327712
rect 284996 327700 285002 327752
rect 110598 327020 110604 327072
rect 110656 327060 110662 327072
rect 136818 327060 136824 327072
rect 110656 327032 136824 327060
rect 110656 327020 110662 327032
rect 136818 327020 136824 327032
rect 136876 327060 136882 327072
rect 137094 327060 137100 327072
rect 136876 327032 137100 327060
rect 136876 327020 136882 327032
rect 137094 327020 137100 327032
rect 137152 327020 137158 327072
rect 65978 326340 65984 326392
rect 66036 326380 66042 326392
rect 115290 326380 115296 326392
rect 66036 326352 115296 326380
rect 66036 326340 66042 326352
rect 115290 326340 115296 326352
rect 115348 326340 115354 326392
rect 72418 325660 72424 325712
rect 72476 325700 72482 325712
rect 108298 325700 108304 325712
rect 72476 325672 108304 325700
rect 72476 325660 72482 325672
rect 108298 325660 108304 325672
rect 108356 325660 108362 325712
rect 111242 325592 111248 325644
rect 111300 325632 111306 325644
rect 132678 325632 132684 325644
rect 111300 325604 132684 325632
rect 111300 325592 111306 325604
rect 132678 325592 132684 325604
rect 132736 325632 132742 325644
rect 133782 325632 133788 325644
rect 132736 325604 133788 325632
rect 132736 325592 132742 325604
rect 133782 325592 133788 325604
rect 133840 325592 133846 325644
rect 106182 325048 106188 325100
rect 106240 325088 106246 325100
rect 115934 325088 115940 325100
rect 106240 325060 115940 325088
rect 106240 325048 106246 325060
rect 115934 325048 115940 325060
rect 115992 325048 115998 325100
rect 80698 324980 80704 325032
rect 80756 325020 80762 325032
rect 197998 325020 198004 325032
rect 80756 324992 198004 325020
rect 80756 324980 80762 324992
rect 197998 324980 198004 324992
rect 198056 324980 198062 325032
rect 48038 324912 48044 324964
rect 48096 324952 48102 324964
rect 107654 324952 107660 324964
rect 48096 324924 107660 324952
rect 48096 324912 48102 324924
rect 107654 324912 107660 324924
rect 107712 324912 107718 324964
rect 133782 324912 133788 324964
rect 133840 324952 133846 324964
rect 340138 324952 340144 324964
rect 133840 324924 340144 324952
rect 133840 324912 133846 324924
rect 340138 324912 340144 324924
rect 340196 324912 340202 324964
rect 14458 324300 14464 324352
rect 14516 324340 14522 324352
rect 48038 324340 48044 324352
rect 14516 324312 48044 324340
rect 14516 324300 14522 324312
rect 48038 324300 48044 324312
rect 48096 324300 48102 324352
rect 67450 323688 67456 323740
rect 67508 323728 67514 323740
rect 121454 323728 121460 323740
rect 67508 323700 121460 323728
rect 67508 323688 67514 323700
rect 121454 323688 121460 323700
rect 121512 323688 121518 323740
rect 93302 323620 93308 323672
rect 93360 323660 93366 323672
rect 265618 323660 265624 323672
rect 93360 323632 265624 323660
rect 93360 323620 93366 323632
rect 265618 323620 265624 323632
rect 265676 323620 265682 323672
rect 76650 323552 76656 323604
rect 76708 323592 76714 323604
rect 345658 323592 345664 323604
rect 76708 323564 345664 323592
rect 76708 323552 76714 323564
rect 345658 323552 345664 323564
rect 345716 323552 345722 323604
rect 86218 322260 86224 322312
rect 86276 322300 86282 322312
rect 147766 322300 147772 322312
rect 86276 322272 147772 322300
rect 86276 322260 86282 322272
rect 147766 322260 147772 322272
rect 147824 322260 147830 322312
rect 88978 322192 88984 322244
rect 89036 322232 89042 322244
rect 217318 322232 217324 322244
rect 89036 322204 217324 322232
rect 89036 322192 89042 322204
rect 217318 322192 217324 322204
rect 217376 322192 217382 322244
rect 105446 321512 105452 321564
rect 105504 321552 105510 321564
rect 133874 321552 133880 321564
rect 105504 321524 133880 321552
rect 105504 321512 105510 321524
rect 133874 321512 133880 321524
rect 133932 321552 133938 321564
rect 135162 321552 135168 321564
rect 133932 321524 135168 321552
rect 133932 321512 133938 321524
rect 135162 321512 135168 321524
rect 135220 321512 135226 321564
rect 67266 320900 67272 320952
rect 67324 320940 67330 320952
rect 207658 320940 207664 320952
rect 67324 320912 207664 320940
rect 67324 320900 67330 320912
rect 207658 320900 207664 320912
rect 207716 320900 207722 320952
rect 65978 320832 65984 320884
rect 66036 320872 66042 320884
rect 112438 320872 112444 320884
rect 66036 320844 112444 320872
rect 66036 320832 66042 320844
rect 112438 320832 112444 320844
rect 112496 320832 112502 320884
rect 135162 320832 135168 320884
rect 135220 320872 135226 320884
rect 349798 320872 349804 320884
rect 135220 320844 349804 320872
rect 135220 320832 135226 320844
rect 349798 320832 349804 320844
rect 349856 320832 349862 320884
rect 100018 320084 100024 320136
rect 100076 320124 100082 320136
rect 131298 320124 131304 320136
rect 100076 320096 131304 320124
rect 100076 320084 100082 320096
rect 131298 320084 131304 320096
rect 131356 320124 131362 320136
rect 131666 320124 131672 320136
rect 131356 320096 131672 320124
rect 131356 320084 131362 320096
rect 131666 320084 131672 320096
rect 131724 320084 131730 320136
rect 75178 319472 75184 319524
rect 75236 319512 75242 319524
rect 115382 319512 115388 319524
rect 75236 319484 115388 319512
rect 75236 319472 75242 319484
rect 115382 319472 115388 319484
rect 115440 319472 115446 319524
rect 69198 319404 69204 319456
rect 69256 319444 69262 319456
rect 121638 319444 121644 319456
rect 69256 319416 121644 319444
rect 69256 319404 69262 319416
rect 121638 319404 121644 319416
rect 121696 319404 121702 319456
rect 106090 318112 106096 318164
rect 106148 318152 106154 318164
rect 113818 318152 113824 318164
rect 106148 318124 113824 318152
rect 106148 318112 106154 318124
rect 113818 318112 113824 318124
rect 113876 318112 113882 318164
rect 83458 318044 83464 318096
rect 83516 318084 83522 318096
rect 351914 318084 351920 318096
rect 83516 318056 351920 318084
rect 83516 318044 83522 318056
rect 351914 318044 351920 318056
rect 351972 318044 351978 318096
rect 59998 316752 60004 316804
rect 60056 316792 60062 316804
rect 128630 316792 128636 316804
rect 60056 316764 128636 316792
rect 60056 316752 60062 316764
rect 128630 316752 128636 316764
rect 128688 316752 128694 316804
rect 84286 316684 84292 316736
rect 84344 316724 84350 316736
rect 113910 316724 113916 316736
rect 84344 316696 113916 316724
rect 84344 316684 84350 316696
rect 113910 316684 113916 316696
rect 113968 316684 113974 316736
rect 115198 316684 115204 316736
rect 115256 316724 115262 316736
rect 204990 316724 204996 316736
rect 115256 316696 204996 316724
rect 115256 316684 115262 316696
rect 204990 316684 204996 316696
rect 205048 316684 205054 316736
rect 91922 315936 91928 315988
rect 91980 315976 91986 315988
rect 124398 315976 124404 315988
rect 91980 315948 124404 315976
rect 91980 315936 91986 315948
rect 124398 315936 124404 315948
rect 124456 315936 124462 315988
rect 73154 315256 73160 315308
rect 73212 315296 73218 315308
rect 116026 315296 116032 315308
rect 73212 315268 116032 315296
rect 73212 315256 73218 315268
rect 116026 315256 116032 315268
rect 116084 315256 116090 315308
rect 69106 313896 69112 313948
rect 69164 313936 69170 313948
rect 282270 313936 282276 313948
rect 69164 313908 282276 313936
rect 69164 313896 69170 313908
rect 282270 313896 282276 313908
rect 282328 313896 282334 313948
rect 69014 313284 69020 313336
rect 69072 313324 69078 313336
rect 122558 313324 122564 313336
rect 69072 313296 122564 313324
rect 69072 313284 69078 313296
rect 122558 313284 122564 313296
rect 122616 313324 122622 313336
rect 395338 313324 395344 313336
rect 122616 313296 395344 313324
rect 122616 313284 122622 313296
rect 395338 313284 395344 313296
rect 395396 313284 395402 313336
rect 102226 313216 102232 313268
rect 102284 313256 102290 313268
rect 127250 313256 127256 313268
rect 102284 313228 127256 313256
rect 102284 313216 102290 313228
rect 127250 313216 127256 313228
rect 127308 313216 127314 313268
rect 71130 312536 71136 312588
rect 71188 312576 71194 312588
rect 129826 312576 129832 312588
rect 71188 312548 129832 312576
rect 71188 312536 71194 312548
rect 129826 312536 129832 312548
rect 129884 312576 129890 312588
rect 410518 312576 410524 312588
rect 129884 312548 410524 312576
rect 129884 312536 129890 312548
rect 410518 312536 410524 312548
rect 410576 312536 410582 312588
rect 81434 311856 81440 311908
rect 81492 311896 81498 311908
rect 356054 311896 356060 311908
rect 81492 311868 356060 311896
rect 81492 311856 81498 311868
rect 356054 311856 356060 311868
rect 356112 311856 356118 311908
rect 102870 311788 102876 311840
rect 102928 311828 102934 311840
rect 135438 311828 135444 311840
rect 102928 311800 135444 311828
rect 102928 311788 102934 311800
rect 135438 311788 135444 311800
rect 135496 311828 135502 311840
rect 136542 311828 136548 311840
rect 135496 311800 136548 311828
rect 135496 311788 135502 311800
rect 136542 311788 136548 311800
rect 136600 311788 136606 311840
rect 117958 311720 117964 311772
rect 118016 311760 118022 311772
rect 125502 311760 125508 311772
rect 118016 311732 125508 311760
rect 118016 311720 118022 311732
rect 125502 311720 125508 311732
rect 125560 311720 125566 311772
rect 79318 311312 79324 311364
rect 79376 311352 79382 311364
rect 120166 311352 120172 311364
rect 79376 311324 120172 311352
rect 79376 311312 79382 311324
rect 120166 311312 120172 311324
rect 120224 311312 120230 311364
rect 91094 311244 91100 311296
rect 91152 311284 91158 311296
rect 121546 311284 121552 311296
rect 91152 311256 121552 311284
rect 91152 311244 91158 311256
rect 121546 311244 121552 311256
rect 121604 311284 121610 311296
rect 159358 311284 159364 311296
rect 121604 311256 159364 311284
rect 121604 311244 121610 311256
rect 159358 311244 159364 311256
rect 159416 311244 159422 311296
rect 70302 311176 70308 311228
rect 70360 311216 70366 311228
rect 104158 311216 104164 311228
rect 70360 311188 104164 311216
rect 70360 311176 70366 311188
rect 104158 311176 104164 311188
rect 104216 311176 104222 311228
rect 136542 311176 136548 311228
rect 136600 311216 136606 311228
rect 273898 311216 273904 311228
rect 136600 311188 273904 311216
rect 136600 311176 136606 311188
rect 273898 311176 273904 311188
rect 273956 311176 273962 311228
rect 114462 311108 114468 311160
rect 114520 311148 114526 311160
rect 141418 311148 141424 311160
rect 114520 311120 141424 311148
rect 114520 311108 114526 311120
rect 141418 311108 141424 311120
rect 141476 311148 141482 311160
rect 464338 311148 464344 311160
rect 141476 311120 464344 311148
rect 141476 311108 141482 311120
rect 464338 311108 464344 311120
rect 464396 311108 464402 311160
rect 539502 311108 539508 311160
rect 539560 311148 539566 311160
rect 580166 311148 580172 311160
rect 539560 311120 580172 311148
rect 539560 311108 539566 311120
rect 580166 311108 580172 311120
rect 580224 311108 580230 311160
rect 124306 310496 124312 310548
rect 124364 310536 124370 310548
rect 125502 310536 125508 310548
rect 124364 310508 125508 310536
rect 124364 310496 124370 310508
rect 125502 310496 125508 310508
rect 125560 310536 125566 310548
rect 538214 310536 538220 310548
rect 125560 310508 538220 310536
rect 125560 310496 125566 310508
rect 538214 310496 538220 310508
rect 538272 310536 538278 310548
rect 539502 310536 539508 310548
rect 538272 310508 539508 310536
rect 538272 310496 538278 310508
rect 539502 310496 539508 310508
rect 539560 310496 539566 310548
rect 3418 310428 3424 310480
rect 3476 310468 3482 310480
rect 48130 310468 48136 310480
rect 3476 310440 48136 310468
rect 3476 310428 3482 310440
rect 48130 310428 48136 310440
rect 48188 310428 48194 310480
rect 80054 309884 80060 309936
rect 80112 309924 80118 309936
rect 91094 309924 91100 309936
rect 80112 309896 91100 309924
rect 80112 309884 80118 309896
rect 91094 309884 91100 309896
rect 91152 309884 91158 309936
rect 107654 309884 107660 309936
rect 107712 309924 107718 309936
rect 134518 309924 134524 309936
rect 107712 309896 134524 309924
rect 107712 309884 107718 309896
rect 134518 309884 134524 309896
rect 134576 309924 134582 309936
rect 135162 309924 135168 309936
rect 134576 309896 135168 309924
rect 134576 309884 134582 309896
rect 135162 309884 135168 309896
rect 135220 309884 135226 309936
rect 76558 309816 76564 309868
rect 76616 309856 76622 309868
rect 192478 309856 192484 309868
rect 76616 309828 192484 309856
rect 76616 309816 76622 309828
rect 192478 309816 192484 309828
rect 192536 309816 192542 309868
rect 48130 309748 48136 309800
rect 48188 309788 48194 309800
rect 116670 309788 116676 309800
rect 48188 309760 116676 309788
rect 48188 309748 48194 309760
rect 116670 309748 116676 309760
rect 116728 309748 116734 309800
rect 135162 309748 135168 309800
rect 135220 309788 135226 309800
rect 521654 309788 521660 309800
rect 135220 309760 521660 309788
rect 135220 309748 135226 309760
rect 521654 309748 521660 309760
rect 521712 309748 521718 309800
rect 75178 309204 75184 309256
rect 75236 309244 75242 309256
rect 228450 309244 228456 309256
rect 75236 309216 228456 309244
rect 75236 309204 75242 309216
rect 228450 309204 228456 309216
rect 228508 309204 228514 309256
rect 89714 309136 89720 309188
rect 89772 309176 89778 309188
rect 304258 309176 304264 309188
rect 89772 309148 304264 309176
rect 89772 309136 89778 309148
rect 304258 309136 304264 309148
rect 304316 309136 304322 309188
rect 108298 309068 108304 309120
rect 108356 309108 108362 309120
rect 142154 309108 142160 309120
rect 108356 309080 142160 309108
rect 108356 309068 108362 309080
rect 142154 309068 142160 309080
rect 142212 309108 142218 309120
rect 143442 309108 143448 309120
rect 142212 309080 143448 309108
rect 142212 309068 142218 309080
rect 143442 309068 143448 309080
rect 143500 309068 143506 309120
rect 75914 308456 75920 308508
rect 75972 308496 75978 308508
rect 216030 308496 216036 308508
rect 75972 308468 216036 308496
rect 75972 308456 75978 308468
rect 216030 308456 216036 308468
rect 216088 308456 216094 308508
rect 84378 308388 84384 308440
rect 84436 308428 84442 308440
rect 114462 308428 114468 308440
rect 84436 308400 114468 308428
rect 84436 308388 84442 308400
rect 114462 308388 114468 308400
rect 114520 308388 114526 308440
rect 143442 308388 143448 308440
rect 143500 308428 143506 308440
rect 475378 308428 475384 308440
rect 143500 308400 475384 308428
rect 143500 308388 143506 308400
rect 475378 308388 475384 308400
rect 475436 308388 475442 308440
rect 102042 307776 102048 307828
rect 102100 307816 102106 307828
rect 103698 307816 103704 307828
rect 102100 307788 103704 307816
rect 102100 307776 102106 307788
rect 103698 307776 103704 307788
rect 103756 307816 103762 307828
rect 467098 307816 467104 307828
rect 103756 307788 467104 307816
rect 103756 307776 103762 307788
rect 467098 307776 467104 307788
rect 467156 307776 467162 307828
rect 93670 307028 93676 307080
rect 93728 307068 93734 307080
rect 279418 307068 279424 307080
rect 93728 307040 279424 307068
rect 93728 307028 93734 307040
rect 279418 307028 279424 307040
rect 279476 307028 279482 307080
rect 86954 306484 86960 306536
rect 87012 306524 87018 306536
rect 213270 306524 213276 306536
rect 87012 306496 213276 306524
rect 87012 306484 87018 306496
rect 213270 306484 213276 306496
rect 213328 306484 213334 306536
rect 85574 306416 85580 306468
rect 85632 306456 85638 306468
rect 240778 306456 240784 306468
rect 85632 306428 240784 306456
rect 85632 306416 85638 306428
rect 240778 306416 240784 306428
rect 240836 306416 240842 306468
rect 106274 306348 106280 306400
rect 106332 306388 106338 306400
rect 118878 306388 118884 306400
rect 106332 306360 118884 306388
rect 106332 306348 106338 306360
rect 118878 306348 118884 306360
rect 118936 306388 118942 306400
rect 514754 306388 514760 306400
rect 118936 306360 514760 306388
rect 118936 306348 118942 306360
rect 514754 306348 514760 306360
rect 514812 306348 514818 306400
rect 3418 306212 3424 306264
rect 3476 306252 3482 306264
rect 7558 306252 7564 306264
rect 3476 306224 7564 306252
rect 3476 306212 3482 306224
rect 7558 306212 7564 306224
rect 7616 306212 7622 306264
rect 59078 305736 59084 305788
rect 59136 305776 59142 305788
rect 123662 305776 123668 305788
rect 59136 305748 123668 305776
rect 59136 305736 59142 305748
rect 123662 305736 123668 305748
rect 123720 305736 123726 305788
rect 90358 305668 90364 305720
rect 90416 305708 90422 305720
rect 275278 305708 275284 305720
rect 90416 305680 275284 305708
rect 90416 305668 90422 305680
rect 275278 305668 275284 305680
rect 275336 305668 275342 305720
rect 93118 305600 93124 305652
rect 93176 305640 93182 305652
rect 294598 305640 294604 305652
rect 93176 305612 294604 305640
rect 93176 305600 93182 305612
rect 294598 305600 294604 305612
rect 294656 305600 294662 305652
rect 81894 305056 81900 305108
rect 81952 305096 81958 305108
rect 221458 305096 221464 305108
rect 81952 305068 221464 305096
rect 81952 305056 81958 305068
rect 221458 305056 221464 305068
rect 221516 305056 221522 305108
rect 367738 305028 367744 305040
rect 78600 305000 367744 305028
rect 49418 304920 49424 304972
rect 49476 304960 49482 304972
rect 77386 304960 77392 304972
rect 49476 304932 77392 304960
rect 49476 304920 49482 304932
rect 77386 304920 77392 304932
rect 77444 304960 77450 304972
rect 78600 304960 78628 305000
rect 367738 304988 367744 305000
rect 367796 304988 367802 305040
rect 77444 304932 78628 304960
rect 77444 304920 77450 304932
rect 107562 304308 107568 304360
rect 107620 304348 107626 304360
rect 127618 304348 127624 304360
rect 107620 304320 127624 304348
rect 107620 304308 107626 304320
rect 127618 304308 127624 304320
rect 127676 304308 127682 304360
rect 60642 304240 60648 304292
rect 60700 304280 60706 304292
rect 124858 304280 124864 304292
rect 60700 304252 124864 304280
rect 60700 304240 60706 304252
rect 124858 304240 124864 304252
rect 124916 304240 124922 304292
rect 146938 303900 146944 303952
rect 146996 303940 147002 303952
rect 196710 303940 196716 303952
rect 146996 303912 196716 303940
rect 146996 303900 147002 303912
rect 196710 303900 196716 303912
rect 196768 303900 196774 303952
rect 233878 303872 233884 303884
rect 95068 303844 233884 303872
rect 95068 303816 95096 303844
rect 233878 303832 233884 303844
rect 233936 303832 233942 303884
rect 94498 303764 94504 303816
rect 94556 303804 94562 303816
rect 95050 303804 95056 303816
rect 94556 303776 95056 303804
rect 94556 303764 94562 303776
rect 95050 303764 95056 303776
rect 95108 303764 95114 303816
rect 96614 303764 96620 303816
rect 96672 303804 96678 303816
rect 315298 303804 315304 303816
rect 96672 303776 315304 303804
rect 96672 303764 96678 303776
rect 315298 303764 315304 303776
rect 315356 303764 315362 303816
rect 86310 303696 86316 303748
rect 86368 303736 86374 303748
rect 318058 303736 318064 303748
rect 86368 303708 318064 303736
rect 86368 303696 86374 303708
rect 318058 303696 318064 303708
rect 318116 303696 318122 303748
rect 482278 303668 482284 303680
rect 67560 303640 482284 303668
rect 56502 303560 56508 303612
rect 56560 303600 56566 303612
rect 66898 303600 66904 303612
rect 56560 303572 66904 303600
rect 56560 303560 56566 303572
rect 66898 303560 66904 303572
rect 66956 303600 66962 303612
rect 67560 303600 67588 303640
rect 482278 303628 482284 303640
rect 482336 303628 482342 303680
rect 66956 303572 67588 303600
rect 66956 303560 66962 303572
rect 93946 302880 93952 302932
rect 94004 302920 94010 302932
rect 122834 302920 122840 302932
rect 94004 302892 122840 302920
rect 94004 302880 94010 302892
rect 122834 302880 122840 302892
rect 122892 302880 122898 302932
rect 90266 302472 90272 302524
rect 90324 302512 90330 302524
rect 135898 302512 135904 302524
rect 90324 302484 135904 302512
rect 90324 302472 90330 302484
rect 135898 302472 135904 302484
rect 135956 302472 135962 302524
rect 66162 302404 66168 302456
rect 66220 302444 66226 302456
rect 169018 302444 169024 302456
rect 66220 302416 169024 302444
rect 66220 302404 66226 302416
rect 169018 302404 169024 302416
rect 169076 302404 169082 302456
rect 115934 302336 115940 302388
rect 115992 302376 115998 302388
rect 116670 302376 116676 302388
rect 115992 302348 116676 302376
rect 115992 302336 115998 302348
rect 116670 302336 116676 302348
rect 116728 302376 116734 302388
rect 232590 302376 232596 302388
rect 116728 302348 232596 302376
rect 116728 302336 116734 302348
rect 232590 302336 232596 302348
rect 232648 302336 232654 302388
rect 75914 302268 75920 302320
rect 75972 302308 75978 302320
rect 193858 302308 193864 302320
rect 75972 302280 193864 302308
rect 75972 302268 75978 302280
rect 193858 302268 193864 302280
rect 193916 302268 193922 302320
rect 71774 302200 71780 302252
rect 71832 302240 71838 302252
rect 325694 302240 325700 302252
rect 71832 302212 325700 302240
rect 71832 302200 71838 302212
rect 325694 302200 325700 302212
rect 325752 302200 325758 302252
rect 105630 301520 105636 301572
rect 105688 301560 105694 301572
rect 105688 301532 142154 301560
rect 105688 301520 105694 301532
rect 43898 301452 43904 301504
rect 43956 301492 43962 301504
rect 124398 301492 124404 301504
rect 43956 301464 124404 301492
rect 43956 301452 43962 301464
rect 124398 301452 124404 301464
rect 124456 301452 124462 301504
rect 142126 301492 142154 301532
rect 145098 301492 145104 301504
rect 142126 301464 145104 301492
rect 145098 301452 145104 301464
rect 145156 301492 145162 301504
rect 238018 301492 238024 301504
rect 145156 301464 238024 301492
rect 145156 301452 145162 301464
rect 238018 301452 238024 301464
rect 238076 301452 238082 301504
rect 104894 301384 104900 301436
rect 104952 301424 104958 301436
rect 106182 301424 106188 301436
rect 104952 301396 106188 301424
rect 104952 301384 104958 301396
rect 106182 301384 106188 301396
rect 106240 301384 106246 301436
rect 106182 301044 106188 301096
rect 106240 301084 106246 301096
rect 187050 301084 187056 301096
rect 106240 301056 187056 301084
rect 106240 301044 106246 301056
rect 187050 301044 187056 301056
rect 187108 301044 187114 301096
rect 79318 300976 79324 301028
rect 79376 301016 79382 301028
rect 214650 301016 214656 301028
rect 79376 300988 214656 301016
rect 79376 300976 79382 300988
rect 214650 300976 214656 300988
rect 214708 300976 214714 301028
rect 88334 300908 88340 300960
rect 88392 300948 88398 300960
rect 347774 300948 347780 300960
rect 88392 300920 347780 300948
rect 88392 300908 88398 300920
rect 347774 300908 347780 300920
rect 347832 300908 347838 300960
rect 88426 300840 88432 300892
rect 88484 300880 88490 300892
rect 350534 300880 350540 300892
rect 88484 300852 350540 300880
rect 88484 300840 88490 300852
rect 350534 300840 350540 300852
rect 350592 300840 350598 300892
rect 226978 300200 226984 300212
rect 74506 300172 226984 300200
rect 59262 300092 59268 300144
rect 59320 300132 59326 300144
rect 70302 300132 70308 300144
rect 59320 300104 70308 300132
rect 59320 300092 59326 300104
rect 70302 300092 70308 300104
rect 70360 300132 70366 300144
rect 74506 300132 74534 300172
rect 226978 300160 226984 300172
rect 227036 300160 227042 300212
rect 70360 300104 74534 300132
rect 70360 300092 70366 300104
rect 87598 300092 87604 300144
rect 87656 300132 87662 300144
rect 344278 300132 344284 300144
rect 87656 300104 344284 300132
rect 87656 300092 87662 300104
rect 344278 300092 344284 300104
rect 344336 300092 344342 300144
rect 94038 300024 94044 300076
rect 94096 300064 94102 300076
rect 95142 300064 95148 300076
rect 94096 300036 95148 300064
rect 94096 300024 94102 300036
rect 95142 300024 95148 300036
rect 95200 300024 95206 300076
rect 113910 299684 113916 299736
rect 113968 299724 113974 299736
rect 130378 299724 130384 299736
rect 113968 299696 130384 299724
rect 113968 299684 113974 299696
rect 130378 299684 130384 299696
rect 130436 299684 130442 299736
rect 95142 299616 95148 299668
rect 95200 299656 95206 299668
rect 166258 299656 166264 299668
rect 95200 299628 166264 299656
rect 95200 299616 95206 299628
rect 166258 299616 166264 299628
rect 166316 299616 166322 299668
rect 110414 299548 110420 299600
rect 110472 299588 110478 299600
rect 266354 299588 266360 299600
rect 110472 299560 266360 299588
rect 110472 299548 110478 299560
rect 266354 299548 266360 299560
rect 266412 299548 266418 299600
rect 109034 299480 109040 299532
rect 109092 299520 109098 299532
rect 331858 299520 331864 299532
rect 109092 299492 331864 299520
rect 109092 299480 109098 299492
rect 331858 299480 331864 299492
rect 331916 299480 331922 299532
rect 74442 298732 74448 298784
rect 74500 298772 74506 298784
rect 128538 298772 128544 298784
rect 74500 298744 128544 298772
rect 74500 298732 74506 298744
rect 128538 298732 128544 298744
rect 128596 298772 128602 298784
rect 195330 298772 195336 298784
rect 128596 298744 195336 298772
rect 128596 298732 128602 298744
rect 195330 298732 195336 298744
rect 195388 298732 195394 298784
rect 419534 298732 419540 298784
rect 419592 298772 419598 298784
rect 580258 298772 580264 298784
rect 419592 298744 580264 298772
rect 419592 298732 419598 298744
rect 580258 298732 580264 298744
rect 580316 298732 580322 298784
rect 83550 298392 83556 298444
rect 83608 298432 83614 298444
rect 147030 298432 147036 298444
rect 83608 298404 147036 298432
rect 83608 298392 83614 298404
rect 147030 298392 147036 298404
rect 147088 298392 147094 298444
rect 117682 298324 117688 298376
rect 117740 298364 117746 298376
rect 191190 298364 191196 298376
rect 117740 298336 191196 298364
rect 117740 298324 117746 298336
rect 191190 298324 191196 298336
rect 191248 298324 191254 298376
rect 67542 298256 67548 298308
rect 67600 298296 67606 298308
rect 220078 298296 220084 298308
rect 67600 298268 220084 298296
rect 67600 298256 67606 298268
rect 220078 298256 220084 298268
rect 220136 298256 220142 298308
rect 93210 298188 93216 298240
rect 93268 298228 93274 298240
rect 246298 298228 246304 298240
rect 93268 298200 246304 298228
rect 93268 298188 93274 298200
rect 246298 298188 246304 298200
rect 246356 298188 246362 298240
rect 102870 298120 102876 298172
rect 102928 298160 102934 298172
rect 276014 298160 276020 298172
rect 102928 298132 276020 298160
rect 102928 298120 102934 298132
rect 276014 298120 276020 298132
rect 276072 298120 276078 298172
rect 91922 297032 91928 297084
rect 91980 297072 91986 297084
rect 133138 297072 133144 297084
rect 91980 297044 133144 297072
rect 91980 297032 91986 297044
rect 133138 297032 133144 297044
rect 133196 297032 133202 297084
rect 98638 296964 98644 297016
rect 98696 297004 98702 297016
rect 160830 297004 160836 297016
rect 98696 296976 160836 297004
rect 98696 296964 98702 296976
rect 160830 296964 160836 296976
rect 160888 296964 160894 297016
rect 67634 296896 67640 296948
rect 67692 296936 67698 296948
rect 224310 296936 224316 296948
rect 67692 296908 224316 296936
rect 67692 296896 67698 296908
rect 224310 296896 224316 296908
rect 224368 296896 224374 296948
rect 82906 296828 82912 296880
rect 82964 296868 82970 296880
rect 249794 296868 249800 296880
rect 82964 296840 249800 296868
rect 82964 296828 82970 296840
rect 249794 296828 249800 296840
rect 249852 296828 249858 296880
rect 75178 296760 75184 296812
rect 75236 296800 75242 296812
rect 251818 296800 251824 296812
rect 75236 296772 251824 296800
rect 75236 296760 75242 296772
rect 251818 296760 251824 296772
rect 251876 296760 251882 296812
rect 113450 296692 113456 296744
rect 113508 296732 113514 296744
rect 113818 296732 113824 296744
rect 113508 296704 113824 296732
rect 113508 296692 113514 296704
rect 113818 296692 113824 296704
rect 113876 296732 113882 296744
rect 378778 296732 378784 296744
rect 113876 296704 378784 296732
rect 113876 296692 113882 296704
rect 378778 296692 378784 296704
rect 378836 296692 378842 296744
rect 69106 295944 69112 295996
rect 69164 295984 69170 295996
rect 94498 295984 94504 295996
rect 69164 295956 94504 295984
rect 69164 295944 69170 295956
rect 94498 295944 94504 295956
rect 94556 295944 94562 295996
rect 92566 295672 92572 295724
rect 92624 295712 92630 295724
rect 93762 295712 93768 295724
rect 92624 295684 93768 295712
rect 92624 295672 92630 295684
rect 93762 295672 93768 295684
rect 93820 295712 93826 295724
rect 125686 295712 125692 295724
rect 93820 295684 125692 295712
rect 93820 295672 93826 295684
rect 125686 295672 125692 295684
rect 125744 295672 125750 295724
rect 99650 295604 99656 295656
rect 99708 295644 99714 295656
rect 144178 295644 144184 295656
rect 99708 295616 144184 295644
rect 99708 295604 99714 295616
rect 144178 295604 144184 295616
rect 144236 295604 144242 295656
rect 88058 295536 88064 295588
rect 88116 295576 88122 295588
rect 155218 295576 155224 295588
rect 88116 295548 155224 295576
rect 88116 295536 88122 295548
rect 155218 295536 155224 295548
rect 155276 295536 155282 295588
rect 74534 295468 74540 295520
rect 74592 295508 74598 295520
rect 225598 295508 225604 295520
rect 74592 295480 225604 295508
rect 74592 295468 74598 295480
rect 225598 295468 225604 295480
rect 225656 295468 225662 295520
rect 69842 295400 69848 295452
rect 69900 295440 69906 295452
rect 244918 295440 244924 295452
rect 69900 295412 244924 295440
rect 69900 295400 69906 295412
rect 244918 295400 244924 295412
rect 244976 295400 244982 295452
rect 106734 295332 106740 295384
rect 106792 295372 106798 295384
rect 333974 295372 333980 295384
rect 106792 295344 333980 295372
rect 106792 295332 106798 295344
rect 333974 295332 333980 295344
rect 334032 295332 334038 295384
rect 70026 295196 70032 295248
rect 70084 295236 70090 295248
rect 75086 295236 75092 295248
rect 70084 295208 75092 295236
rect 70084 295196 70090 295208
rect 75086 295196 75092 295208
rect 75144 295196 75150 295248
rect 99006 294720 99012 294772
rect 99064 294760 99070 294772
rect 113174 294760 113180 294772
rect 99064 294732 113180 294760
rect 99064 294720 99070 294732
rect 113174 294720 113180 294732
rect 113232 294720 113238 294772
rect 84194 294652 84200 294704
rect 84252 294692 84258 294704
rect 113910 294692 113916 294704
rect 84252 294664 113916 294692
rect 84252 294652 84258 294664
rect 113910 294652 113916 294664
rect 113968 294652 113974 294704
rect 119614 294652 119620 294704
rect 119672 294692 119678 294704
rect 146938 294692 146944 294704
rect 119672 294664 146944 294692
rect 119672 294652 119678 294664
rect 146938 294652 146944 294664
rect 146996 294652 147002 294704
rect 511994 294652 512000 294704
rect 512052 294692 512058 294704
rect 580902 294692 580908 294704
rect 512052 294664 580908 294692
rect 512052 294652 512058 294664
rect 580902 294652 580908 294664
rect 580960 294652 580966 294704
rect 109954 294584 109960 294636
rect 110012 294624 110018 294636
rect 152090 294624 152096 294636
rect 110012 294596 152096 294624
rect 110012 294584 110018 294596
rect 152090 294584 152096 294596
rect 152148 294624 152154 294636
rect 525794 294624 525800 294636
rect 152148 294596 525800 294624
rect 152148 294584 152154 294596
rect 525794 294584 525800 294596
rect 525852 294584 525858 294636
rect 71314 294380 71320 294432
rect 71372 294420 71378 294432
rect 72418 294420 72424 294432
rect 71372 294392 72424 294420
rect 71372 294380 71378 294392
rect 72418 294380 72424 294392
rect 72476 294380 72482 294432
rect 73154 294312 73160 294364
rect 73212 294352 73218 294364
rect 73614 294352 73620 294364
rect 73212 294324 73620 294352
rect 73212 294312 73218 294324
rect 73614 294312 73620 294324
rect 73672 294312 73678 294364
rect 77294 294312 77300 294364
rect 77352 294352 77358 294364
rect 78030 294352 78036 294364
rect 77352 294324 78036 294352
rect 77352 294312 77358 294324
rect 78030 294312 78036 294324
rect 78088 294312 78094 294364
rect 84286 294312 84292 294364
rect 84344 294352 84350 294364
rect 85206 294352 85212 294364
rect 84344 294324 85212 294352
rect 84344 294312 84350 294324
rect 85206 294312 85212 294324
rect 85264 294312 85270 294364
rect 88334 294312 88340 294364
rect 88392 294352 88398 294364
rect 89070 294352 89076 294364
rect 88392 294324 89076 294352
rect 88392 294312 88398 294324
rect 89070 294312 89076 294324
rect 89128 294312 89134 294364
rect 93946 294312 93952 294364
rect 94004 294352 94010 294364
rect 94774 294352 94780 294364
rect 94004 294324 94780 294352
rect 94004 294312 94010 294324
rect 94774 294312 94780 294324
rect 94832 294312 94838 294364
rect 72602 294244 72608 294296
rect 72660 294284 72666 294296
rect 74442 294284 74448 294296
rect 72660 294256 74448 294284
rect 72660 294244 72666 294256
rect 74442 294244 74448 294256
rect 74500 294244 74506 294296
rect 115106 294244 115112 294296
rect 115164 294284 115170 294296
rect 115382 294284 115388 294296
rect 115164 294256 115388 294284
rect 115164 294244 115170 294256
rect 115382 294244 115388 294256
rect 115440 294284 115446 294296
rect 123570 294284 123576 294296
rect 115440 294256 123576 294284
rect 115440 294244 115446 294256
rect 123570 294244 123576 294256
rect 123628 294244 123634 294296
rect 103514 294176 103520 294228
rect 103572 294216 103578 294228
rect 117222 294216 117228 294228
rect 103572 294188 117228 294216
rect 103572 294176 103578 294188
rect 117222 294176 117228 294188
rect 117280 294176 117286 294228
rect 115290 294108 115296 294160
rect 115348 294148 115354 294160
rect 123754 294148 123760 294160
rect 115348 294120 123760 294148
rect 115348 294108 115354 294120
rect 123754 294108 123760 294120
rect 123812 294108 123818 294160
rect 57790 294040 57796 294092
rect 57848 294080 57854 294092
rect 79042 294080 79048 294092
rect 57848 294052 79048 294080
rect 57848 294040 57854 294052
rect 79042 294040 79048 294052
rect 79100 294040 79106 294092
rect 80974 294040 80980 294092
rect 81032 294080 81038 294092
rect 117130 294080 117136 294092
rect 81032 294052 117136 294080
rect 81032 294040 81038 294052
rect 117130 294040 117136 294052
rect 117188 294040 117194 294092
rect 44082 293972 44088 294024
rect 44140 294012 44146 294024
rect 96430 294012 96436 294024
rect 44140 293984 96436 294012
rect 44140 293972 44146 293984
rect 96430 293972 96436 293984
rect 96488 293972 96494 294024
rect 113818 293972 113824 294024
rect 113876 294012 113882 294024
rect 357526 294012 357532 294024
rect 113876 293984 357532 294012
rect 113876 293972 113882 293984
rect 357526 293972 357532 293984
rect 357584 293972 357590 294024
rect 3050 293904 3056 293956
rect 3108 293944 3114 293956
rect 14458 293944 14464 293956
rect 3108 293916 14464 293944
rect 3108 293904 3114 293916
rect 14458 293904 14464 293916
rect 14516 293904 14522 293956
rect 113082 293360 113088 293412
rect 113140 293400 113146 293412
rect 126238 293400 126244 293412
rect 113140 293372 126244 293400
rect 113140 293360 113174 293372
rect 126238 293360 126244 293372
rect 126296 293360 126302 293412
rect 77110 293292 77116 293344
rect 77168 293332 77174 293344
rect 113146 293332 113174 293360
rect 77168 293304 113174 293332
rect 77168 293292 77174 293304
rect 116578 293292 116584 293344
rect 116636 293332 116642 293344
rect 131114 293332 131120 293344
rect 116636 293304 131120 293332
rect 116636 293292 116642 293304
rect 131114 293292 131120 293304
rect 131172 293292 131178 293344
rect 21358 293224 21364 293276
rect 21416 293264 21422 293276
rect 53190 293264 53196 293276
rect 21416 293236 53196 293264
rect 21416 293224 21422 293236
rect 53190 293224 53196 293236
rect 53248 293264 53254 293276
rect 97074 293264 97080 293276
rect 53248 293236 97080 293264
rect 53248 293224 53254 293236
rect 97074 293224 97080 293236
rect 97132 293224 97138 293276
rect 117222 293224 117228 293276
rect 117280 293264 117286 293276
rect 311158 293264 311164 293276
rect 117280 293236 311164 293264
rect 117280 293224 117286 293236
rect 311158 293224 311164 293236
rect 311216 293224 311222 293276
rect 93854 292680 93860 292732
rect 93912 292720 93918 292732
rect 142798 292720 142804 292732
rect 93912 292692 142804 292720
rect 93912 292680 93918 292692
rect 142798 292680 142804 292692
rect 142856 292680 142862 292732
rect 112530 292612 112536 292664
rect 112588 292652 112594 292664
rect 220170 292652 220176 292664
rect 112588 292624 220176 292652
rect 112588 292612 112594 292624
rect 220170 292612 220176 292624
rect 220228 292612 220234 292664
rect 102226 292544 102232 292596
rect 102284 292584 102290 292596
rect 229738 292584 229744 292596
rect 102284 292556 229744 292584
rect 102284 292544 102290 292556
rect 229738 292544 229744 292556
rect 229796 292544 229802 292596
rect 118326 292476 118332 292528
rect 118384 292516 118390 292528
rect 119798 292516 119804 292528
rect 118384 292488 119804 292516
rect 118384 292476 118390 292488
rect 119798 292476 119804 292488
rect 119856 292516 119862 292528
rect 135346 292516 135352 292528
rect 119856 292488 135352 292516
rect 119856 292476 119862 292488
rect 135346 292476 135352 292488
rect 135404 292476 135410 292528
rect 117130 291932 117136 291984
rect 117188 291972 117194 291984
rect 117188 291944 122834 291972
rect 117188 291932 117194 291944
rect 103974 291864 103980 291916
rect 104032 291904 104038 291916
rect 104032 291876 113174 291904
rect 104032 291864 104038 291876
rect 4062 291796 4068 291848
rect 4120 291836 4126 291848
rect 57790 291836 57796 291848
rect 4120 291808 57796 291836
rect 4120 291796 4126 291808
rect 57790 291796 57796 291808
rect 57848 291796 57854 291848
rect 113146 291360 113174 291876
rect 117222 291864 117228 291916
rect 117280 291864 117286 291916
rect 119338 291864 119344 291916
rect 119396 291904 119402 291916
rect 119982 291904 119988 291916
rect 119396 291876 119988 291904
rect 119396 291864 119402 291876
rect 119982 291864 119988 291876
rect 120040 291864 120046 291916
rect 117240 291836 117268 291864
rect 119890 291836 119896 291848
rect 117240 291808 119896 291836
rect 119890 291796 119896 291808
rect 119948 291796 119954 291848
rect 122806 291836 122834 291944
rect 224218 291836 224224 291848
rect 122806 291808 224224 291836
rect 224218 291796 224224 291808
rect 224276 291796 224282 291848
rect 121546 291728 121552 291780
rect 121604 291768 121610 291780
rect 123478 291768 123484 291780
rect 121604 291740 123484 291768
rect 121604 291728 121610 291740
rect 123478 291728 123484 291740
rect 123536 291768 123542 291780
rect 124858 291768 124864 291780
rect 123536 291740 124864 291768
rect 123536 291728 123542 291740
rect 124858 291728 124864 291740
rect 124916 291728 124922 291780
rect 231210 291360 231216 291372
rect 113146 291332 231216 291360
rect 231210 291320 231216 291332
rect 231268 291320 231274 291372
rect 119982 291252 119988 291304
rect 120040 291292 120046 291304
rect 345106 291292 345112 291304
rect 120040 291264 345112 291292
rect 120040 291252 120046 291264
rect 345106 291252 345112 291264
rect 345164 291252 345170 291304
rect 119890 291184 119896 291236
rect 119948 291224 119954 291236
rect 353386 291224 353392 291236
rect 119948 291196 353392 291224
rect 119948 291184 119954 291196
rect 353386 291184 353392 291196
rect 353444 291184 353450 291236
rect 22738 290436 22744 290488
rect 22796 290476 22802 290488
rect 65978 290476 65984 290488
rect 22796 290448 65984 290476
rect 22796 290436 22802 290448
rect 65978 290436 65984 290448
rect 66036 290476 66042 290488
rect 67726 290476 67732 290488
rect 66036 290448 67732 290476
rect 66036 290436 66042 290448
rect 67726 290436 67732 290448
rect 67784 290436 67790 290488
rect 121546 289824 121552 289876
rect 121604 289864 121610 289876
rect 214558 289864 214564 289876
rect 121604 289836 214564 289864
rect 121604 289824 121610 289836
rect 214558 289824 214564 289836
rect 214616 289824 214622 289876
rect 123478 289756 123484 289808
rect 123536 289796 123542 289808
rect 123662 289796 123668 289808
rect 123536 289768 123668 289796
rect 123536 289756 123542 289768
rect 123662 289756 123668 289768
rect 123720 289756 123726 289808
rect 123478 289076 123484 289128
rect 123536 289116 123542 289128
rect 511994 289116 512000 289128
rect 123536 289088 512000 289116
rect 123536 289076 123542 289088
rect 511994 289076 512000 289088
rect 512052 289076 512058 289128
rect 122374 288464 122380 288516
rect 122432 288504 122438 288516
rect 222838 288504 222844 288516
rect 122432 288476 222844 288504
rect 122432 288464 122438 288476
rect 222838 288464 222844 288476
rect 222896 288464 222902 288516
rect 39942 288396 39948 288448
rect 40000 288436 40006 288448
rect 67634 288436 67640 288448
rect 40000 288408 67640 288436
rect 40000 288396 40006 288408
rect 67634 288396 67640 288408
rect 67692 288396 67698 288448
rect 121730 288396 121736 288448
rect 121788 288436 121794 288448
rect 328454 288436 328460 288448
rect 121788 288408 328460 288436
rect 121788 288396 121794 288408
rect 328454 288396 328460 288408
rect 328512 288396 328518 288448
rect 65610 288328 65616 288380
rect 65668 288368 65674 288380
rect 67818 288368 67824 288380
rect 65668 288340 67824 288368
rect 65668 288328 65674 288340
rect 67818 288328 67824 288340
rect 67876 288328 67882 288380
rect 121546 288328 121552 288380
rect 121604 288368 121610 288380
rect 142430 288368 142436 288380
rect 121604 288340 142436 288368
rect 121604 288328 121610 288340
rect 142430 288328 142436 288340
rect 142488 288368 142494 288380
rect 143442 288368 143448 288380
rect 142488 288340 143448 288368
rect 142488 288328 142494 288340
rect 143442 288328 143448 288340
rect 143500 288328 143506 288380
rect 143442 287648 143448 287700
rect 143500 287688 143506 287700
rect 507854 287688 507860 287700
rect 143500 287660 507860 287688
rect 143500 287648 143506 287660
rect 507854 287648 507860 287660
rect 507912 287648 507918 287700
rect 65518 287376 65524 287428
rect 65576 287416 65582 287428
rect 67818 287416 67824 287428
rect 65576 287388 67824 287416
rect 65576 287376 65582 287388
rect 67818 287376 67824 287388
rect 67876 287376 67882 287428
rect 121822 287036 121828 287088
rect 121880 287076 121886 287088
rect 325786 287076 325792 287088
rect 121880 287048 325792 287076
rect 121880 287036 121886 287048
rect 325786 287036 325792 287048
rect 325844 287036 325850 287088
rect 121546 286968 121552 287020
rect 121604 287008 121610 287020
rect 134058 287008 134064 287020
rect 121604 286980 134064 287008
rect 121604 286968 121610 286980
rect 134058 286968 134064 286980
rect 134116 286968 134122 287020
rect 124398 286764 124404 286816
rect 124456 286804 124462 286816
rect 128538 286804 128544 286816
rect 124456 286776 128544 286804
rect 124456 286764 124462 286776
rect 128538 286764 128544 286776
rect 128596 286764 128602 286816
rect 122742 286356 122748 286408
rect 122800 286396 122806 286408
rect 125778 286396 125784 286408
rect 122800 286368 125784 286396
rect 122800 286356 122806 286368
rect 125778 286356 125784 286368
rect 125836 286356 125842 286408
rect 121546 286288 121552 286340
rect 121604 286328 121610 286340
rect 124398 286328 124404 286340
rect 121604 286300 124404 286328
rect 121604 286288 121610 286300
rect 124398 286288 124404 286300
rect 124456 286288 124462 286340
rect 134058 286288 134064 286340
rect 134116 286328 134122 286340
rect 382918 286328 382924 286340
rect 134116 286300 382924 286328
rect 134116 286288 134122 286300
rect 382918 286288 382924 286300
rect 382976 286288 382982 286340
rect 121546 284384 121552 284436
rect 121604 284424 121610 284436
rect 322934 284424 322940 284436
rect 121604 284396 322940 284424
rect 121604 284384 121610 284396
rect 322934 284384 322940 284396
rect 322992 284384 322998 284436
rect 121638 284316 121644 284368
rect 121696 284356 121702 284368
rect 495434 284356 495440 284368
rect 121696 284328 495440 284356
rect 121696 284316 121702 284328
rect 495434 284316 495440 284328
rect 495492 284316 495498 284368
rect 50798 284248 50804 284300
rect 50856 284288 50862 284300
rect 67634 284288 67640 284300
rect 50856 284260 67640 284288
rect 50856 284248 50862 284260
rect 67634 284248 67640 284260
rect 67692 284248 67698 284300
rect 121546 283568 121552 283620
rect 121604 283608 121610 283620
rect 124950 283608 124956 283620
rect 121604 283580 124956 283608
rect 121604 283568 121610 283580
rect 124950 283568 124956 283580
rect 125008 283568 125014 283620
rect 121546 282888 121552 282940
rect 121604 282928 121610 282940
rect 342346 282928 342352 282940
rect 121604 282900 342352 282928
rect 121604 282888 121610 282900
rect 342346 282888 342352 282900
rect 342404 282888 342410 282940
rect 128538 282140 128544 282192
rect 128596 282180 128602 282192
rect 448514 282180 448520 282192
rect 128596 282152 448520 282180
rect 128596 282140 128602 282152
rect 448514 282140 448520 282152
rect 448572 282140 448578 282192
rect 121638 281596 121644 281648
rect 121696 281636 121702 281648
rect 246390 281636 246396 281648
rect 121696 281608 246396 281636
rect 121696 281596 121702 281608
rect 246390 281596 246396 281608
rect 246448 281596 246454 281648
rect 121546 281528 121552 281580
rect 121604 281568 121610 281580
rect 249058 281568 249064 281580
rect 121604 281540 249064 281568
rect 121604 281528 121610 281540
rect 249058 281528 249064 281540
rect 249116 281528 249122 281580
rect 122742 280780 122748 280832
rect 122800 280820 122806 280832
rect 407758 280820 407764 280832
rect 122800 280792 407764 280820
rect 122800 280780 122806 280792
rect 407758 280780 407764 280792
rect 407816 280780 407822 280832
rect 56502 280236 56508 280288
rect 56560 280276 56566 280288
rect 67726 280276 67732 280288
rect 56560 280248 67732 280276
rect 56560 280236 56566 280248
rect 67726 280236 67732 280248
rect 67784 280236 67790 280288
rect 121546 280236 121552 280288
rect 121604 280276 121610 280288
rect 240870 280276 240876 280288
rect 121604 280248 240876 280276
rect 121604 280236 121610 280248
rect 240870 280236 240876 280248
rect 240928 280236 240934 280288
rect 45462 280168 45468 280220
rect 45520 280208 45526 280220
rect 67634 280208 67640 280220
rect 45520 280180 67640 280208
rect 45520 280168 45526 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121638 280168 121644 280220
rect 121696 280208 121702 280220
rect 353294 280208 353300 280220
rect 121696 280180 353300 280208
rect 121696 280168 121702 280180
rect 353294 280168 353300 280180
rect 353352 280168 353358 280220
rect 44174 280100 44180 280152
rect 44232 280140 44238 280152
rect 45370 280140 45376 280152
rect 44232 280112 45376 280140
rect 44232 280100 44238 280112
rect 45370 280100 45376 280112
rect 45428 280140 45434 280152
rect 68002 280140 68008 280152
rect 45428 280112 68008 280140
rect 45428 280100 45434 280112
rect 68002 280100 68008 280112
rect 68060 280100 68066 280152
rect 55122 280032 55128 280084
rect 55180 280072 55186 280084
rect 67634 280072 67640 280084
rect 55180 280044 67640 280072
rect 55180 280032 55186 280044
rect 67634 280032 67640 280044
rect 67692 280032 67698 280084
rect 35158 279420 35164 279472
rect 35216 279460 35222 279472
rect 44174 279460 44180 279472
rect 35216 279432 44180 279460
rect 35216 279420 35222 279432
rect 44174 279420 44180 279432
rect 44232 279420 44238 279472
rect 121546 278808 121552 278860
rect 121604 278848 121610 278860
rect 236638 278848 236644 278860
rect 121604 278820 236644 278848
rect 121604 278808 121610 278820
rect 236638 278808 236644 278820
rect 236696 278808 236702 278860
rect 121638 278740 121644 278792
rect 121696 278780 121702 278792
rect 319438 278780 319444 278792
rect 121696 278752 319444 278780
rect 121696 278740 121702 278752
rect 319438 278740 319444 278752
rect 319496 278740 319502 278792
rect 123754 277992 123760 278044
rect 123812 278032 123818 278044
rect 496814 278032 496820 278044
rect 123812 278004 496820 278032
rect 123812 277992 123818 278004
rect 496814 277992 496820 278004
rect 496872 277992 496878 278044
rect 47946 277448 47952 277500
rect 48004 277488 48010 277500
rect 67634 277488 67640 277500
rect 48004 277460 67640 277488
rect 48004 277448 48010 277460
rect 67634 277448 67640 277460
rect 67692 277448 67698 277500
rect 42702 277380 42708 277432
rect 42760 277420 42766 277432
rect 67726 277420 67732 277432
rect 42760 277392 67732 277420
rect 42760 277380 42766 277392
rect 67726 277380 67732 277392
rect 67784 277380 67790 277432
rect 121546 277380 121552 277432
rect 121604 277420 121610 277432
rect 316678 277420 316684 277432
rect 121604 277392 316684 277420
rect 121604 277380 121610 277392
rect 316678 277380 316684 277392
rect 316736 277380 316742 277432
rect 63310 276088 63316 276140
rect 63368 276128 63374 276140
rect 67634 276128 67640 276140
rect 63368 276100 67640 276128
rect 63368 276088 63374 276100
rect 67634 276088 67640 276100
rect 67692 276088 67698 276140
rect 52178 276020 52184 276072
rect 52236 276060 52242 276072
rect 67726 276060 67732 276072
rect 52236 276032 67732 276060
rect 52236 276020 52242 276032
rect 67726 276020 67732 276032
rect 67784 276020 67790 276072
rect 121546 276020 121552 276072
rect 121604 276060 121610 276072
rect 335354 276060 335360 276072
rect 121604 276032 335360 276060
rect 121604 276020 121610 276032
rect 335354 276020 335360 276032
rect 335412 276020 335418 276072
rect 121638 275952 121644 276004
rect 121696 275992 121702 276004
rect 131114 275992 131120 276004
rect 121696 275964 131120 275992
rect 121696 275952 121702 275964
rect 131114 275952 131120 275964
rect 131172 275952 131178 276004
rect 121730 275340 121736 275392
rect 121788 275380 121794 275392
rect 406378 275380 406384 275392
rect 121788 275352 406384 275380
rect 121788 275340 121794 275352
rect 406378 275340 406384 275352
rect 406436 275340 406442 275392
rect 131114 275272 131120 275324
rect 131172 275312 131178 275324
rect 493318 275312 493324 275324
rect 131172 275284 493324 275312
rect 131172 275272 131178 275284
rect 493318 275272 493324 275284
rect 493376 275272 493382 275324
rect 55122 274728 55128 274780
rect 55180 274768 55186 274780
rect 67726 274768 67732 274780
rect 55180 274740 67732 274768
rect 55180 274728 55186 274740
rect 67726 274728 67732 274740
rect 67784 274728 67790 274780
rect 50798 274660 50804 274712
rect 50856 274700 50862 274712
rect 67634 274700 67640 274712
rect 50856 274672 67640 274700
rect 50856 274660 50862 274672
rect 67634 274660 67640 274672
rect 67692 274660 67698 274712
rect 121546 274660 121552 274712
rect 121604 274700 121610 274712
rect 222930 274700 222936 274712
rect 121604 274672 222936 274700
rect 121604 274660 121610 274672
rect 222930 274660 222936 274672
rect 222988 274660 222994 274712
rect 39758 274592 39764 274644
rect 39816 274632 39822 274644
rect 68002 274632 68008 274644
rect 39816 274604 68008 274632
rect 39816 274592 39822 274604
rect 68002 274592 68008 274604
rect 68060 274592 68066 274644
rect 121546 274524 121552 274576
rect 121604 274564 121610 274576
rect 124306 274564 124312 274576
rect 121604 274536 124312 274564
rect 121604 274524 121610 274536
rect 124306 274524 124312 274536
rect 124364 274524 124370 274576
rect 48130 273232 48136 273284
rect 48188 273272 48194 273284
rect 67634 273272 67640 273284
rect 48188 273244 67640 273272
rect 48188 273232 48194 273244
rect 67634 273232 67640 273244
rect 67692 273232 67698 273284
rect 121546 273232 121552 273284
rect 121604 273272 121610 273284
rect 267734 273272 267740 273284
rect 121604 273244 267740 273272
rect 121604 273232 121610 273244
rect 267734 273232 267740 273244
rect 267792 273232 267798 273284
rect 124950 273164 124956 273216
rect 125008 273204 125014 273216
rect 150434 273204 150440 273216
rect 125008 273176 150440 273204
rect 125008 273164 125014 273176
rect 150434 273164 150440 273176
rect 150492 273164 150498 273216
rect 121546 273096 121552 273148
rect 121604 273136 121610 273148
rect 129826 273136 129832 273148
rect 121604 273108 129832 273136
rect 121604 273096 121610 273108
rect 129826 273096 129832 273108
rect 129884 273096 129890 273148
rect 129826 272552 129832 272604
rect 129884 272592 129890 272604
rect 251910 272592 251916 272604
rect 129884 272564 251916 272592
rect 129884 272552 129890 272564
rect 251910 272552 251916 272564
rect 251968 272552 251974 272604
rect 150434 272484 150440 272536
rect 150492 272524 150498 272536
rect 417418 272524 417424 272536
rect 150492 272496 417424 272524
rect 150492 272484 150498 272496
rect 417418 272484 417424 272496
rect 417476 272484 417482 272536
rect 66070 271940 66076 271992
rect 66128 271980 66134 271992
rect 68186 271980 68192 271992
rect 66128 271952 68192 271980
rect 66128 271940 66134 271952
rect 68186 271940 68192 271952
rect 68244 271940 68250 271992
rect 64506 271872 64512 271924
rect 64564 271912 64570 271924
rect 67634 271912 67640 271924
rect 64564 271884 67640 271912
rect 64564 271872 64570 271884
rect 67634 271872 67640 271884
rect 67692 271872 67698 271924
rect 121546 271872 121552 271924
rect 121604 271912 121610 271924
rect 164878 271912 164884 271924
rect 121604 271884 164884 271912
rect 121604 271872 121610 271884
rect 164878 271872 164884 271884
rect 164936 271872 164942 271924
rect 419442 271872 419448 271924
rect 419500 271912 419506 271924
rect 579798 271912 579804 271924
rect 419500 271884 579804 271912
rect 419500 271872 419506 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 160830 271124 160836 271176
rect 160888 271164 160894 271176
rect 447778 271164 447784 271176
rect 160888 271136 447784 271164
rect 160888 271124 160894 271136
rect 447778 271124 447784 271136
rect 447836 271124 447842 271176
rect 43898 270512 43904 270564
rect 43956 270552 43962 270564
rect 67634 270552 67640 270564
rect 43956 270524 67640 270552
rect 43956 270512 43962 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 121546 270512 121552 270564
rect 121604 270552 121610 270564
rect 233970 270552 233976 270564
rect 121604 270524 233976 270552
rect 121604 270512 121610 270524
rect 233970 270512 233976 270524
rect 234028 270512 234034 270564
rect 46750 269764 46756 269816
rect 46808 269804 46814 269816
rect 68278 269804 68284 269816
rect 46808 269776 68284 269804
rect 46808 269764 46814 269776
rect 68278 269764 68284 269776
rect 68336 269764 68342 269816
rect 49510 269152 49516 269204
rect 49568 269192 49574 269204
rect 67726 269192 67732 269204
rect 49568 269164 67732 269192
rect 49568 269152 49574 269164
rect 67726 269152 67732 269164
rect 67784 269152 67790 269204
rect 121546 269152 121552 269204
rect 121604 269192 121610 269204
rect 231118 269192 231124 269204
rect 121604 269164 231124 269192
rect 121604 269152 121610 269164
rect 231118 269152 231124 269164
rect 231176 269152 231182 269204
rect 45370 269084 45376 269136
rect 45428 269124 45434 269136
rect 67634 269124 67640 269136
rect 45428 269096 67640 269124
rect 45428 269084 45434 269096
rect 67634 269084 67640 269096
rect 67692 269084 67698 269136
rect 121638 269084 121644 269136
rect 121696 269124 121702 269136
rect 252554 269124 252560 269136
rect 121696 269096 252560 269124
rect 121696 269084 121702 269096
rect 252554 269084 252560 269096
rect 252612 269084 252618 269136
rect 53650 269016 53656 269068
rect 53708 269056 53714 269068
rect 54938 269056 54944 269068
rect 53708 269028 54944 269056
rect 53708 269016 53714 269028
rect 54938 269016 54944 269028
rect 54996 269016 55002 269068
rect 129642 268404 129648 268456
rect 129700 268444 129706 268456
rect 139578 268444 139584 268456
rect 129700 268416 139584 268444
rect 129700 268404 129706 268416
rect 139578 268404 139584 268416
rect 139636 268404 139642 268456
rect 119982 268336 119988 268388
rect 120040 268376 120046 268388
rect 434714 268376 434720 268388
rect 120040 268348 434720 268376
rect 120040 268336 120046 268348
rect 434714 268336 434720 268348
rect 434772 268336 434778 268388
rect 61930 267792 61936 267844
rect 61988 267832 61994 267844
rect 67726 267832 67732 267844
rect 61988 267804 67732 267832
rect 61988 267792 61994 267804
rect 67726 267792 67732 267804
rect 67784 267792 67790 267844
rect 121638 267792 121644 267844
rect 121696 267832 121702 267844
rect 129642 267832 129648 267844
rect 121696 267804 129648 267832
rect 121696 267792 121702 267804
rect 129642 267792 129648 267804
rect 129700 267792 129706 267844
rect 67634 267764 67640 267776
rect 52288 267736 67640 267764
rect 39574 267656 39580 267708
rect 39632 267696 39638 267708
rect 51718 267696 51724 267708
rect 39632 267668 51724 267696
rect 39632 267656 39638 267668
rect 51718 267656 51724 267668
rect 51776 267696 51782 267708
rect 52288 267696 52316 267736
rect 67634 267724 67640 267736
rect 67692 267724 67698 267776
rect 121546 267724 121552 267776
rect 121604 267764 121610 267776
rect 338114 267764 338120 267776
rect 121604 267736 338120 267764
rect 121604 267724 121610 267736
rect 338114 267724 338120 267736
rect 338172 267724 338178 267776
rect 51776 267668 52316 267696
rect 51776 267656 51782 267668
rect 52362 267044 52368 267096
rect 52420 267084 52426 267096
rect 59170 267084 59176 267096
rect 52420 267056 59176 267084
rect 52420 267044 52426 267056
rect 59170 267044 59176 267056
rect 59228 267044 59234 267096
rect 54938 266976 54944 267028
rect 54996 267016 55002 267028
rect 67634 267016 67640 267028
rect 54996 266988 67640 267016
rect 54996 266976 55002 266988
rect 67634 266976 67640 266988
rect 67692 266976 67698 267028
rect 320818 266976 320824 267028
rect 320876 267016 320882 267028
rect 351178 267016 351184 267028
rect 320876 266988 351184 267016
rect 320876 266976 320882 266988
rect 351178 266976 351184 266988
rect 351236 266976 351242 267028
rect 121546 266432 121552 266484
rect 121604 266472 121610 266484
rect 312538 266472 312544 266484
rect 121604 266444 312544 266472
rect 121604 266432 121610 266444
rect 312538 266432 312544 266444
rect 312596 266432 312602 266484
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 25498 266404 25504 266416
rect 3108 266376 25504 266404
rect 3108 266364 3114 266376
rect 25498 266364 25504 266376
rect 25556 266364 25562 266416
rect 59170 266364 59176 266416
rect 59228 266404 59234 266416
rect 67634 266404 67640 266416
rect 59228 266376 67640 266404
rect 59228 266364 59234 266376
rect 67634 266364 67640 266376
rect 67692 266364 67698 266416
rect 121638 266364 121644 266416
rect 121696 266404 121702 266416
rect 349246 266404 349252 266416
rect 121696 266376 349252 266404
rect 121696 266364 121702 266376
rect 349246 266364 349252 266376
rect 349304 266364 349310 266416
rect 59262 266296 59268 266348
rect 59320 266336 59326 266348
rect 67818 266336 67824 266348
rect 59320 266308 67824 266336
rect 59320 266296 59326 266308
rect 67818 266296 67824 266308
rect 67876 266296 67882 266348
rect 123570 265616 123576 265668
rect 123628 265656 123634 265668
rect 489914 265656 489920 265668
rect 123628 265628 489920 265656
rect 123628 265616 123634 265628
rect 489914 265616 489920 265628
rect 489972 265616 489978 265668
rect 60550 264936 60556 264988
rect 60608 264976 60614 264988
rect 67726 264976 67732 264988
rect 60608 264948 67732 264976
rect 60608 264936 60614 264948
rect 67726 264936 67732 264948
rect 67784 264936 67790 264988
rect 121546 264936 121552 264988
rect 121604 264976 121610 264988
rect 300118 264976 300124 264988
rect 121604 264948 300124 264976
rect 121604 264936 121610 264948
rect 300118 264936 300124 264948
rect 300176 264936 300182 264988
rect 48222 264868 48228 264920
rect 48280 264908 48286 264920
rect 67634 264908 67640 264920
rect 48280 264880 67640 264908
rect 48280 264868 48286 264880
rect 67634 264868 67640 264880
rect 67692 264868 67698 264920
rect 36630 264188 36636 264240
rect 36688 264228 36694 264240
rect 48222 264228 48228 264240
rect 36688 264200 48228 264228
rect 36688 264188 36694 264200
rect 48222 264188 48228 264200
rect 48280 264188 48286 264240
rect 121638 264188 121644 264240
rect 121696 264228 121702 264240
rect 321554 264228 321560 264240
rect 121696 264200 321560 264228
rect 121696 264188 121702 264200
rect 321554 264188 321560 264200
rect 321612 264188 321618 264240
rect 121546 263644 121552 263696
rect 121604 263684 121610 263696
rect 270494 263684 270500 263696
rect 121604 263656 270500 263684
rect 121604 263644 121610 263656
rect 270494 263644 270500 263656
rect 270552 263644 270558 263696
rect 50706 263576 50712 263628
rect 50764 263616 50770 263628
rect 67634 263616 67640 263628
rect 50764 263588 67640 263616
rect 50764 263576 50770 263588
rect 67634 263576 67640 263588
rect 67692 263576 67698 263628
rect 137278 263576 137284 263628
rect 137336 263616 137342 263628
rect 388438 263616 388444 263628
rect 137336 263588 388444 263616
rect 137336 263576 137342 263588
rect 388438 263576 388444 263588
rect 388496 263576 388502 263628
rect 121546 263508 121552 263560
rect 121604 263548 121610 263560
rect 140774 263548 140780 263560
rect 121604 263520 140780 263548
rect 121604 263508 121610 263520
rect 140774 263508 140780 263520
rect 140832 263508 140838 263560
rect 121730 263440 121736 263492
rect 121788 263480 121794 263492
rect 128630 263480 128636 263492
rect 121788 263452 128636 263480
rect 121788 263440 121794 263452
rect 128630 263440 128636 263452
rect 128688 263480 128694 263492
rect 128906 263480 128912 263492
rect 128688 263452 128912 263480
rect 128688 263440 128694 263452
rect 128906 263440 128912 263452
rect 128964 263440 128970 263492
rect 43990 262896 43996 262948
rect 44048 262936 44054 262948
rect 52454 262936 52460 262948
rect 44048 262908 52460 262936
rect 44048 262896 44054 262908
rect 52454 262896 52460 262908
rect 52512 262896 52518 262948
rect 128906 262896 128912 262948
rect 128964 262936 128970 262948
rect 414658 262936 414664 262948
rect 128964 262908 414664 262936
rect 128964 262896 128970 262908
rect 414658 262896 414664 262908
rect 414716 262896 414722 262948
rect 53558 262828 53564 262880
rect 53616 262868 53622 262880
rect 65518 262868 65524 262880
rect 53616 262840 65524 262868
rect 53616 262828 53622 262840
rect 65518 262828 65524 262840
rect 65576 262828 65582 262880
rect 140774 262828 140780 262880
rect 140832 262868 140838 262880
rect 471238 262868 471244 262880
rect 140832 262840 471244 262868
rect 140832 262828 140838 262840
rect 471238 262828 471244 262840
rect 471296 262828 471302 262880
rect 52454 262284 52460 262336
rect 52512 262324 52518 262336
rect 53650 262324 53656 262336
rect 52512 262296 53656 262324
rect 52512 262284 52518 262296
rect 53650 262284 53656 262296
rect 53708 262324 53714 262336
rect 67726 262324 67732 262336
rect 53708 262296 67732 262324
rect 53708 262284 53714 262296
rect 67726 262284 67732 262296
rect 67784 262284 67790 262336
rect 48222 262216 48228 262268
rect 48280 262256 48286 262268
rect 67634 262256 67640 262268
rect 48280 262228 67640 262256
rect 48280 262216 48286 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 121546 262216 121552 262268
rect 121604 262256 121610 262268
rect 327074 262256 327080 262268
rect 121604 262228 327080 262256
rect 121604 262216 121610 262228
rect 327074 262216 327080 262228
rect 327132 262216 327138 262268
rect 121638 262148 121644 262200
rect 121696 262188 121702 262200
rect 137278 262188 137284 262200
rect 121696 262160 137284 262188
rect 121696 262148 121702 262160
rect 137278 262148 137284 262160
rect 137336 262148 137342 262200
rect 66162 260924 66168 260976
rect 66220 260964 66226 260976
rect 67634 260964 67640 260976
rect 66220 260936 67640 260964
rect 66220 260924 66226 260936
rect 67634 260924 67640 260936
rect 67692 260924 67698 260976
rect 57882 260856 57888 260908
rect 57940 260896 57946 260908
rect 67726 260896 67732 260908
rect 57940 260868 67732 260896
rect 57940 260856 57946 260868
rect 67726 260856 67732 260868
rect 67784 260856 67790 260908
rect 134610 260856 134616 260908
rect 134668 260896 134674 260908
rect 134886 260896 134892 260908
rect 134668 260868 134892 260896
rect 134668 260856 134674 260868
rect 134886 260856 134892 260868
rect 134944 260896 134950 260908
rect 232498 260896 232504 260908
rect 134944 260868 232504 260896
rect 134944 260856 134950 260868
rect 232498 260856 232504 260868
rect 232556 260856 232562 260908
rect 60642 260788 60648 260840
rect 60700 260828 60706 260840
rect 67634 260828 67640 260840
rect 60700 260800 67640 260828
rect 60700 260788 60706 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 121546 260788 121552 260840
rect 121604 260828 121610 260840
rect 146294 260828 146300 260840
rect 121604 260800 146300 260828
rect 121604 260788 121610 260800
rect 146294 260788 146300 260800
rect 146352 260828 146358 260840
rect 146754 260828 146760 260840
rect 146352 260800 146760 260828
rect 146352 260788 146358 260800
rect 146754 260788 146760 260800
rect 146812 260788 146818 260840
rect 121730 260176 121736 260228
rect 121788 260216 121794 260228
rect 323026 260216 323032 260228
rect 121788 260188 323032 260216
rect 121788 260176 121794 260188
rect 323026 260176 323032 260188
rect 323084 260176 323090 260228
rect 146754 260108 146760 260160
rect 146812 260148 146818 260160
rect 517606 260148 517612 260160
rect 146812 260120 517612 260148
rect 146812 260108 146818 260120
rect 517606 260108 517612 260120
rect 517664 260108 517670 260160
rect 52362 259428 52368 259480
rect 52420 259468 52426 259480
rect 67634 259468 67640 259480
rect 52420 259440 67640 259468
rect 52420 259428 52426 259440
rect 67634 259428 67640 259440
rect 67692 259428 67698 259480
rect 121546 259428 121552 259480
rect 121604 259468 121610 259480
rect 245010 259468 245016 259480
rect 121604 259440 245016 259468
rect 121604 259428 121610 259440
rect 245010 259428 245016 259440
rect 245068 259428 245074 259480
rect 121638 259360 121644 259412
rect 121696 259400 121702 259412
rect 134886 259400 134892 259412
rect 121696 259372 134892 259400
rect 121696 259360 121702 259372
rect 134886 259360 134892 259372
rect 134944 259360 134950 259412
rect 126238 258680 126244 258732
rect 126296 258720 126302 258732
rect 547874 258720 547880 258732
rect 126296 258692 547880 258720
rect 126296 258680 126302 258692
rect 547874 258680 547880 258692
rect 547932 258680 547938 258732
rect 57790 258136 57796 258188
rect 57848 258176 57854 258188
rect 67726 258176 67732 258188
rect 57848 258148 67732 258176
rect 57848 258136 57854 258148
rect 67726 258136 67732 258148
rect 67784 258136 67790 258188
rect 56318 258068 56324 258120
rect 56376 258108 56382 258120
rect 67634 258108 67640 258120
rect 56376 258080 67640 258108
rect 56376 258068 56382 258080
rect 67634 258068 67640 258080
rect 67692 258068 67698 258120
rect 121546 258068 121552 258120
rect 121604 258108 121610 258120
rect 349154 258108 349160 258120
rect 121604 258080 349160 258108
rect 121604 258068 121610 258080
rect 349154 258068 349160 258080
rect 349212 258068 349218 258120
rect 547874 258068 547880 258120
rect 547932 258108 547938 258120
rect 580166 258108 580172 258120
rect 547932 258080 580172 258108
rect 547932 258068 547938 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 36538 258000 36544 258052
rect 36596 258040 36602 258052
rect 67910 258040 67916 258052
rect 36596 258012 67916 258040
rect 36596 258000 36602 258012
rect 67910 258000 67916 258012
rect 67968 258000 67974 258052
rect 15838 257320 15844 257372
rect 15896 257360 15902 257372
rect 36538 257360 36544 257372
rect 15896 257332 36544 257360
rect 15896 257320 15902 257332
rect 36538 257320 36544 257332
rect 36596 257320 36602 257372
rect 124858 257320 124864 257372
rect 124916 257360 124922 257372
rect 485774 257360 485780 257372
rect 124916 257332 485780 257360
rect 124916 257320 124922 257332
rect 485774 257320 485780 257332
rect 485832 257320 485838 257372
rect 59262 256708 59268 256760
rect 59320 256748 59326 256760
rect 67634 256748 67640 256760
rect 59320 256720 67640 256748
rect 59320 256708 59326 256720
rect 67634 256708 67640 256720
rect 67692 256708 67698 256760
rect 121638 256708 121644 256760
rect 121696 256748 121702 256760
rect 260834 256748 260840 256760
rect 121696 256720 260840 256748
rect 121696 256708 121702 256720
rect 260834 256708 260840 256720
rect 260892 256708 260898 256760
rect 121546 256640 121552 256692
rect 121604 256680 121610 256692
rect 154574 256680 154580 256692
rect 121604 256652 154580 256680
rect 121604 256640 121610 256652
rect 154574 256640 154580 256652
rect 154632 256640 154638 256692
rect 154574 256028 154580 256080
rect 154632 256068 154638 256080
rect 399478 256068 399484 256080
rect 154632 256040 399484 256068
rect 154632 256028 154638 256040
rect 399478 256028 399484 256040
rect 399536 256028 399542 256080
rect 159358 255960 159364 256012
rect 159416 256000 159422 256012
rect 520918 256000 520924 256012
rect 159416 255972 520924 256000
rect 159416 255960 159422 255972
rect 520918 255960 520924 255972
rect 520976 255960 520982 256012
rect 65978 255348 65984 255400
rect 66036 255388 66042 255400
rect 67634 255388 67640 255400
rect 66036 255360 67640 255388
rect 66036 255348 66042 255360
rect 67634 255348 67640 255360
rect 67692 255348 67698 255400
rect 53374 255280 53380 255332
rect 53432 255320 53438 255332
rect 67726 255320 67732 255332
rect 53432 255292 67732 255320
rect 53432 255280 53438 255292
rect 67726 255280 67732 255292
rect 67784 255280 67790 255332
rect 3418 255212 3424 255264
rect 3476 255252 3482 255264
rect 33134 255252 33140 255264
rect 3476 255224 33140 255252
rect 3476 255212 3482 255224
rect 33134 255212 33140 255224
rect 33192 255212 33198 255264
rect 57606 255212 57612 255264
rect 57664 255252 57670 255264
rect 67634 255252 67640 255264
rect 57664 255224 67640 255252
rect 57664 255212 57670 255224
rect 67634 255212 67640 255224
rect 67692 255212 67698 255264
rect 33134 254532 33140 254584
rect 33192 254572 33198 254584
rect 34422 254572 34428 254584
rect 33192 254544 34428 254572
rect 33192 254532 33198 254544
rect 34422 254532 34428 254544
rect 34480 254572 34486 254584
rect 58618 254572 58624 254584
rect 34480 254544 58624 254572
rect 34480 254532 34486 254544
rect 58618 254532 58624 254544
rect 58676 254532 58682 254584
rect 187050 254532 187056 254584
rect 187108 254572 187114 254584
rect 508498 254572 508504 254584
rect 187108 254544 508504 254572
rect 187108 254532 187114 254544
rect 508498 254532 508504 254544
rect 508556 254532 508562 254584
rect 67634 253960 67640 253972
rect 60016 253932 67640 253960
rect 60016 253904 60044 253932
rect 67634 253920 67640 253932
rect 67692 253920 67698 253972
rect 121546 253920 121552 253972
rect 121604 253960 121610 253972
rect 284294 253960 284300 253972
rect 121604 253932 284300 253960
rect 121604 253920 121610 253932
rect 284294 253920 284300 253932
rect 284352 253920 284358 253972
rect 53742 253852 53748 253904
rect 53800 253892 53806 253904
rect 59998 253892 60004 253904
rect 53800 253864 60004 253892
rect 53800 253852 53806 253864
rect 59998 253852 60004 253864
rect 60056 253852 60062 253904
rect 17218 253172 17224 253224
rect 17276 253212 17282 253224
rect 35710 253212 35716 253224
rect 17276 253184 35716 253212
rect 17276 253172 17282 253184
rect 35710 253172 35716 253184
rect 35768 253212 35774 253224
rect 56226 253212 56232 253224
rect 35768 253184 56232 253212
rect 35768 253172 35774 253184
rect 56226 253172 56232 253184
rect 56284 253172 56290 253224
rect 121638 253172 121644 253224
rect 121696 253212 121702 253224
rect 400858 253212 400864 253224
rect 121696 253184 400864 253212
rect 121696 253172 121702 253184
rect 400858 253172 400864 253184
rect 400916 253172 400922 253224
rect 121546 252628 121552 252680
rect 121604 252668 121610 252680
rect 258074 252668 258080 252680
rect 121604 252640 258080 252668
rect 121604 252628 121610 252640
rect 258074 252628 258080 252640
rect 258132 252628 258138 252680
rect 56226 252560 56232 252612
rect 56284 252600 56290 252612
rect 67634 252600 67640 252612
rect 56284 252572 67640 252600
rect 56284 252560 56290 252572
rect 67634 252560 67640 252572
rect 67692 252560 67698 252612
rect 121638 252560 121644 252612
rect 121696 252600 121702 252612
rect 316770 252600 316776 252612
rect 121696 252572 316776 252600
rect 121696 252560 121702 252572
rect 316770 252560 316776 252572
rect 316828 252560 316834 252612
rect 121546 252492 121552 252544
rect 121604 252532 121610 252544
rect 143718 252532 143724 252544
rect 121604 252504 143724 252532
rect 121604 252492 121610 252504
rect 143718 252492 143724 252504
rect 143776 252532 143782 252544
rect 144822 252532 144828 252544
rect 143776 252504 144828 252532
rect 143776 252492 143782 252504
rect 144822 252492 144828 252504
rect 144880 252492 144886 252544
rect 144822 251812 144828 251864
rect 144880 251852 144886 251864
rect 472618 251852 472624 251864
rect 144880 251824 472624 251852
rect 144880 251812 144886 251824
rect 472618 251812 472624 251824
rect 472676 251812 472682 251864
rect 61838 251268 61844 251320
rect 61896 251308 61902 251320
rect 67634 251308 67640 251320
rect 61896 251280 67640 251308
rect 61896 251268 61902 251280
rect 67634 251268 67640 251280
rect 67692 251268 67698 251320
rect 53466 251200 53472 251252
rect 53524 251240 53530 251252
rect 67726 251240 67732 251252
rect 53524 251212 67732 251240
rect 53524 251200 53530 251212
rect 67726 251200 67732 251212
rect 67784 251200 67790 251252
rect 121546 251200 121552 251252
rect 121604 251240 121610 251252
rect 327258 251240 327264 251252
rect 121604 251212 327264 251240
rect 121604 251200 121610 251212
rect 327258 251200 327264 251212
rect 327316 251200 327322 251252
rect 129642 250452 129648 250504
rect 129700 250492 129706 250504
rect 478874 250492 478880 250504
rect 129700 250464 478880 250492
rect 129700 250452 129706 250464
rect 478874 250452 478880 250464
rect 478932 250452 478938 250504
rect 122098 249840 122104 249892
rect 122156 249880 122162 249892
rect 124306 249880 124312 249892
rect 122156 249852 124312 249880
rect 122156 249840 122162 249852
rect 124306 249840 124312 249852
rect 124364 249840 124370 249892
rect 60458 249772 60464 249824
rect 60516 249812 60522 249824
rect 67634 249812 67640 249824
rect 60516 249784 67640 249812
rect 60516 249772 60522 249784
rect 67634 249772 67640 249784
rect 67692 249772 67698 249824
rect 121546 249772 121552 249824
rect 121604 249812 121610 249824
rect 243538 249812 243544 249824
rect 121604 249784 243544 249812
rect 121604 249772 121610 249784
rect 243538 249772 243544 249784
rect 243596 249772 243602 249824
rect 41138 249024 41144 249076
rect 41196 249064 41202 249076
rect 57698 249064 57704 249076
rect 41196 249036 57704 249064
rect 41196 249024 41202 249036
rect 57698 249024 57704 249036
rect 57756 249024 57762 249076
rect 169018 249024 169024 249076
rect 169076 249064 169082 249076
rect 517514 249064 517520 249076
rect 169076 249036 517520 249064
rect 169076 249024 169082 249036
rect 517514 249024 517520 249036
rect 517572 249024 517578 249076
rect 57698 248480 57704 248532
rect 57756 248520 57762 248532
rect 67726 248520 67732 248532
rect 57756 248492 67732 248520
rect 57756 248480 57762 248492
rect 67726 248480 67732 248492
rect 67784 248480 67790 248532
rect 54846 248412 54852 248464
rect 54904 248452 54910 248464
rect 67634 248452 67640 248464
rect 54904 248424 67640 248452
rect 54904 248412 54910 248424
rect 67634 248412 67640 248424
rect 67692 248412 67698 248464
rect 121546 248412 121552 248464
rect 121604 248452 121610 248464
rect 345198 248452 345204 248464
rect 121604 248424 345204 248452
rect 121604 248412 121610 248424
rect 345198 248412 345204 248424
rect 345256 248412 345262 248464
rect 121454 248344 121460 248396
rect 121512 248384 121518 248396
rect 121730 248384 121736 248396
rect 121512 248356 121736 248384
rect 121512 248344 121518 248356
rect 121730 248344 121736 248356
rect 121788 248344 121794 248396
rect 63218 247120 63224 247172
rect 63276 247160 63282 247172
rect 67634 247160 67640 247172
rect 63276 247132 67640 247160
rect 63276 247120 63282 247132
rect 67634 247120 67640 247132
rect 67692 247120 67698 247172
rect 121454 247120 121460 247172
rect 121512 247160 121518 247172
rect 235258 247160 235264 247172
rect 121512 247132 235264 247160
rect 121512 247120 121518 247132
rect 235258 247120 235264 247132
rect 235316 247120 235322 247172
rect 60642 247052 60648 247104
rect 60700 247092 60706 247104
rect 67726 247092 67732 247104
rect 60700 247064 67732 247092
rect 60700 247052 60706 247064
rect 67726 247052 67732 247064
rect 67784 247052 67790 247104
rect 124030 247052 124036 247104
rect 124088 247092 124094 247104
rect 494238 247092 494244 247104
rect 124088 247064 494244 247092
rect 124088 247052 124094 247064
rect 494238 247052 494244 247064
rect 494296 247052 494302 247104
rect 124306 246372 124312 246424
rect 124364 246412 124370 246424
rect 442994 246412 443000 246424
rect 124364 246384 443000 246412
rect 124364 246372 124370 246384
rect 442994 246372 443000 246384
rect 443052 246372 443058 246424
rect 121638 246304 121644 246356
rect 121696 246344 121702 246356
rect 499666 246344 499672 246356
rect 121696 246316 499672 246344
rect 121696 246304 121702 246316
rect 499666 246304 499672 246316
rect 499724 246304 499730 246356
rect 63402 245692 63408 245744
rect 63460 245732 63466 245744
rect 67634 245732 67640 245744
rect 63460 245704 67640 245732
rect 63460 245692 63466 245704
rect 67634 245692 67640 245704
rect 67692 245692 67698 245744
rect 121546 245692 121552 245744
rect 121604 245732 121610 245744
rect 159358 245732 159364 245744
rect 121604 245704 159364 245732
rect 121604 245692 121610 245704
rect 159358 245692 159364 245704
rect 159416 245692 159422 245744
rect 61378 245664 61384 245676
rect 60752 245636 61384 245664
rect 55030 245556 55036 245608
rect 55088 245596 55094 245608
rect 60752 245596 60780 245636
rect 61378 245624 61384 245636
rect 61436 245664 61442 245676
rect 67726 245664 67732 245676
rect 61436 245636 67732 245664
rect 61436 245624 61442 245636
rect 67726 245624 67732 245636
rect 67784 245624 67790 245676
rect 121454 245624 121460 245676
rect 121512 245664 121518 245676
rect 269114 245664 269120 245676
rect 121512 245636 269120 245664
rect 121512 245624 121518 245636
rect 269114 245624 269120 245636
rect 269172 245624 269178 245676
rect 55088 245568 60780 245596
rect 55088 245556 55094 245568
rect 135898 244944 135904 244996
rect 135956 244984 135962 244996
rect 227070 244984 227076 244996
rect 135956 244956 227076 244984
rect 135956 244944 135962 244956
rect 227070 244944 227076 244956
rect 227128 244944 227134 244996
rect 122282 244876 122288 244928
rect 122340 244916 122346 244928
rect 328546 244916 328552 244928
rect 122340 244888 328552 244916
rect 122340 244876 122346 244888
rect 328546 244876 328552 244888
rect 328604 244876 328610 244928
rect 263594 244264 263600 244316
rect 263652 244304 263658 244316
rect 579614 244304 579620 244316
rect 263652 244276 579620 244304
rect 263652 244264 263658 244276
rect 579614 244264 579620 244276
rect 579672 244304 579678 244316
rect 579982 244304 579988 244316
rect 579672 244276 579988 244304
rect 579672 244264 579678 244276
rect 579982 244264 579988 244276
rect 580040 244264 580046 244316
rect 62022 244196 62028 244248
rect 62080 244236 62086 244248
rect 65886 244236 65892 244248
rect 62080 244208 65892 244236
rect 62080 244196 62086 244208
rect 65886 244196 65892 244208
rect 65944 244196 65950 244248
rect 231210 243652 231216 243704
rect 231268 243692 231274 243704
rect 318150 243692 318156 243704
rect 231268 243664 318156 243692
rect 231268 243652 231274 243664
rect 318150 243652 318156 243664
rect 318208 243652 318214 243704
rect 232590 243584 232596 243636
rect 232648 243624 232654 243636
rect 370498 243624 370504 243636
rect 232648 243596 370504 243624
rect 232648 243584 232654 243596
rect 370498 243584 370504 243596
rect 370556 243584 370562 243636
rect 121730 243516 121736 243568
rect 121788 243556 121794 243568
rect 498286 243556 498292 243568
rect 121788 243528 498292 243556
rect 121788 243516 121794 243528
rect 498286 243516 498292 243528
rect 498344 243516 498350 243568
rect 67634 243012 67640 243024
rect 55186 242984 67640 243012
rect 48038 242836 48044 242888
rect 48096 242876 48102 242888
rect 54478 242876 54484 242888
rect 48096 242848 54484 242876
rect 48096 242836 48102 242848
rect 54478 242836 54484 242848
rect 54536 242876 54542 242888
rect 55186 242876 55214 242984
rect 67634 242972 67640 242984
rect 67692 242972 67698 243024
rect 121454 242972 121460 243024
rect 121512 243012 121518 243024
rect 206370 243012 206376 243024
rect 121512 242984 206376 243012
rect 121512 242972 121518 242984
rect 206370 242972 206376 242984
rect 206428 242972 206434 243024
rect 127618 242904 127624 242956
rect 127676 242944 127682 242956
rect 231302 242944 231308 242956
rect 127676 242916 231308 242944
rect 127676 242904 127682 242916
rect 231302 242904 231308 242916
rect 231360 242904 231366 242956
rect 54536 242848 55214 242876
rect 54536 242836 54542 242848
rect 121454 242836 121460 242888
rect 121512 242876 121518 242888
rect 147674 242876 147680 242888
rect 121512 242848 147680 242876
rect 121512 242836 121518 242848
rect 147674 242836 147680 242848
rect 147732 242876 147738 242888
rect 263594 242876 263600 242888
rect 147732 242848 263600 242876
rect 147732 242836 147738 242848
rect 263594 242836 263600 242848
rect 263652 242836 263658 242888
rect 121546 242768 121552 242820
rect 121604 242808 121610 242820
rect 140774 242808 140780 242820
rect 121604 242780 140780 242808
rect 121604 242768 121610 242780
rect 140774 242768 140780 242780
rect 140832 242768 140838 242820
rect 140774 242156 140780 242208
rect 140832 242196 140838 242208
rect 413278 242196 413284 242208
rect 140832 242168 413284 242196
rect 140832 242156 140838 242168
rect 413278 242156 413284 242168
rect 413336 242156 413342 242208
rect 62022 241476 62028 241528
rect 62080 241516 62086 241528
rect 67634 241516 67640 241528
rect 62080 241488 67640 241516
rect 62080 241476 62086 241488
rect 67634 241476 67640 241488
rect 67692 241476 67698 241528
rect 121638 240728 121644 240780
rect 121696 240768 121702 240780
rect 321646 240768 321652 240780
rect 121696 240740 321652 240768
rect 121696 240728 121702 240740
rect 321646 240728 321652 240740
rect 321704 240728 321710 240780
rect 121454 240184 121460 240236
rect 121512 240224 121518 240236
rect 238110 240224 238116 240236
rect 121512 240196 238116 240224
rect 121512 240184 121518 240196
rect 238110 240184 238116 240196
rect 238168 240184 238174 240236
rect 119890 240116 119896 240168
rect 119948 240156 119954 240168
rect 331214 240156 331220 240168
rect 119948 240128 331220 240156
rect 119948 240116 119954 240128
rect 331214 240116 331220 240128
rect 331272 240116 331278 240168
rect 3142 240048 3148 240100
rect 3200 240088 3206 240100
rect 33594 240088 33600 240100
rect 3200 240060 33600 240088
rect 3200 240048 3206 240060
rect 33594 240048 33600 240060
rect 33652 240048 33658 240100
rect 75914 239776 75920 239828
rect 75972 239816 75978 239828
rect 77098 239816 77104 239828
rect 75972 239788 77104 239816
rect 75972 239776 75978 239788
rect 77098 239776 77104 239788
rect 77156 239776 77162 239828
rect 80054 239776 80060 239828
rect 80112 239816 80118 239828
rect 80962 239816 80968 239828
rect 80112 239788 80968 239816
rect 80112 239776 80118 239788
rect 80962 239776 80968 239788
rect 81020 239776 81026 239828
rect 92474 239776 92480 239828
rect 92532 239816 92538 239828
rect 93198 239816 93204 239828
rect 92532 239788 93204 239816
rect 92532 239776 92538 239788
rect 93198 239776 93204 239788
rect 93256 239776 93262 239828
rect 95234 239776 95240 239828
rect 95292 239816 95298 239828
rect 96418 239816 96424 239828
rect 95292 239788 96424 239816
rect 95292 239776 95298 239788
rect 96418 239776 96424 239788
rect 96476 239776 96482 239828
rect 96614 239776 96620 239828
rect 96672 239816 96678 239828
rect 97706 239816 97712 239828
rect 96672 239788 97712 239816
rect 96672 239776 96678 239788
rect 97706 239776 97712 239788
rect 97764 239776 97770 239828
rect 100754 239776 100760 239828
rect 100812 239816 100818 239828
rect 101570 239816 101576 239828
rect 100812 239788 101576 239816
rect 100812 239776 100818 239788
rect 101570 239776 101576 239788
rect 101628 239776 101634 239828
rect 104894 239776 104900 239828
rect 104952 239816 104958 239828
rect 106078 239816 106084 239828
rect 104952 239788 106084 239816
rect 104952 239776 104958 239788
rect 106078 239776 106084 239788
rect 106136 239776 106142 239828
rect 114554 239776 114560 239828
rect 114612 239816 114618 239828
rect 115738 239816 115744 239828
rect 114612 239788 115744 239816
rect 114612 239776 114618 239788
rect 115738 239776 115744 239788
rect 115796 239776 115802 239828
rect 117314 239776 117320 239828
rect 117372 239816 117378 239828
rect 118326 239816 118332 239828
rect 117372 239788 118332 239816
rect 117372 239776 117378 239788
rect 118326 239776 118332 239788
rect 118384 239816 118390 239828
rect 124214 239816 124220 239828
rect 118384 239788 124220 239816
rect 118384 239776 118390 239788
rect 124214 239776 124220 239788
rect 124272 239776 124278 239828
rect 63402 239504 63408 239556
rect 63460 239544 63466 239556
rect 72418 239544 72424 239556
rect 63460 239516 72424 239544
rect 63460 239504 63466 239516
rect 72418 239504 72424 239516
rect 72476 239504 72482 239556
rect 61930 239436 61936 239488
rect 61988 239476 61994 239488
rect 98638 239476 98644 239488
rect 61988 239448 98644 239476
rect 61988 239436 61994 239448
rect 98638 239436 98644 239448
rect 98696 239436 98702 239488
rect 33594 239368 33600 239420
rect 33652 239408 33658 239420
rect 34330 239408 34336 239420
rect 33652 239380 34336 239408
rect 33652 239368 33658 239380
rect 34330 239368 34336 239380
rect 34388 239408 34394 239420
rect 92658 239408 92664 239420
rect 34388 239380 92664 239408
rect 34388 239368 34394 239380
rect 92658 239368 92664 239380
rect 92716 239368 92722 239420
rect 113174 239300 113180 239352
rect 113232 239340 113238 239352
rect 114462 239340 114468 239352
rect 113232 239312 114468 239340
rect 113232 239300 113238 239312
rect 114462 239300 114468 239312
rect 114520 239300 114526 239352
rect 65886 238824 65892 238876
rect 65944 238864 65950 238876
rect 76006 238864 76012 238876
rect 65944 238836 76012 238864
rect 65944 238824 65950 238836
rect 76006 238824 76012 238836
rect 76064 238864 76070 238876
rect 76466 238864 76472 238876
rect 76064 238836 76472 238864
rect 76064 238824 76070 238836
rect 76466 238824 76472 238836
rect 76524 238824 76530 238876
rect 58618 238756 58624 238808
rect 58676 238796 58682 238808
rect 112530 238796 112536 238808
rect 58676 238768 112536 238796
rect 58676 238756 58682 238768
rect 112530 238756 112536 238768
rect 112588 238756 112594 238808
rect 121454 238756 121460 238808
rect 121512 238796 121518 238808
rect 346394 238796 346400 238808
rect 121512 238768 346400 238796
rect 121512 238756 121518 238768
rect 346394 238756 346400 238768
rect 346452 238756 346458 238808
rect 50890 238688 50896 238740
rect 50948 238728 50954 238740
rect 98362 238728 98368 238740
rect 50948 238700 98368 238728
rect 50948 238688 50954 238700
rect 98362 238688 98368 238700
rect 98420 238688 98426 238740
rect 25498 238620 25504 238672
rect 25556 238660 25562 238672
rect 56410 238660 56416 238672
rect 25556 238632 56416 238660
rect 25556 238620 25562 238632
rect 56410 238620 56416 238632
rect 56468 238660 56474 238672
rect 86770 238660 86776 238672
rect 56468 238632 86776 238660
rect 56468 238620 56474 238632
rect 86770 238620 86776 238632
rect 86828 238620 86834 238672
rect 91922 238620 91928 238672
rect 91980 238660 91986 238672
rect 123478 238660 123484 238672
rect 91980 238632 123484 238660
rect 91980 238620 91986 238632
rect 123478 238620 123484 238632
rect 123536 238620 123542 238672
rect 92658 238552 92664 238604
rect 92716 238592 92722 238604
rect 103514 238592 103520 238604
rect 92716 238564 103520 238592
rect 92716 238552 92722 238564
rect 103514 238552 103520 238564
rect 103572 238552 103578 238604
rect 105446 238212 105452 238264
rect 105504 238252 105510 238264
rect 181438 238252 181444 238264
rect 105504 238224 181444 238252
rect 105504 238212 105510 238224
rect 181438 238212 181444 238224
rect 181496 238212 181502 238264
rect 251910 238212 251916 238264
rect 251968 238252 251974 238264
rect 381538 238252 381544 238264
rect 251968 238224 381544 238252
rect 251968 238212 251974 238224
rect 381538 238212 381544 238224
rect 381596 238212 381602 238264
rect 67450 238144 67456 238196
rect 67508 238184 67514 238196
rect 259454 238184 259460 238196
rect 67508 238156 259460 238184
rect 67508 238144 67514 238156
rect 259454 238144 259460 238156
rect 259512 238144 259518 238196
rect 69934 238076 69940 238128
rect 69992 238116 69998 238128
rect 77938 238116 77944 238128
rect 69992 238088 77944 238116
rect 69992 238076 69998 238088
rect 77938 238076 77944 238088
rect 77996 238076 78002 238128
rect 102226 238076 102232 238128
rect 102284 238116 102290 238128
rect 339586 238116 339592 238128
rect 102284 238088 339592 238116
rect 102284 238076 102290 238088
rect 339586 238076 339592 238088
rect 339644 238076 339650 238128
rect 73890 238008 73896 238060
rect 73948 238048 73954 238060
rect 332594 238048 332600 238060
rect 73948 238020 332600 238048
rect 73948 238008 73954 238020
rect 332594 238008 332600 238020
rect 332652 238008 332658 238060
rect 86218 237464 86224 237516
rect 86276 237504 86282 237516
rect 86770 237504 86776 237516
rect 86276 237476 86776 237504
rect 86276 237464 86282 237476
rect 86770 237464 86776 237476
rect 86828 237464 86834 237516
rect 85482 237396 85488 237448
rect 85540 237436 85546 237448
rect 86310 237436 86316 237448
rect 85540 237408 86316 237436
rect 85540 237396 85546 237408
rect 86310 237396 86316 237408
rect 86368 237396 86374 237448
rect 89990 237396 89996 237448
rect 90048 237436 90054 237448
rect 91738 237436 91744 237448
rect 90048 237408 91744 237436
rect 90048 237396 90054 237408
rect 91738 237396 91744 237408
rect 91796 237396 91802 237448
rect 103514 237396 103520 237448
rect 103572 237436 103578 237448
rect 104158 237436 104164 237448
rect 103572 237408 104164 237436
rect 103572 237396 103578 237408
rect 104158 237396 104164 237408
rect 104216 237396 104222 237448
rect 116578 237396 116584 237448
rect 116636 237436 116642 237448
rect 117682 237436 117688 237448
rect 116636 237408 117688 237436
rect 116636 237396 116642 237408
rect 117682 237396 117688 237408
rect 117740 237396 117746 237448
rect 69198 237328 69204 237380
rect 69256 237368 69262 237380
rect 150526 237368 150532 237380
rect 69256 237340 150532 237368
rect 69256 237328 69262 237340
rect 150526 237328 150532 237340
rect 150584 237328 150590 237380
rect 52270 237260 52276 237312
rect 52328 237300 52334 237312
rect 116578 237300 116584 237312
rect 52328 237272 116584 237300
rect 52328 237260 52334 237272
rect 116578 237260 116584 237272
rect 116636 237260 116642 237312
rect 50982 237192 50988 237244
rect 51040 237232 51046 237244
rect 81618 237232 81624 237244
rect 51040 237204 81624 237232
rect 51040 237192 51046 237204
rect 81618 237192 81624 237204
rect 81676 237192 81682 237244
rect 110598 237192 110604 237244
rect 110656 237232 110662 237244
rect 132494 237232 132500 237244
rect 110656 237204 132500 237232
rect 110656 237192 110662 237204
rect 132494 237192 132500 237204
rect 132552 237192 132558 237244
rect 58986 237124 58992 237176
rect 59044 237164 59050 237176
rect 86126 237164 86132 237176
rect 59044 237136 86132 237164
rect 59044 237124 59050 237136
rect 86126 237124 86132 237136
rect 86184 237124 86190 237176
rect 150526 236648 150532 236700
rect 150584 236688 150590 236700
rect 452654 236688 452660 236700
rect 150584 236660 452660 236688
rect 150584 236648 150590 236660
rect 452654 236648 452660 236660
rect 452712 236648 452718 236700
rect 81618 235968 81624 236020
rect 81676 236008 81682 236020
rect 82078 236008 82084 236020
rect 81676 235980 82084 236008
rect 81676 235968 81682 235980
rect 82078 235968 82084 235980
rect 82136 235968 82142 236020
rect 110598 235968 110604 236020
rect 110656 236008 110662 236020
rect 111058 236008 111064 236020
rect 110656 235980 111064 236008
rect 110656 235968 110662 235980
rect 111058 235968 111064 235980
rect 111116 235968 111122 236020
rect 89622 235900 89628 235952
rect 89680 235940 89686 235952
rect 125594 235940 125600 235952
rect 89680 235912 125600 235940
rect 89680 235900 89686 235912
rect 125594 235900 125600 235912
rect 125652 235900 125658 235952
rect 63218 235356 63224 235408
rect 63276 235396 63282 235408
rect 239398 235396 239404 235408
rect 63276 235368 239404 235396
rect 63276 235356 63282 235368
rect 239398 235356 239404 235368
rect 239456 235356 239462 235408
rect 251818 235356 251824 235408
rect 251876 235396 251882 235408
rect 277394 235396 277400 235408
rect 251876 235368 277400 235396
rect 251876 235356 251882 235368
rect 277394 235356 277400 235368
rect 277452 235356 277458 235408
rect 60458 235288 60464 235340
rect 60516 235328 60522 235340
rect 278774 235328 278780 235340
rect 60516 235300 278780 235328
rect 60516 235288 60522 235300
rect 278774 235288 278780 235300
rect 278832 235288 278838 235340
rect 113266 235220 113272 235272
rect 113324 235260 113330 235272
rect 340966 235260 340972 235272
rect 113324 235232 340972 235260
rect 113324 235220 113330 235232
rect 340966 235220 340972 235232
rect 341024 235220 341030 235272
rect 46842 234540 46848 234592
rect 46900 234580 46906 234592
rect 109678 234580 109684 234592
rect 46900 234552 109684 234580
rect 46900 234540 46906 234552
rect 109678 234540 109684 234552
rect 109736 234540 109742 234592
rect 61838 234064 61844 234116
rect 61896 234104 61902 234116
rect 182818 234104 182824 234116
rect 61896 234076 182824 234104
rect 61896 234064 61902 234076
rect 182818 234064 182824 234076
rect 182876 234064 182882 234116
rect 65978 233996 65984 234048
rect 66036 234036 66042 234048
rect 251266 234036 251272 234048
rect 66036 234008 251272 234036
rect 66036 233996 66042 234008
rect 251266 233996 251272 234008
rect 251324 233996 251330 234048
rect 112530 233928 112536 233980
rect 112588 233968 112594 233980
rect 445754 233968 445760 233980
rect 112588 233940 445760 233968
rect 112588 233928 112594 233940
rect 445754 233928 445760 233940
rect 445812 233928 445818 233980
rect 86126 233860 86132 233912
rect 86184 233900 86190 233912
rect 502334 233900 502340 233912
rect 86184 233872 502340 233900
rect 86184 233860 86190 233872
rect 502334 233860 502340 233872
rect 502392 233860 502398 233912
rect 93854 233724 93860 233776
rect 93912 233764 93918 233776
rect 94038 233764 94044 233776
rect 93912 233736 94044 233764
rect 93912 233724 93918 233736
rect 94038 233724 94044 233736
rect 94096 233724 94102 233776
rect 77754 232568 77760 232620
rect 77812 232608 77818 232620
rect 352006 232608 352012 232620
rect 77812 232580 352012 232608
rect 77812 232568 77818 232580
rect 352006 232568 352012 232580
rect 352064 232568 352070 232620
rect 56226 232500 56232 232552
rect 56284 232540 56290 232552
rect 403618 232540 403624 232552
rect 56284 232512 403624 232540
rect 56284 232500 56290 232512
rect 403618 232500 403624 232512
rect 403676 232500 403682 232552
rect 515398 232500 515404 232552
rect 515456 232540 515462 232552
rect 579614 232540 579620 232552
rect 515456 232512 579620 232540
rect 515456 232500 515462 232512
rect 579614 232500 579620 232512
rect 579672 232500 579678 232552
rect 49602 231752 49608 231804
rect 49660 231792 49666 231804
rect 107286 231792 107292 231804
rect 49660 231764 107292 231792
rect 49660 231752 49666 231764
rect 107286 231752 107292 231764
rect 107344 231752 107350 231804
rect 95326 231684 95332 231736
rect 95384 231724 95390 231736
rect 126974 231724 126980 231736
rect 95384 231696 126980 231724
rect 95384 231684 95390 231696
rect 126974 231684 126980 231696
rect 127032 231724 127038 231736
rect 127434 231724 127440 231736
rect 127032 231696 127440 231724
rect 127032 231684 127038 231696
rect 127434 231684 127440 231696
rect 127492 231684 127498 231736
rect 95050 231140 95056 231192
rect 95108 231180 95114 231192
rect 347866 231180 347872 231192
rect 95108 231152 347872 231180
rect 95108 231140 95114 231152
rect 347866 231140 347872 231152
rect 347924 231140 347930 231192
rect 127434 231072 127440 231124
rect 127492 231112 127498 231124
rect 393958 231112 393964 231124
rect 127492 231084 393964 231112
rect 127492 231072 127498 231084
rect 393958 231072 393964 231084
rect 394016 231072 394022 231124
rect 84194 229916 84200 229968
rect 84252 229956 84258 229968
rect 84470 229956 84476 229968
rect 84252 229928 84476 229956
rect 84252 229916 84258 229928
rect 84470 229916 84476 229928
rect 84528 229916 84534 229968
rect 66070 229848 66076 229900
rect 66128 229888 66134 229900
rect 251358 229888 251364 229900
rect 66128 229860 251364 229888
rect 66128 229848 66134 229860
rect 251358 229848 251364 229860
rect 251416 229848 251422 229900
rect 108574 229780 108580 229832
rect 108632 229820 108638 229832
rect 331306 229820 331312 229832
rect 108632 229792 331312 229820
rect 108632 229780 108638 229792
rect 331306 229780 331312 229792
rect 331364 229780 331370 229832
rect 59998 229712 60004 229764
rect 60056 229752 60062 229764
rect 468478 229752 468484 229764
rect 60056 229724 468484 229752
rect 60056 229712 60062 229724
rect 468478 229712 468484 229724
rect 468536 229712 468542 229764
rect 83458 229032 83464 229084
rect 83516 229072 83522 229084
rect 149054 229072 149060 229084
rect 83516 229044 149060 229072
rect 83516 229032 83522 229044
rect 149054 229032 149060 229044
rect 149112 229032 149118 229084
rect 82814 228964 82820 229016
rect 82872 229004 82878 229016
rect 128354 229004 128360 229016
rect 82872 228976 128360 229004
rect 82872 228964 82878 228976
rect 128354 228964 128360 228976
rect 128412 228964 128418 229016
rect 149054 228556 149060 228608
rect 149112 228596 149118 228608
rect 171778 228596 171784 228608
rect 149112 228568 171784 228596
rect 149112 228556 149118 228568
rect 171778 228556 171784 228568
rect 171836 228556 171842 228608
rect 57882 228488 57888 228540
rect 57940 228528 57946 228540
rect 314010 228528 314016 228540
rect 57940 228500 314016 228528
rect 57940 228488 57946 228500
rect 314010 228488 314016 228500
rect 314068 228488 314074 228540
rect 53466 228420 53472 228472
rect 53524 228460 53530 228472
rect 339494 228460 339500 228472
rect 53524 228432 339500 228460
rect 53524 228420 53530 228432
rect 339494 228420 339500 228432
rect 339552 228420 339558 228472
rect 128354 228352 128360 228404
rect 128412 228392 128418 228404
rect 513374 228392 513380 228404
rect 128412 228364 513380 228392
rect 128412 228352 128418 228364
rect 513374 228352 513380 228364
rect 513432 228352 513438 228404
rect 91094 227672 91100 227724
rect 91152 227712 91158 227724
rect 131206 227712 131212 227724
rect 91152 227684 131212 227712
rect 91152 227672 91158 227684
rect 131206 227672 131212 227684
rect 131264 227712 131270 227724
rect 131758 227712 131764 227724
rect 131264 227684 131764 227712
rect 131264 227672 131270 227684
rect 131758 227672 131764 227684
rect 131816 227672 131822 227724
rect 71222 227060 71228 227112
rect 71280 227100 71286 227112
rect 255406 227100 255412 227112
rect 71280 227072 255412 227100
rect 71280 227060 71286 227072
rect 255406 227060 255412 227072
rect 255464 227060 255470 227112
rect 131206 226992 131212 227044
rect 131264 227032 131270 227044
rect 342990 227032 342996 227044
rect 131264 227004 342996 227032
rect 131264 226992 131270 227004
rect 342990 226992 342996 227004
rect 343048 226992 343054 227044
rect 64506 225632 64512 225684
rect 64564 225672 64570 225684
rect 251174 225672 251180 225684
rect 64564 225644 251180 225672
rect 64564 225632 64570 225644
rect 251174 225632 251180 225644
rect 251232 225632 251238 225684
rect 80054 225564 80060 225616
rect 80112 225604 80118 225616
rect 328638 225604 328644 225616
rect 80112 225576 328644 225604
rect 80112 225564 80118 225576
rect 328638 225564 328644 225576
rect 328696 225564 328702 225616
rect 75730 224884 75736 224936
rect 75788 224924 75794 224936
rect 142246 224924 142252 224936
rect 75788 224896 142252 224924
rect 75788 224884 75794 224896
rect 142246 224884 142252 224896
rect 142304 224924 142310 224936
rect 143442 224924 143448 224936
rect 142304 224896 143448 224924
rect 142304 224884 142310 224896
rect 143442 224884 143448 224896
rect 143500 224884 143506 224936
rect 55122 224340 55128 224392
rect 55180 224380 55186 224392
rect 151078 224380 151084 224392
rect 55180 224352 151084 224380
rect 55180 224340 55186 224352
rect 151078 224340 151084 224352
rect 151136 224340 151142 224392
rect 90082 224272 90088 224324
rect 90140 224312 90146 224324
rect 255590 224312 255596 224324
rect 90140 224284 255596 224312
rect 90140 224272 90146 224284
rect 255590 224272 255596 224284
rect 255648 224272 255654 224324
rect 143442 224204 143448 224256
rect 143500 224244 143506 224256
rect 333330 224244 333336 224256
rect 143500 224216 333336 224244
rect 143500 224204 143506 224216
rect 333330 224204 333336 224216
rect 333388 224204 333394 224256
rect 109678 223592 109684 223644
rect 109736 223632 109742 223644
rect 457438 223632 457444 223644
rect 109736 223604 457444 223632
rect 109736 223592 109742 223604
rect 457438 223592 457444 223604
rect 457496 223592 457502 223644
rect 47946 222844 47952 222896
rect 48004 222884 48010 222896
rect 276106 222884 276112 222896
rect 48004 222856 276112 222884
rect 48004 222844 48010 222856
rect 276106 222844 276112 222856
rect 276164 222844 276170 222896
rect 103606 221552 103612 221604
rect 103664 221592 103670 221604
rect 327166 221592 327172 221604
rect 103664 221564 327172 221592
rect 103664 221552 103670 221564
rect 327166 221552 327172 221564
rect 327224 221552 327230 221604
rect 61378 221484 61384 221536
rect 61436 221524 61442 221536
rect 371878 221524 371884 221536
rect 61436 221496 371884 221524
rect 61436 221484 61442 221496
rect 371878 221484 371884 221496
rect 371936 221484 371942 221536
rect 4798 221416 4804 221468
rect 4856 221456 4862 221468
rect 83458 221456 83464 221468
rect 4856 221428 83464 221456
rect 4856 221416 4862 221428
rect 83458 221416 83464 221428
rect 83516 221416 83522 221468
rect 104158 221416 104164 221468
rect 104216 221456 104222 221468
rect 466454 221456 466460 221468
rect 104216 221428 466460 221456
rect 104216 221416 104222 221428
rect 466454 221416 466460 221428
rect 466512 221416 466518 221468
rect 74626 220056 74632 220108
rect 74684 220096 74690 220108
rect 281534 220096 281540 220108
rect 74684 220068 281540 220096
rect 74684 220056 74690 220068
rect 281534 220056 281540 220068
rect 281592 220056 281598 220108
rect 57698 218764 57704 218816
rect 57756 218804 57762 218816
rect 489178 218804 489184 218816
rect 57756 218776 489184 218804
rect 57756 218764 57762 218776
rect 489178 218764 489184 218776
rect 489236 218764 489242 218816
rect 54938 218696 54944 218748
rect 54996 218736 55002 218748
rect 503714 218736 503720 218748
rect 54996 218708 503720 218736
rect 54996 218696 55002 218708
rect 503714 218696 503720 218708
rect 503772 218696 503778 218748
rect 520918 218696 520924 218748
rect 520976 218736 520982 218748
rect 580166 218736 580172 218748
rect 520976 218708 580172 218736
rect 520976 218696 520982 218708
rect 580166 218696 580172 218708
rect 580224 218696 580230 218748
rect 54846 217336 54852 217388
rect 54904 217376 54910 217388
rect 246482 217376 246488 217388
rect 54904 217348 246488 217376
rect 54904 217336 54910 217348
rect 246482 217336 246488 217348
rect 246540 217336 246546 217388
rect 59078 217268 59084 217320
rect 59136 217308 59142 217320
rect 488534 217308 488540 217320
rect 59136 217280 488540 217308
rect 59136 217268 59142 217280
rect 488534 217268 488540 217280
rect 488592 217268 488598 217320
rect 81526 216588 81532 216640
rect 81584 216628 81590 216640
rect 151814 216628 151820 216640
rect 81584 216600 151820 216628
rect 81584 216588 81590 216600
rect 151814 216588 151820 216600
rect 151872 216628 151878 216640
rect 153102 216628 153108 216640
rect 151872 216600 153108 216628
rect 151872 216588 151878 216600
rect 153102 216588 153108 216600
rect 153160 216588 153166 216640
rect 77938 215976 77944 216028
rect 77996 216016 78002 216028
rect 315390 216016 315396 216028
rect 77996 215988 315396 216016
rect 77996 215976 78002 215988
rect 315390 215976 315396 215988
rect 315448 215976 315454 216028
rect 153102 215908 153108 215960
rect 153160 215948 153166 215960
rect 473354 215948 473360 215960
rect 153160 215920 473360 215948
rect 153160 215908 153166 215920
rect 473354 215908 473360 215920
rect 473412 215908 473418 215960
rect 113174 215228 113180 215280
rect 113232 215268 113238 215280
rect 147766 215268 147772 215280
rect 113232 215240 147772 215268
rect 113232 215228 113238 215240
rect 147766 215228 147772 215240
rect 147824 215228 147830 215280
rect 78766 214684 78772 214736
rect 78824 214724 78830 214736
rect 314102 214724 314108 214736
rect 78824 214696 314108 214724
rect 78824 214684 78830 214696
rect 314102 214684 314108 214696
rect 314160 214684 314166 214736
rect 147766 214616 147772 214668
rect 147824 214656 147830 214668
rect 501046 214656 501052 214668
rect 147824 214628 501052 214656
rect 147824 214616 147830 214628
rect 501046 214616 501052 214628
rect 501104 214616 501110 214668
rect 3418 214548 3424 214600
rect 3476 214588 3482 214600
rect 36630 214588 36636 214600
rect 3476 214560 36636 214588
rect 3476 214548 3482 214560
rect 36630 214548 36636 214560
rect 36688 214588 36694 214600
rect 396718 214588 396724 214600
rect 36688 214560 396724 214588
rect 36688 214548 36694 214560
rect 396718 214548 396724 214560
rect 396776 214548 396782 214600
rect 71774 213324 71780 213376
rect 71832 213364 71838 213376
rect 329926 213364 329932 213376
rect 71832 213336 329932 213364
rect 71832 213324 71838 213336
rect 329926 213324 329932 213336
rect 329984 213324 329990 213376
rect 42702 213256 42708 213308
rect 42760 213296 42766 213308
rect 304350 213296 304356 213308
rect 42760 213268 304356 213296
rect 42760 213256 42766 213268
rect 304350 213256 304356 213268
rect 304408 213256 304414 213308
rect 93946 213188 93952 213240
rect 94004 213228 94010 213240
rect 232590 213228 232596 213240
rect 94004 213200 232596 213228
rect 94004 213188 94010 213200
rect 232590 213188 232596 213200
rect 232648 213188 232654 213240
rect 238018 213188 238024 213240
rect 238076 213228 238082 213240
rect 512086 213228 512092 213240
rect 238076 213200 512092 213228
rect 238076 213188 238082 213200
rect 512086 213188 512092 213200
rect 512144 213188 512150 213240
rect 62022 211896 62028 211948
rect 62080 211936 62086 211948
rect 267826 211936 267832 211948
rect 62080 211908 267832 211936
rect 62080 211896 62086 211908
rect 267826 211896 267832 211908
rect 267884 211896 267890 211948
rect 76006 211828 76012 211880
rect 76064 211868 76070 211880
rect 336090 211868 336096 211880
rect 76064 211840 336096 211868
rect 76064 211828 76070 211840
rect 336090 211828 336096 211840
rect 336148 211828 336154 211880
rect 52362 211760 52368 211812
rect 52420 211800 52426 211812
rect 338206 211800 338212 211812
rect 52420 211772 338212 211800
rect 52420 211760 52426 211772
rect 338206 211760 338212 211772
rect 338264 211760 338270 211812
rect 114554 210536 114560 210588
rect 114612 210576 114618 210588
rect 325878 210576 325884 210588
rect 114612 210548 325884 210576
rect 114612 210536 114618 210548
rect 325878 210536 325884 210548
rect 325936 210536 325942 210588
rect 53558 210468 53564 210520
rect 53616 210508 53622 210520
rect 273254 210508 273260 210520
rect 53616 210480 273260 210508
rect 53616 210468 53622 210480
rect 273254 210468 273260 210480
rect 273312 210468 273318 210520
rect 75914 210400 75920 210452
rect 75972 210440 75978 210452
rect 330110 210440 330116 210452
rect 75972 210412 330116 210440
rect 75972 210400 75978 210412
rect 330110 210400 330116 210412
rect 330168 210400 330174 210452
rect 100846 209176 100852 209228
rect 100904 209216 100910 209228
rect 252646 209216 252652 209228
rect 100904 209188 252652 209216
rect 100904 209176 100910 209188
rect 252646 209176 252652 209188
rect 252704 209176 252710 209228
rect 74534 209108 74540 209160
rect 74592 209148 74598 209160
rect 323118 209148 323124 209160
rect 74592 209120 323124 209148
rect 74592 209108 74598 209120
rect 323118 209108 323124 209120
rect 323176 209108 323182 209160
rect 53650 209040 53656 209092
rect 53708 209080 53714 209092
rect 480254 209080 480260 209092
rect 53708 209052 480260 209080
rect 53708 209040 53714 209052
rect 480254 209040 480260 209052
rect 480312 209040 480318 209092
rect 106274 208292 106280 208344
rect 106332 208332 106338 208344
rect 138014 208332 138020 208344
rect 106332 208304 138020 208332
rect 106332 208292 106338 208304
rect 138014 208292 138020 208304
rect 138072 208292 138078 208344
rect 87046 207748 87052 207800
rect 87104 207788 87110 207800
rect 249886 207788 249892 207800
rect 87104 207760 249892 207788
rect 87104 207748 87110 207760
rect 249886 207748 249892 207760
rect 249944 207748 249950 207800
rect 60642 207680 60648 207732
rect 60700 207720 60706 207732
rect 263594 207720 263600 207732
rect 60700 207692 263600 207720
rect 60700 207680 60706 207692
rect 263594 207680 263600 207692
rect 263652 207680 263658 207732
rect 138014 207612 138020 207664
rect 138072 207652 138078 207664
rect 354030 207652 354036 207664
rect 138072 207624 354036 207652
rect 138072 207612 138078 207624
rect 354030 207612 354036 207624
rect 354088 207612 354094 207664
rect 86310 206320 86316 206372
rect 86368 206360 86374 206372
rect 264974 206360 264980 206372
rect 86368 206332 264980 206360
rect 86368 206320 86374 206332
rect 264974 206320 264980 206332
rect 265032 206320 265038 206372
rect 86218 206252 86224 206304
rect 86276 206292 86282 206304
rect 498378 206292 498384 206304
rect 86276 206264 498384 206292
rect 86276 206252 86282 206264
rect 498378 206252 498384 206264
rect 498436 206252 498442 206304
rect 508498 206252 508504 206304
rect 508556 206292 508562 206304
rect 580166 206292 580172 206304
rect 508556 206264 580172 206292
rect 508556 206252 508562 206264
rect 580166 206252 580172 206264
rect 580224 206252 580230 206304
rect 98086 205572 98092 205624
rect 98144 205612 98150 205624
rect 143534 205612 143540 205624
rect 98144 205584 143540 205612
rect 98144 205572 98150 205584
rect 143534 205572 143540 205584
rect 143592 205612 143598 205624
rect 144822 205612 144828 205624
rect 143592 205584 144828 205612
rect 143592 205572 143598 205584
rect 144822 205572 144828 205584
rect 144880 205572 144886 205624
rect 3234 204960 3240 205012
rect 3292 205000 3298 205012
rect 120166 205000 120172 205012
rect 3292 204972 120172 205000
rect 3292 204960 3298 204972
rect 120166 204960 120172 204972
rect 120224 204960 120230 205012
rect 144822 204960 144828 205012
rect 144880 205000 144886 205012
rect 392578 205000 392584 205012
rect 144880 204972 392584 205000
rect 144880 204960 144886 204972
rect 392578 204960 392584 204972
rect 392636 204960 392642 205012
rect 50706 204892 50712 204944
rect 50764 204932 50770 204944
rect 312630 204932 312636 204944
rect 50764 204904 312636 204932
rect 50764 204892 50770 204904
rect 312630 204892 312636 204904
rect 312688 204892 312694 204944
rect 100754 203736 100760 203788
rect 100812 203776 100818 203788
rect 254210 203776 254216 203788
rect 100812 203748 254216 203776
rect 100812 203736 100818 203748
rect 254210 203736 254216 203748
rect 254268 203736 254274 203788
rect 91738 203668 91744 203720
rect 91796 203708 91802 203720
rect 263686 203708 263692 203720
rect 91796 203680 263692 203708
rect 91796 203668 91802 203680
rect 263686 203668 263692 203680
rect 263744 203668 263750 203720
rect 90358 203600 90364 203652
rect 90416 203640 90422 203652
rect 349338 203640 349344 203652
rect 90416 203612 349344 203640
rect 90416 203600 90422 203612
rect 349338 203600 349344 203612
rect 349396 203600 349402 203652
rect 195330 203532 195336 203584
rect 195388 203572 195394 203584
rect 501230 203572 501236 203584
rect 195388 203544 501236 203572
rect 195388 203532 195394 203544
rect 501230 203532 501236 203544
rect 501288 203532 501294 203584
rect 99466 202240 99472 202292
rect 99524 202280 99530 202292
rect 255498 202280 255504 202292
rect 99524 202252 255504 202280
rect 99524 202240 99530 202252
rect 255498 202240 255504 202252
rect 255556 202240 255562 202292
rect 98638 202172 98644 202224
rect 98696 202212 98702 202224
rect 269206 202212 269212 202224
rect 98696 202184 269212 202212
rect 98696 202172 98702 202184
rect 269206 202172 269212 202184
rect 269264 202172 269270 202224
rect 7558 202104 7564 202156
rect 7616 202144 7622 202156
rect 125686 202144 125692 202156
rect 7616 202116 125692 202144
rect 7616 202104 7622 202116
rect 125686 202104 125692 202116
rect 125744 202144 125750 202156
rect 465074 202144 465080 202156
rect 125744 202116 465080 202144
rect 125744 202104 125750 202116
rect 465074 202104 465080 202116
rect 465132 202104 465138 202156
rect 50798 200880 50804 200932
rect 50856 200920 50862 200932
rect 259638 200920 259644 200932
rect 50856 200892 259644 200920
rect 50856 200880 50862 200892
rect 259638 200880 259644 200892
rect 259696 200880 259702 200932
rect 117314 200812 117320 200864
rect 117372 200852 117378 200864
rect 337470 200852 337476 200864
rect 117372 200824 337476 200852
rect 117372 200812 117378 200824
rect 337470 200812 337476 200824
rect 337528 200812 337534 200864
rect 70394 200744 70400 200796
rect 70452 200784 70458 200796
rect 334158 200784 334164 200796
rect 70452 200756 334164 200784
rect 70452 200744 70458 200756
rect 334158 200744 334164 200756
rect 334216 200744 334222 200796
rect 133138 199656 133144 199708
rect 133196 199696 133202 199708
rect 262306 199696 262312 199708
rect 133196 199668 262312 199696
rect 133196 199656 133202 199668
rect 262306 199656 262312 199668
rect 262364 199656 262370 199708
rect 115934 199588 115940 199640
rect 115992 199628 115998 199640
rect 249978 199628 249984 199640
rect 115992 199600 249984 199628
rect 115992 199588 115998 199600
rect 249978 199588 249984 199600
rect 250036 199588 250042 199640
rect 77294 199520 77300 199572
rect 77352 199560 77358 199572
rect 266446 199560 266452 199572
rect 77352 199532 266452 199560
rect 77352 199520 77358 199532
rect 266446 199520 266452 199532
rect 266504 199520 266510 199572
rect 45370 199452 45376 199504
rect 45428 199492 45434 199504
rect 318242 199492 318248 199504
rect 45428 199464 318248 199492
rect 45428 199452 45434 199464
rect 318242 199452 318248 199464
rect 318300 199452 318306 199504
rect 403618 199452 403624 199504
rect 403676 199492 403682 199504
rect 459554 199492 459560 199504
rect 403676 199464 459560 199492
rect 403676 199452 403682 199464
rect 459554 199452 459560 199464
rect 459612 199452 459618 199504
rect 233878 199384 233884 199436
rect 233936 199424 233942 199436
rect 509234 199424 509240 199436
rect 233936 199396 509240 199424
rect 233936 199384 233942 199396
rect 509234 199384 509240 199396
rect 509292 199384 509298 199436
rect 92566 198092 92572 198144
rect 92624 198132 92630 198144
rect 259546 198132 259552 198144
rect 92624 198104 259552 198132
rect 92624 198092 92630 198104
rect 259546 198092 259552 198104
rect 259604 198092 259610 198144
rect 52178 198024 52184 198076
rect 52236 198064 52242 198076
rect 238018 198064 238024 198076
rect 52236 198036 238024 198064
rect 52236 198024 52242 198036
rect 238018 198024 238024 198036
rect 238076 198024 238082 198076
rect 231302 197956 231308 198008
rect 231360 197996 231366 198008
rect 510614 197996 510620 198008
rect 231360 197968 510620 197996
rect 231360 197956 231366 197968
rect 510614 197956 510620 197968
rect 510672 197956 510678 198008
rect 111794 196800 111800 196852
rect 111852 196840 111858 196852
rect 254026 196840 254032 196852
rect 111852 196812 254032 196840
rect 111852 196800 111858 196812
rect 254026 196800 254032 196812
rect 254084 196800 254090 196852
rect 57790 196732 57796 196784
rect 57848 196772 57854 196784
rect 271874 196772 271880 196784
rect 57848 196744 271880 196772
rect 57848 196732 57854 196744
rect 271874 196732 271880 196744
rect 271932 196732 271938 196784
rect 92474 196664 92480 196716
rect 92532 196704 92538 196716
rect 328730 196704 328736 196716
rect 92532 196676 328736 196704
rect 92532 196664 92538 196676
rect 328730 196664 328736 196676
rect 328788 196664 328794 196716
rect 69014 196596 69020 196648
rect 69072 196636 69078 196648
rect 496906 196636 496912 196648
rect 69072 196608 496912 196636
rect 69072 196596 69078 196608
rect 496906 196596 496912 196608
rect 496964 196596 496970 196648
rect 56318 195440 56324 195492
rect 56376 195480 56382 195492
rect 260926 195480 260932 195492
rect 56376 195452 260932 195480
rect 56376 195440 56382 195452
rect 260926 195440 260932 195452
rect 260984 195440 260990 195492
rect 103698 195372 103704 195424
rect 103756 195412 103762 195424
rect 321738 195412 321744 195424
rect 103756 195384 321744 195412
rect 103756 195372 103762 195384
rect 321738 195372 321744 195384
rect 321796 195372 321802 195424
rect 49510 195304 49516 195356
rect 49568 195344 49574 195356
rect 273346 195344 273352 195356
rect 49568 195316 273352 195344
rect 49568 195304 49574 195316
rect 273346 195304 273352 195316
rect 273404 195304 273410 195356
rect 89622 195236 89628 195288
rect 89680 195276 89686 195288
rect 506566 195276 506572 195288
rect 89680 195248 506572 195276
rect 89680 195236 89686 195248
rect 506566 195236 506572 195248
rect 506624 195236 506630 195288
rect 102134 193876 102140 193928
rect 102192 193916 102198 193928
rect 252830 193916 252836 193928
rect 102192 193888 252836 193916
rect 102192 193876 102198 193888
rect 252830 193876 252836 193888
rect 252888 193876 252894 193928
rect 93854 193808 93860 193860
rect 93912 193848 93918 193860
rect 352098 193848 352104 193860
rect 93912 193820 352104 193848
rect 93912 193808 93918 193820
rect 352098 193808 352104 193820
rect 352156 193808 352162 193860
rect 3418 193196 3424 193248
rect 3476 193236 3482 193248
rect 4062 193236 4068 193248
rect 3476 193208 4068 193236
rect 3476 193196 3482 193208
rect 4062 193196 4068 193208
rect 4120 193236 4126 193248
rect 509326 193236 509332 193248
rect 4120 193208 509332 193236
rect 4120 193196 4126 193208
rect 509326 193196 509332 193208
rect 509384 193196 509390 193248
rect 221458 192720 221464 192772
rect 221516 192760 221522 192772
rect 280154 192760 280160 192772
rect 221516 192732 280160 192760
rect 221516 192720 221522 192732
rect 280154 192720 280160 192732
rect 280212 192720 280218 192772
rect 43898 192652 43904 192704
rect 43956 192692 43962 192704
rect 199378 192692 199384 192704
rect 43956 192664 199384 192692
rect 43956 192652 43962 192664
rect 199378 192652 199384 192664
rect 199436 192652 199442 192704
rect 214650 192652 214656 192704
rect 214708 192692 214714 192704
rect 277486 192692 277492 192704
rect 214708 192664 277492 192692
rect 214708 192652 214714 192664
rect 277486 192652 277492 192664
rect 277544 192652 277550 192704
rect 196710 192584 196716 192636
rect 196768 192624 196774 192636
rect 471974 192624 471980 192636
rect 196768 192596 471980 192624
rect 196768 192584 196774 192596
rect 471974 192584 471980 192596
rect 472032 192584 472038 192636
rect 53374 192516 53380 192568
rect 53432 192556 53438 192568
rect 346486 192556 346492 192568
rect 53432 192528 346492 192556
rect 53432 192516 53438 192528
rect 346486 192516 346492 192528
rect 346544 192516 346550 192568
rect 54478 192448 54484 192500
rect 54536 192488 54542 192500
rect 469214 192488 469220 192500
rect 54536 192460 469220 192488
rect 54536 192448 54542 192460
rect 469214 192448 469220 192460
rect 469272 192448 469278 192500
rect 224310 191292 224316 191344
rect 224368 191332 224374 191344
rect 276198 191332 276204 191344
rect 224368 191304 276204 191332
rect 224368 191292 224374 191304
rect 276198 191292 276204 191304
rect 276256 191292 276262 191344
rect 48130 191224 48136 191276
rect 48188 191264 48194 191276
rect 267918 191264 267924 191276
rect 48188 191236 267924 191264
rect 48188 191224 48194 191236
rect 267918 191224 267924 191236
rect 267976 191224 267982 191276
rect 46750 191156 46756 191208
rect 46808 191196 46814 191208
rect 343634 191196 343640 191208
rect 46808 191168 343640 191196
rect 46808 191156 46814 191168
rect 343634 191156 343640 191168
rect 343692 191156 343698 191208
rect 419626 191156 419632 191208
rect 419684 191196 419690 191208
rect 580166 191196 580172 191208
rect 419684 191168 580172 191196
rect 419684 191156 419690 191168
rect 580166 191156 580172 191168
rect 580224 191156 580230 191208
rect 119338 191088 119344 191140
rect 119396 191128 119402 191140
rect 494330 191128 494336 191140
rect 119396 191100 494336 191128
rect 119396 191088 119402 191100
rect 494330 191088 494336 191100
rect 494388 191088 494394 191140
rect 100662 190544 100668 190596
rect 100720 190584 100726 190596
rect 170490 190584 170496 190596
rect 100720 190556 170496 190584
rect 100720 190544 100726 190556
rect 170490 190544 170496 190556
rect 170548 190544 170554 190596
rect 106182 190476 106188 190528
rect 106240 190516 106246 190528
rect 195330 190516 195336 190528
rect 106240 190488 195336 190516
rect 106240 190476 106246 190488
rect 195330 190476 195336 190488
rect 195388 190476 195394 190528
rect 249058 190000 249064 190052
rect 249116 190040 249122 190052
rect 271966 190040 271972 190052
rect 249116 190012 271972 190040
rect 249116 190000 249122 190012
rect 271966 190000 271972 190012
rect 272024 190000 272030 190052
rect 155218 189932 155224 189984
rect 155276 189972 155282 189984
rect 265158 189972 265164 189984
rect 155276 189944 265164 189972
rect 155276 189932 155282 189944
rect 265158 189932 265164 189944
rect 265216 189932 265222 189984
rect 78674 189864 78680 189916
rect 78732 189904 78738 189916
rect 258166 189904 258172 189916
rect 78732 189876 258172 189904
rect 78732 189864 78738 189876
rect 258166 189864 258172 189876
rect 258224 189864 258230 189916
rect 59262 189796 59268 189848
rect 59320 189836 59326 189848
rect 350626 189836 350632 189848
rect 59320 189808 350632 189836
rect 59320 189796 59326 189808
rect 350626 189796 350632 189808
rect 350684 189796 350690 189848
rect 116578 189728 116584 189780
rect 116636 189768 116642 189780
rect 505278 189768 505284 189780
rect 116636 189740 505284 189768
rect 116636 189728 116642 189740
rect 505278 189728 505284 189740
rect 505336 189728 505342 189780
rect 102042 189048 102048 189100
rect 102100 189088 102106 189100
rect 173158 189088 173164 189100
rect 102100 189060 173164 189088
rect 102100 189048 102106 189060
rect 173158 189048 173164 189060
rect 173216 189048 173222 189100
rect 3510 188844 3516 188896
rect 3568 188884 3574 188896
rect 7558 188884 7564 188896
rect 3568 188856 7564 188884
rect 3568 188844 3574 188856
rect 7558 188844 7564 188856
rect 7616 188844 7622 188896
rect 213270 188504 213276 188556
rect 213328 188544 213334 188556
rect 274634 188544 274640 188556
rect 213328 188516 274640 188544
rect 213328 188504 213334 188516
rect 274634 188504 274640 188516
rect 274692 188504 274698 188556
rect 130378 188436 130384 188488
rect 130436 188476 130442 188488
rect 249334 188476 249340 188488
rect 130436 188448 249340 188476
rect 130436 188436 130442 188448
rect 249334 188436 249340 188448
rect 249392 188436 249398 188488
rect 99374 188368 99380 188420
rect 99432 188408 99438 188420
rect 327350 188408 327356 188420
rect 99432 188380 327356 188408
rect 99432 188368 99438 188380
rect 327350 188368 327356 188380
rect 327408 188368 327414 188420
rect 63310 188300 63316 188352
rect 63368 188340 63374 188352
rect 324314 188340 324320 188352
rect 63368 188312 324320 188340
rect 63368 188300 63374 188312
rect 324314 188300 324320 188312
rect 324372 188300 324378 188352
rect 135898 187688 135904 187740
rect 135956 187728 135962 187740
rect 214650 187728 214656 187740
rect 135956 187700 214656 187728
rect 135956 187688 135962 187700
rect 214650 187688 214656 187700
rect 214708 187688 214714 187740
rect 229738 187280 229744 187332
rect 229796 187320 229802 187332
rect 256694 187320 256700 187332
rect 229796 187292 256700 187320
rect 229796 187280 229802 187292
rect 256694 187280 256700 187292
rect 256752 187280 256758 187332
rect 222930 187212 222936 187264
rect 222988 187252 222994 187264
rect 274726 187252 274732 187264
rect 222988 187224 274732 187252
rect 222988 187212 222994 187224
rect 274726 187212 274732 187224
rect 274784 187212 274790 187264
rect 88334 187144 88340 187196
rect 88392 187184 88398 187196
rect 325970 187184 325976 187196
rect 88392 187156 325976 187184
rect 88392 187144 88398 187156
rect 325970 187144 325976 187156
rect 326028 187144 326034 187196
rect 73154 187076 73160 187128
rect 73212 187116 73218 187128
rect 321830 187116 321836 187128
rect 73212 187088 321836 187116
rect 73212 187076 73218 187088
rect 321830 187076 321836 187088
rect 321888 187076 321894 187128
rect 104894 187008 104900 187060
rect 104952 187048 104958 187060
rect 354674 187048 354680 187060
rect 104952 187020 354680 187048
rect 104952 187008 104958 187020
rect 354674 187008 354680 187020
rect 354732 187008 354738 187060
rect 72418 186940 72424 186992
rect 72476 186980 72482 186992
rect 345290 186980 345296 186992
rect 72476 186952 345296 186980
rect 72476 186940 72482 186952
rect 345290 186940 345296 186952
rect 345348 186940 345354 186992
rect 419258 186940 419264 186992
rect 419316 186980 419322 186992
rect 580258 186980 580264 186992
rect 419316 186952 580264 186980
rect 419316 186940 419322 186952
rect 580258 186940 580264 186952
rect 580316 186940 580322 186992
rect 133138 186328 133144 186380
rect 133196 186368 133202 186380
rect 209222 186368 209228 186380
rect 133196 186340 209228 186368
rect 133196 186328 133202 186340
rect 209222 186328 209228 186340
rect 209280 186328 209286 186380
rect 227070 185784 227076 185836
rect 227128 185824 227134 185836
rect 270678 185824 270684 185836
rect 227128 185796 270684 185824
rect 227128 185784 227134 185796
rect 270678 185784 270684 185796
rect 270736 185784 270742 185836
rect 151078 185716 151084 185768
rect 151136 185756 151142 185768
rect 336734 185756 336740 185768
rect 151136 185728 336740 185756
rect 151136 185716 151142 185728
rect 336734 185716 336740 185728
rect 336792 185716 336798 185768
rect 48222 185648 48228 185700
rect 48280 185688 48286 185700
rect 247678 185688 247684 185700
rect 48280 185660 247684 185688
rect 48280 185648 48286 185660
rect 247678 185648 247684 185660
rect 247736 185648 247742 185700
rect 67542 185580 67548 185632
rect 67600 185620 67606 185632
rect 318334 185620 318340 185632
rect 67600 185592 318340 185620
rect 67600 185580 67606 185592
rect 318334 185580 318340 185592
rect 318392 185580 318398 185632
rect 422938 185580 422944 185632
rect 422996 185620 423002 185632
rect 450538 185620 450544 185632
rect 422996 185592 450544 185620
rect 422996 185580 423002 185592
rect 450538 185580 450544 185592
rect 450596 185580 450602 185632
rect 124122 184968 124128 185020
rect 124180 185008 124186 185020
rect 167822 185008 167828 185020
rect 124180 184980 167828 185008
rect 124180 184968 124186 184980
rect 167822 184968 167828 184980
rect 167880 184968 167886 185020
rect 126882 184900 126888 184952
rect 126940 184940 126946 184952
rect 214742 184940 214748 184952
rect 126940 184912 214748 184940
rect 126940 184900 126946 184912
rect 214742 184900 214748 184912
rect 214800 184900 214806 184952
rect 429930 184832 429936 184884
rect 429988 184872 429994 184884
rect 430574 184872 430580 184884
rect 429988 184844 430580 184872
rect 429988 184832 429994 184844
rect 430574 184832 430580 184844
rect 430632 184832 430638 184884
rect 152458 184424 152464 184476
rect 152516 184464 152522 184476
rect 187050 184464 187056 184476
rect 152516 184436 187056 184464
rect 152516 184424 152522 184436
rect 187050 184424 187056 184436
rect 187108 184424 187114 184476
rect 225598 184424 225604 184476
rect 225656 184464 225662 184476
rect 269298 184464 269304 184476
rect 225656 184436 269304 184464
rect 225656 184424 225662 184436
rect 269298 184424 269304 184436
rect 269356 184424 269362 184476
rect 86954 184356 86960 184408
rect 87012 184396 87018 184408
rect 196802 184396 196808 184408
rect 87012 184368 196808 184396
rect 87012 184356 87018 184368
rect 196802 184356 196808 184368
rect 196860 184356 196866 184408
rect 206370 184356 206376 184408
rect 206428 184396 206434 184408
rect 335446 184396 335452 184408
rect 206428 184368 335452 184396
rect 206428 184356 206434 184368
rect 335446 184356 335452 184368
rect 335504 184356 335510 184408
rect 96706 184288 96712 184340
rect 96764 184328 96770 184340
rect 263778 184328 263784 184340
rect 96764 184300 263784 184328
rect 96764 184288 96770 184300
rect 263778 184288 263784 184300
rect 263836 184288 263842 184340
rect 467098 184288 467104 184340
rect 467156 184328 467162 184340
rect 499758 184328 499764 184340
rect 467156 184300 499764 184328
rect 467156 184288 467162 184300
rect 499758 184288 499764 184300
rect 499816 184288 499822 184340
rect 95234 184220 95240 184272
rect 95292 184260 95298 184272
rect 321278 184260 321284 184272
rect 95292 184232 321284 184260
rect 95292 184220 95298 184232
rect 321278 184220 321284 184232
rect 321336 184220 321342 184272
rect 472618 184220 472624 184272
rect 472676 184260 472682 184272
rect 506658 184260 506664 184272
rect 472676 184232 506664 184260
rect 472676 184220 472682 184232
rect 506658 184220 506664 184232
rect 506716 184220 506722 184272
rect 107654 184152 107660 184204
rect 107712 184192 107718 184204
rect 338298 184192 338304 184204
rect 107712 184164 338304 184192
rect 107712 184152 107718 184164
rect 338298 184152 338304 184164
rect 338356 184152 338362 184204
rect 464338 184152 464344 184204
rect 464396 184192 464402 184204
rect 512178 184192 512184 184204
rect 464396 184164 512184 184192
rect 464396 184152 464402 184164
rect 512178 184152 512184 184164
rect 512236 184152 512242 184204
rect 345014 184016 345020 184068
rect 345072 184056 345078 184068
rect 345658 184056 345664 184068
rect 345072 184028 345664 184056
rect 345072 184016 345078 184028
rect 345658 184016 345664 184028
rect 345716 184016 345722 184068
rect 121362 183540 121368 183592
rect 121420 183580 121426 183592
rect 166350 183580 166356 183592
rect 121420 183552 166356 183580
rect 121420 183540 121426 183552
rect 166350 183540 166356 183552
rect 166408 183540 166414 183592
rect 345658 183540 345664 183592
rect 345716 183580 345722 183592
rect 499850 183580 499856 183592
rect 345716 183552 499856 183580
rect 345716 183540 345722 183552
rect 499850 183540 499856 183552
rect 499908 183540 499914 183592
rect 240778 183132 240784 183184
rect 240836 183172 240842 183184
rect 261110 183172 261116 183184
rect 240836 183144 261116 183172
rect 240836 183132 240842 183144
rect 261110 183132 261116 183144
rect 261168 183132 261174 183184
rect 220170 183064 220176 183116
rect 220228 183104 220234 183116
rect 268010 183104 268016 183116
rect 220228 183076 268016 183104
rect 220228 183064 220234 183076
rect 268010 183064 268016 183076
rect 268068 183064 268074 183116
rect 142798 182996 142804 183048
rect 142856 183036 142862 183048
rect 245378 183036 245384 183048
rect 142856 183008 245384 183036
rect 142856 182996 142862 183008
rect 245378 182996 245384 183008
rect 245436 182996 245442 183048
rect 110414 182928 110420 182980
rect 110472 182968 110478 182980
rect 252738 182968 252744 182980
rect 110472 182940 252744 182968
rect 110472 182928 110478 182940
rect 252738 182928 252744 182940
rect 252796 182928 252802 182980
rect 45462 182860 45468 182912
rect 45520 182900 45526 182912
rect 265066 182900 265072 182912
rect 45520 182872 265072 182900
rect 45520 182860 45526 182872
rect 265066 182860 265072 182872
rect 265124 182860 265130 182912
rect 316678 182860 316684 182912
rect 316736 182900 316742 182912
rect 339678 182900 339684 182912
rect 316736 182872 339684 182900
rect 316736 182860 316742 182872
rect 339678 182860 339684 182872
rect 339736 182860 339742 182912
rect 96614 182792 96620 182844
rect 96672 182832 96678 182844
rect 206370 182832 206376 182844
rect 96672 182804 206376 182832
rect 96672 182792 96678 182804
rect 206370 182792 206376 182804
rect 206428 182792 206434 182844
rect 232498 182792 232504 182844
rect 232556 182832 232562 182844
rect 502518 182832 502524 182844
rect 232556 182804 502524 182832
rect 232556 182792 232562 182804
rect 502518 182792 502524 182804
rect 502576 182792 502582 182844
rect 130746 182248 130752 182300
rect 130804 182288 130810 182300
rect 166534 182288 166540 182300
rect 130804 182260 166540 182288
rect 130804 182248 130810 182260
rect 166534 182248 166540 182260
rect 166592 182248 166598 182300
rect 110690 182180 110696 182232
rect 110748 182220 110754 182232
rect 169018 182220 169024 182232
rect 110748 182192 169024 182220
rect 110748 182180 110754 182192
rect 169018 182180 169024 182192
rect 169076 182180 169082 182232
rect 457438 182112 457444 182164
rect 457496 182152 457502 182164
rect 458174 182152 458180 182164
rect 457496 182124 458180 182152
rect 457496 182112 457502 182124
rect 458174 182112 458180 182124
rect 458232 182112 458238 182164
rect 475378 182112 475384 182164
rect 475436 182152 475442 182164
rect 476574 182152 476580 182164
rect 475436 182124 476580 182152
rect 475436 182112 475442 182124
rect 476574 182112 476580 182124
rect 476632 182112 476638 182164
rect 160738 181704 160744 181756
rect 160796 181744 160802 181756
rect 203518 181744 203524 181756
rect 160796 181716 203524 181744
rect 160796 181704 160802 181716
rect 203518 181704 203524 181716
rect 203576 181704 203582 181756
rect 233970 181704 233976 181756
rect 234028 181744 234034 181756
rect 256878 181744 256884 181756
rect 234028 181716 256884 181744
rect 234028 181704 234034 181716
rect 256878 181704 256884 181716
rect 256936 181704 256942 181756
rect 489178 181704 489184 181756
rect 489236 181744 489242 181756
rect 492858 181744 492864 181756
rect 489236 181716 492864 181744
rect 489236 181704 489242 181716
rect 492858 181704 492864 181716
rect 492916 181704 492922 181756
rect 202230 181636 202236 181688
rect 202288 181676 202294 181688
rect 334066 181676 334072 181688
rect 202288 181648 334072 181676
rect 202288 181636 202294 181648
rect 334066 181636 334072 181648
rect 334124 181636 334130 181688
rect 483658 181636 483664 181688
rect 483716 181676 483722 181688
rect 502426 181676 502432 181688
rect 483716 181648 502432 181676
rect 483716 181636 483722 181648
rect 502426 181636 502432 181648
rect 502484 181636 502490 181688
rect 171778 181568 171784 181620
rect 171836 181608 171842 181620
rect 439406 181608 439412 181620
rect 171836 181580 439412 181608
rect 171836 181568 171842 181580
rect 439406 181568 439412 181580
rect 439464 181568 439470 181620
rect 482278 181568 482284 181620
rect 482336 181608 482342 181620
rect 502610 181608 502616 181620
rect 482336 181580 502616 181608
rect 482336 181568 482342 181580
rect 502610 181568 502616 181580
rect 502668 181568 502674 181620
rect 56502 181500 56508 181552
rect 56560 181540 56566 181552
rect 343726 181540 343732 181552
rect 56560 181512 343732 181540
rect 56560 181500 56566 181512
rect 343726 181500 343732 181512
rect 343784 181500 343790 181552
rect 471238 181500 471244 181552
rect 471296 181540 471302 181552
rect 508038 181540 508044 181552
rect 471296 181512 508044 181540
rect 471296 181500 471302 181512
rect 508038 181500 508044 181512
rect 508096 181500 508102 181552
rect 166258 181432 166264 181484
rect 166316 181472 166322 181484
rect 483566 181472 483572 181484
rect 166316 181444 483572 181472
rect 166316 181432 166322 181444
rect 483566 181432 483572 181444
rect 483624 181432 483630 181484
rect 485038 181432 485044 181484
rect 485096 181472 485102 181484
rect 505186 181472 505192 181484
rect 485096 181444 505192 181472
rect 485096 181432 485102 181444
rect 505186 181432 505192 181444
rect 505244 181432 505250 181484
rect 447778 181296 447784 181348
rect 447836 181336 447842 181348
rect 451366 181336 451372 181348
rect 447836 181308 451372 181336
rect 447836 181296 447842 181308
rect 451366 181296 451372 181308
rect 451424 181296 451430 181348
rect 132402 181024 132408 181076
rect 132460 181064 132466 181076
rect 164970 181064 164976 181076
rect 132460 181036 164976 181064
rect 132460 181024 132466 181036
rect 164970 181024 164976 181036
rect 165028 181024 165034 181076
rect 118510 180956 118516 181008
rect 118568 180996 118574 181008
rect 171870 180996 171876 181008
rect 118568 180968 171876 180996
rect 118568 180956 118574 180968
rect 171870 180956 171876 180968
rect 171928 180956 171934 181008
rect 114370 180888 114376 180940
rect 114428 180928 114434 180940
rect 167730 180928 167736 180940
rect 114428 180900 167736 180928
rect 114428 180888 114434 180900
rect 167730 180888 167736 180900
rect 167788 180888 167794 180940
rect 97074 180820 97080 180872
rect 97132 180860 97138 180872
rect 170582 180860 170588 180872
rect 97132 180832 170588 180860
rect 97132 180820 97138 180832
rect 170582 180820 170588 180832
rect 170640 180820 170646 180872
rect 385678 180820 385684 180872
rect 385736 180860 385742 180872
rect 491294 180860 491300 180872
rect 385736 180832 491300 180860
rect 385736 180820 385742 180832
rect 491294 180820 491300 180832
rect 491352 180820 491358 180872
rect 246390 180412 246396 180464
rect 246448 180452 246454 180464
rect 249058 180452 249064 180464
rect 246448 180424 249064 180452
rect 246448 180412 246454 180424
rect 249058 180412 249064 180424
rect 249116 180412 249122 180464
rect 314010 180412 314016 180464
rect 314068 180452 314074 180464
rect 331490 180452 331496 180464
rect 314068 180424 331496 180452
rect 314068 180412 314074 180424
rect 331490 180412 331496 180424
rect 331548 180412 331554 180464
rect 236638 180344 236644 180396
rect 236696 180384 236702 180396
rect 249426 180384 249432 180396
rect 236696 180356 249432 180384
rect 236696 180344 236702 180356
rect 249426 180344 249432 180356
rect 249484 180344 249490 180396
rect 316770 180344 316776 180396
rect 316828 180384 316834 180396
rect 341150 180384 341156 180396
rect 316828 180356 341156 180384
rect 316828 180344 316834 180356
rect 341150 180344 341156 180356
rect 341208 180344 341214 180396
rect 232590 180276 232596 180328
rect 232648 180316 232654 180328
rect 256786 180316 256792 180328
rect 232648 180288 256792 180316
rect 232648 180276 232654 180288
rect 256786 180276 256792 180288
rect 256844 180276 256850 180328
rect 305730 180276 305736 180328
rect 305788 180316 305794 180328
rect 333238 180316 333244 180328
rect 305788 180288 333244 180316
rect 305788 180276 305794 180288
rect 333238 180276 333244 180288
rect 333296 180276 333302 180328
rect 159358 180208 159364 180260
rect 159416 180248 159422 180260
rect 259730 180248 259736 180260
rect 159416 180220 259736 180248
rect 159416 180208 159422 180220
rect 259730 180208 259736 180220
rect 259788 180208 259794 180260
rect 311158 180208 311164 180260
rect 311216 180248 311222 180260
rect 343818 180248 343824 180260
rect 311216 180220 343824 180248
rect 311216 180208 311222 180220
rect 343818 180208 343824 180220
rect 343876 180208 343882 180260
rect 493318 180208 493324 180260
rect 493376 180248 493382 180260
rect 507946 180248 507952 180260
rect 493376 180220 507952 180248
rect 493376 180208 493382 180220
rect 507946 180208 507952 180220
rect 508004 180208 508010 180260
rect 29638 180140 29644 180192
rect 29696 180180 29702 180192
rect 109678 180180 109684 180192
rect 29696 180152 109684 180180
rect 29696 180140 29702 180152
rect 109678 180140 109684 180152
rect 109736 180140 109742 180192
rect 226978 180140 226984 180192
rect 227036 180180 227042 180192
rect 389818 180180 389824 180192
rect 227036 180152 389824 180180
rect 227036 180140 227042 180152
rect 389818 180140 389824 180152
rect 389876 180140 389882 180192
rect 468478 180140 468484 180192
rect 468536 180180 468542 180192
rect 503898 180180 503904 180192
rect 468536 180152 503904 180180
rect 468536 180140 468542 180152
rect 503898 180140 503904 180152
rect 503956 180140 503962 180192
rect 82078 180072 82084 180124
rect 82136 180112 82142 180124
rect 495618 180112 495624 180124
rect 82136 180084 495624 180112
rect 82136 180072 82142 180084
rect 495618 180072 495624 180084
rect 495676 180072 495682 180124
rect 407758 180004 407764 180056
rect 407816 180044 407822 180056
rect 408402 180044 408408 180056
rect 407816 180016 408408 180044
rect 407816 180004 407822 180016
rect 408402 180004 408408 180016
rect 408460 180004 408466 180056
rect 114002 179528 114008 179580
rect 114060 179568 114066 179580
rect 166258 179568 166264 179580
rect 114060 179540 166264 179568
rect 114060 179528 114066 179540
rect 166258 179528 166264 179540
rect 166316 179528 166322 179580
rect 115842 179460 115848 179512
rect 115900 179500 115906 179512
rect 167914 179500 167920 179512
rect 115900 179472 167920 179500
rect 115900 179460 115906 179472
rect 167914 179460 167920 179472
rect 167972 179460 167978 179512
rect 108114 179392 108120 179444
rect 108172 179432 108178 179444
rect 169202 179432 169208 179444
rect 108172 179404 169208 179432
rect 108172 179392 108178 179404
rect 169202 179392 169208 179404
rect 169260 179392 169266 179444
rect 408402 179392 408408 179444
rect 408460 179432 408466 179444
rect 574738 179432 574744 179444
rect 408460 179404 574744 179432
rect 408460 179392 408466 179404
rect 574738 179392 574744 179404
rect 574796 179392 574802 179444
rect 235258 178984 235264 179036
rect 235316 179024 235322 179036
rect 250070 179024 250076 179036
rect 235316 178996 250076 179024
rect 235316 178984 235322 178996
rect 250070 178984 250076 178996
rect 250128 178984 250134 179036
rect 238110 178916 238116 178968
rect 238168 178956 238174 178968
rect 258350 178956 258356 178968
rect 238168 178928 258356 178956
rect 238168 178916 238174 178928
rect 258350 178916 258356 178928
rect 258408 178916 258414 178968
rect 84194 178848 84200 178900
rect 84252 178888 84258 178900
rect 323210 178888 323216 178900
rect 84252 178860 323216 178888
rect 84252 178848 84258 178860
rect 323210 178848 323216 178860
rect 323268 178848 323274 178900
rect 69106 178780 69112 178832
rect 69164 178820 69170 178832
rect 324406 178820 324412 178832
rect 69164 178792 324412 178820
rect 69164 178780 69170 178792
rect 324406 178780 324412 178792
rect 324464 178780 324470 178832
rect 66162 178712 66168 178764
rect 66220 178752 66226 178764
rect 324498 178752 324504 178764
rect 66220 178724 324504 178752
rect 66220 178712 66226 178724
rect 324498 178712 324504 178724
rect 324556 178712 324562 178764
rect 331858 178712 331864 178764
rect 331916 178752 331922 178764
rect 342438 178752 342444 178764
rect 331916 178724 342444 178752
rect 331916 178712 331922 178724
rect 342438 178712 342444 178724
rect 342496 178712 342502 178764
rect 100754 178644 100760 178696
rect 100812 178684 100818 178696
rect 133874 178684 133880 178696
rect 100812 178656 133880 178684
rect 100812 178644 100818 178656
rect 133874 178644 133880 178656
rect 133932 178684 133938 178696
rect 505094 178684 505100 178696
rect 133932 178656 505100 178684
rect 133932 178644 133938 178656
rect 505094 178644 505100 178656
rect 505152 178644 505158 178696
rect 122098 178032 122104 178084
rect 122156 178072 122162 178084
rect 166442 178072 166448 178084
rect 122156 178044 166448 178072
rect 122156 178032 122162 178044
rect 166442 178032 166448 178044
rect 166500 178032 166506 178084
rect 360930 178032 360936 178084
rect 360988 178072 360994 178084
rect 416774 178072 416780 178084
rect 360988 178044 416780 178072
rect 360988 178032 360994 178044
rect 416774 178032 416780 178044
rect 416832 178032 416838 178084
rect 119522 177964 119528 178016
rect 119580 178004 119586 178016
rect 135898 178004 135904 178016
rect 119580 177976 135904 178004
rect 119580 177964 119586 177976
rect 135898 177964 135904 177976
rect 135956 177964 135962 178016
rect 243538 177964 243544 178016
rect 243596 178004 243602 178016
rect 249150 178004 249156 178016
rect 243596 177976 249156 178004
rect 243596 177964 243602 177976
rect 249150 177964 249156 177976
rect 249208 177964 249214 178016
rect 109954 177896 109960 177948
rect 110012 177936 110018 177948
rect 121454 177936 121460 177948
rect 110012 177908 121460 177936
rect 110012 177896 110018 177908
rect 121454 177896 121460 177908
rect 121512 177896 121518 177948
rect 127894 177896 127900 177948
rect 127952 177936 127958 177948
rect 133138 177936 133144 177948
rect 127952 177908 133144 177936
rect 127952 177896 127958 177908
rect 133138 177896 133144 177908
rect 133196 177896 133202 177948
rect 245378 177896 245384 177948
rect 245436 177936 245442 177948
rect 249242 177936 249248 177948
rect 245436 177908 249248 177936
rect 245436 177896 245442 177908
rect 249242 177896 249248 177908
rect 249300 177896 249306 177948
rect 318334 177556 318340 177608
rect 318392 177596 318398 177608
rect 329834 177596 329840 177608
rect 318392 177568 329840 177596
rect 318392 177556 318398 177568
rect 329834 177556 329840 177568
rect 329892 177556 329898 177608
rect 246298 177488 246304 177540
rect 246356 177528 246362 177540
rect 261018 177528 261024 177540
rect 246356 177500 261024 177528
rect 246356 177488 246362 177500
rect 261018 177488 261024 177500
rect 261076 177488 261082 177540
rect 314102 177488 314108 177540
rect 314160 177528 314166 177540
rect 332686 177528 332692 177540
rect 314160 177500 332692 177528
rect 314160 177488 314166 177500
rect 332686 177488 332692 177500
rect 332744 177488 332750 177540
rect 240870 177420 240876 177472
rect 240928 177460 240934 177472
rect 262490 177460 262496 177472
rect 240928 177432 262496 177460
rect 240928 177420 240934 177432
rect 262490 177420 262496 177432
rect 262548 177420 262554 177472
rect 318150 177420 318156 177472
rect 318208 177460 318214 177472
rect 336826 177460 336832 177472
rect 318208 177432 336832 177460
rect 318208 177420 318214 177432
rect 336826 177420 336832 177432
rect 336884 177420 336890 177472
rect 231118 177352 231124 177404
rect 231176 177392 231182 177404
rect 258258 177392 258264 177404
rect 231176 177364 258264 177392
rect 231176 177352 231182 177364
rect 258258 177352 258264 177364
rect 258316 177352 258322 177404
rect 313918 177352 313924 177404
rect 313976 177392 313982 177404
rect 341058 177392 341064 177404
rect 313976 177364 341064 177392
rect 313976 177352 313982 177364
rect 341058 177352 341064 177364
rect 341116 177352 341122 177404
rect 7558 177284 7564 177336
rect 7616 177324 7622 177336
rect 100754 177324 100760 177336
rect 7616 177296 100760 177324
rect 7616 177284 7622 177296
rect 100754 177284 100760 177296
rect 100812 177284 100818 177336
rect 214558 177284 214564 177336
rect 214616 177324 214622 177336
rect 270586 177324 270592 177336
rect 214616 177296 270592 177324
rect 214616 177284 214622 177296
rect 270586 177284 270592 177296
rect 270644 177284 270650 177336
rect 289078 177284 289084 177336
rect 289136 177324 289142 177336
rect 338758 177324 338764 177336
rect 289136 177296 338764 177324
rect 289136 177284 289142 177296
rect 338758 177284 338764 177296
rect 338816 177284 338822 177336
rect 134426 177012 134432 177064
rect 134484 177052 134490 177064
rect 165522 177052 165528 177064
rect 134484 177024 165528 177052
rect 134484 177012 134490 177024
rect 165522 177012 165528 177024
rect 165580 177012 165586 177064
rect 124490 176944 124496 176996
rect 124548 176984 124554 176996
rect 170674 176984 170680 176996
rect 124548 176956 170680 176984
rect 124548 176944 124554 176956
rect 170674 176944 170680 176956
rect 170732 176944 170738 176996
rect 496998 176944 497004 176996
rect 497056 176984 497062 176996
rect 498470 176984 498476 176996
rect 497056 176956 498476 176984
rect 497056 176944 497062 176956
rect 498470 176944 498476 176956
rect 498528 176944 498534 176996
rect 107010 176876 107016 176928
rect 107068 176916 107074 176928
rect 165246 176916 165252 176928
rect 107068 176888 165252 176916
rect 107068 176876 107074 176888
rect 165246 176876 165252 176888
rect 165304 176876 165310 176928
rect 103330 176808 103336 176860
rect 103388 176848 103394 176860
rect 169110 176848 169116 176860
rect 103388 176820 169116 176848
rect 103388 176808 103394 176820
rect 169110 176808 169116 176820
rect 169168 176808 169174 176860
rect 136082 176740 136088 176792
rect 136140 176780 136146 176792
rect 213914 176780 213920 176792
rect 136140 176752 213920 176780
rect 136140 176740 136146 176752
rect 213914 176740 213920 176752
rect 213972 176740 213978 176792
rect 133138 176672 133144 176724
rect 133196 176712 133202 176724
rect 133196 176684 213500 176712
rect 133196 176672 133202 176684
rect 213472 176644 213500 176684
rect 356698 176672 356704 176724
rect 356756 176712 356762 176724
rect 416774 176712 416780 176724
rect 356756 176684 416780 176712
rect 356756 176672 356762 176684
rect 416774 176672 416780 176684
rect 416832 176672 416838 176724
rect 496998 176672 497004 176724
rect 497056 176712 497062 176724
rect 500954 176712 500960 176724
rect 497056 176684 500960 176712
rect 497056 176672 497062 176684
rect 500954 176672 500960 176684
rect 501012 176672 501018 176724
rect 214006 176644 214012 176656
rect 213472 176616 214012 176644
rect 214006 176604 214012 176616
rect 214064 176604 214070 176656
rect 128170 176264 128176 176316
rect 128228 176304 128234 176316
rect 166994 176304 167000 176316
rect 128228 176276 167000 176304
rect 128228 176264 128234 176276
rect 166994 176264 167000 176276
rect 167052 176264 167058 176316
rect 158898 176196 158904 176248
rect 158956 176236 158962 176248
rect 211890 176236 211896 176248
rect 158956 176208 211896 176236
rect 158956 176196 158962 176208
rect 211890 176196 211896 176208
rect 211948 176196 211954 176248
rect 148226 176128 148232 176180
rect 148284 176168 148290 176180
rect 209130 176168 209136 176180
rect 148284 176140 209136 176168
rect 148284 176128 148290 176140
rect 209130 176128 209136 176140
rect 209188 176128 209194 176180
rect 104618 176060 104624 176112
rect 104676 176100 104682 176112
rect 169294 176100 169300 176112
rect 104676 176072 169300 176100
rect 104676 176060 104682 176072
rect 169294 176060 169300 176072
rect 169352 176060 169358 176112
rect 244918 176060 244924 176112
rect 244976 176100 244982 176112
rect 254118 176100 254124 176112
rect 244976 176072 254124 176100
rect 244976 176060 244982 176072
rect 254118 176060 254124 176072
rect 254176 176060 254182 176112
rect 315390 176060 315396 176112
rect 315448 176100 315454 176112
rect 330018 176100 330024 176112
rect 315448 176072 330024 176100
rect 315448 176060 315454 176072
rect 330018 176060 330024 176072
rect 330076 176060 330082 176112
rect 129458 175992 129464 176044
rect 129516 176032 129522 176044
rect 214098 176032 214104 176044
rect 129516 176004 214104 176032
rect 129516 175992 129522 176004
rect 214098 175992 214104 176004
rect 214156 175992 214162 176044
rect 245010 175992 245016 176044
rect 245068 176032 245074 176044
rect 262398 176032 262404 176044
rect 245068 176004 262404 176032
rect 245068 175992 245074 176004
rect 262398 175992 262404 176004
rect 262456 175992 262462 176044
rect 315298 175992 315304 176044
rect 315356 176032 315362 176044
rect 334250 176032 334256 176044
rect 315356 176004 334256 176032
rect 315356 175992 315362 176004
rect 334250 175992 334256 176004
rect 334308 175992 334314 176044
rect 14458 175924 14464 175976
rect 14516 175964 14522 175976
rect 111058 175964 111064 175976
rect 14516 175936 111064 175964
rect 14516 175924 14522 175936
rect 111058 175924 111064 175936
rect 111116 175924 111122 175976
rect 116946 175924 116952 175976
rect 117004 175964 117010 175976
rect 213362 175964 213368 175976
rect 117004 175936 213368 175964
rect 117004 175924 117010 175936
rect 213362 175924 213368 175936
rect 213420 175924 213426 175976
rect 239398 175924 239404 175976
rect 239456 175964 239462 175976
rect 262214 175964 262220 175976
rect 239456 175936 262220 175964
rect 239456 175924 239462 175936
rect 262214 175924 262220 175936
rect 262272 175924 262278 175976
rect 312538 175924 312544 175976
rect 312596 175964 312602 175976
rect 331398 175964 331404 175976
rect 312596 175936 331404 175964
rect 312596 175924 312602 175936
rect 331398 175924 331404 175936
rect 331456 175924 331462 175976
rect 319438 175584 319444 175636
rect 319496 175624 319502 175636
rect 321462 175624 321468 175636
rect 319496 175596 321468 175624
rect 319496 175584 319502 175596
rect 321462 175584 321468 175596
rect 321520 175584 321526 175636
rect 165522 175176 165528 175228
rect 165580 175216 165586 175228
rect 213914 175216 213920 175228
rect 165580 175188 213920 175216
rect 165580 175176 165586 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 165246 174496 165252 174548
rect 165304 174536 165310 174548
rect 214558 174536 214564 174548
rect 165304 174508 214564 174536
rect 165304 174496 165310 174508
rect 214558 174496 214564 174508
rect 214616 174496 214622 174548
rect 496998 174224 497004 174276
rect 497056 174264 497062 174276
rect 501138 174264 501144 174276
rect 497056 174236 501144 174264
rect 497056 174224 497062 174236
rect 501138 174224 501144 174236
rect 501196 174224 501202 174276
rect 266998 174088 267004 174140
rect 267056 174128 267062 174140
rect 307662 174128 307668 174140
rect 267056 174100 307668 174128
rect 267056 174088 267062 174100
rect 307662 174088 307668 174100
rect 307720 174088 307726 174140
rect 302878 174020 302884 174072
rect 302936 174060 302942 174072
rect 307570 174060 307576 174072
rect 302936 174032 307576 174060
rect 302936 174020 302942 174032
rect 307570 174020 307576 174032
rect 307628 174020 307634 174072
rect 297450 173952 297456 174004
rect 297508 173992 297514 174004
rect 307478 173992 307484 174004
rect 297508 173964 307484 173992
rect 297508 173952 297514 173964
rect 307478 173952 307484 173964
rect 307536 173952 307542 174004
rect 355318 173884 355324 173936
rect 355376 173924 355382 173936
rect 416774 173924 416780 173936
rect 355376 173896 416780 173924
rect 355376 173884 355382 173896
rect 416774 173884 416780 173896
rect 416832 173884 416838 173936
rect 164970 173816 164976 173868
rect 165028 173856 165034 173868
rect 213914 173856 213920 173868
rect 165028 173828 213920 173856
rect 165028 173816 165034 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 324314 173816 324320 173868
rect 324372 173856 324378 173868
rect 333974 173856 333980 173868
rect 324372 173828 333980 173856
rect 324372 173816 324378 173828
rect 333974 173816 333980 173828
rect 334032 173816 334038 173868
rect 166534 173748 166540 173800
rect 166592 173788 166598 173800
rect 214006 173788 214012 173800
rect 166592 173760 214012 173788
rect 166592 173748 166598 173760
rect 214006 173748 214012 173760
rect 214064 173748 214070 173800
rect 285030 172660 285036 172712
rect 285088 172700 285094 172712
rect 307570 172700 307576 172712
rect 285088 172672 307576 172700
rect 285088 172660 285094 172672
rect 307570 172660 307576 172672
rect 307628 172660 307634 172712
rect 271138 172592 271144 172644
rect 271196 172632 271202 172644
rect 307478 172632 307484 172644
rect 271196 172604 307484 172632
rect 271196 172592 271202 172604
rect 307478 172592 307484 172604
rect 307536 172592 307542 172644
rect 264238 172524 264244 172576
rect 264296 172564 264302 172576
rect 307662 172564 307668 172576
rect 264296 172536 307668 172564
rect 264296 172524 264302 172536
rect 307662 172524 307668 172536
rect 307720 172524 307726 172576
rect 166994 172456 167000 172508
rect 167052 172496 167058 172508
rect 213914 172496 213920 172508
rect 167052 172468 213920 172496
rect 167052 172456 167058 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 252462 172456 252468 172508
rect 252520 172496 252526 172508
rect 267734 172496 267740 172508
rect 252520 172468 267740 172496
rect 252520 172456 252526 172468
rect 267734 172456 267740 172468
rect 267792 172456 267798 172508
rect 252370 172388 252376 172440
rect 252428 172428 252434 172440
rect 256878 172428 256884 172440
rect 252428 172400 256884 172428
rect 252428 172388 252434 172400
rect 256878 172388 256884 172400
rect 256936 172388 256942 172440
rect 304442 171232 304448 171284
rect 304500 171272 304506 171284
rect 307662 171272 307668 171284
rect 304500 171244 307668 171272
rect 304500 171232 304506 171244
rect 307662 171232 307668 171244
rect 307720 171232 307726 171284
rect 286410 171164 286416 171216
rect 286468 171204 286474 171216
rect 306558 171204 306564 171216
rect 286468 171176 306564 171204
rect 286468 171164 286474 171176
rect 306558 171164 306564 171176
rect 306616 171164 306622 171216
rect 273990 171096 273996 171148
rect 274048 171136 274054 171148
rect 307294 171136 307300 171148
rect 274048 171108 307300 171136
rect 274048 171096 274054 171108
rect 307294 171096 307300 171108
rect 307352 171096 307358 171148
rect 353938 171096 353944 171148
rect 353996 171136 354002 171148
rect 416774 171136 416780 171148
rect 353996 171108 416780 171136
rect 353996 171096 354002 171108
rect 416774 171096 416780 171108
rect 416832 171096 416838 171148
rect 209222 171028 209228 171080
rect 209280 171068 209286 171080
rect 213914 171068 213920 171080
rect 209280 171040 213920 171068
rect 209280 171028 209286 171040
rect 213914 171028 213920 171040
rect 213972 171028 213978 171080
rect 252370 171028 252376 171080
rect 252428 171068 252434 171080
rect 262214 171068 262220 171080
rect 252428 171040 262220 171068
rect 252428 171028 252434 171040
rect 262214 171028 262220 171040
rect 262272 171028 262278 171080
rect 324314 171028 324320 171080
rect 324372 171068 324378 171080
rect 334250 171068 334256 171080
rect 324372 171040 334256 171068
rect 324372 171028 324378 171040
rect 334250 171028 334256 171040
rect 334308 171028 334314 171080
rect 252462 170960 252468 171012
rect 252520 171000 252526 171012
rect 261110 171000 261116 171012
rect 252520 170972 261116 171000
rect 252520 170960 252526 170972
rect 261110 170960 261116 170972
rect 261168 170960 261174 171012
rect 496998 170756 497004 170808
rect 497056 170796 497062 170808
rect 499850 170796 499856 170808
rect 497056 170768 499856 170796
rect 497056 170756 497062 170768
rect 499850 170756 499856 170768
rect 499908 170756 499914 170808
rect 252462 170076 252468 170128
rect 252520 170116 252526 170128
rect 259638 170116 259644 170128
rect 252520 170088 259644 170116
rect 252520 170076 252526 170088
rect 259638 170076 259644 170088
rect 259696 170076 259702 170128
rect 307018 170076 307024 170128
rect 307076 170116 307082 170128
rect 308582 170116 308588 170128
rect 307076 170088 308588 170116
rect 307076 170076 307082 170088
rect 308582 170076 308588 170088
rect 308640 170076 308646 170128
rect 289262 169872 289268 169924
rect 289320 169912 289326 169924
rect 307294 169912 307300 169924
rect 289320 169884 307300 169912
rect 289320 169872 289326 169884
rect 307294 169872 307300 169884
rect 307352 169872 307358 169924
rect 268562 169804 268568 169856
rect 268620 169844 268626 169856
rect 307570 169844 307576 169856
rect 268620 169816 307576 169844
rect 268620 169804 268626 169816
rect 307570 169804 307576 169816
rect 307628 169804 307634 169856
rect 262858 169736 262864 169788
rect 262916 169776 262922 169788
rect 307662 169776 307668 169788
rect 262916 169748 307668 169776
rect 262916 169736 262922 169748
rect 307662 169736 307668 169748
rect 307720 169736 307726 169788
rect 334618 169736 334624 169788
rect 334676 169776 334682 169788
rect 416774 169776 416780 169788
rect 334676 169748 416780 169776
rect 334676 169736 334682 169748
rect 416774 169736 416780 169748
rect 416832 169736 416838 169788
rect 167822 169668 167828 169720
rect 167880 169708 167886 169720
rect 214006 169708 214012 169720
rect 167880 169680 214012 169708
rect 167880 169668 167886 169680
rect 214006 169668 214012 169680
rect 214064 169668 214070 169720
rect 170674 169600 170680 169652
rect 170732 169640 170738 169652
rect 213914 169640 213920 169652
rect 170732 169612 213920 169640
rect 170732 169600 170738 169612
rect 213914 169600 213920 169612
rect 213972 169600 213978 169652
rect 252462 169600 252468 169652
rect 252520 169640 252526 169652
rect 263778 169640 263784 169652
rect 252520 169612 263784 169640
rect 252520 169600 252526 169612
rect 263778 169600 263784 169612
rect 263836 169600 263842 169652
rect 252370 169532 252376 169584
rect 252428 169572 252434 169584
rect 265158 169572 265164 169584
rect 252428 169544 265164 169572
rect 252428 169532 252434 169544
rect 265158 169532 265164 169544
rect 265216 169532 265222 169584
rect 290550 168988 290556 169040
rect 290608 169028 290614 169040
rect 307110 169028 307116 169040
rect 290608 169000 307116 169028
rect 290608 168988 290614 169000
rect 307110 168988 307116 169000
rect 307168 168988 307174 169040
rect 278222 168444 278228 168496
rect 278280 168484 278286 168496
rect 307662 168484 307668 168496
rect 278280 168456 307668 168484
rect 278280 168444 278286 168456
rect 307662 168444 307668 168456
rect 307720 168444 307726 168496
rect 267090 168376 267096 168428
rect 267148 168416 267154 168428
rect 307478 168416 307484 168428
rect 267148 168388 307484 168416
rect 267148 168376 267154 168388
rect 307478 168376 307484 168388
rect 307536 168376 307542 168428
rect 166442 168308 166448 168360
rect 166500 168348 166506 168360
rect 213914 168348 213920 168360
rect 166500 168320 213920 168348
rect 166500 168308 166506 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 252370 168308 252376 168360
rect 252428 168348 252434 168360
rect 262306 168348 262312 168360
rect 252428 168320 262312 168348
rect 252428 168308 252434 168320
rect 262306 168308 262312 168320
rect 262364 168308 262370 168360
rect 324314 168308 324320 168360
rect 324372 168348 324378 168360
rect 329834 168348 329840 168360
rect 324372 168320 329840 168348
rect 324372 168308 324378 168320
rect 329834 168308 329840 168320
rect 329892 168308 329898 168360
rect 496998 168308 497004 168360
rect 497056 168348 497062 168360
rect 502334 168348 502340 168360
rect 497056 168320 502340 168348
rect 497056 168308 497062 168320
rect 502334 168308 502340 168320
rect 502392 168348 502398 168360
rect 503622 168348 503628 168360
rect 502392 168320 503628 168348
rect 502392 168308 502398 168320
rect 503622 168308 503628 168320
rect 503680 168308 503686 168360
rect 166350 168240 166356 168292
rect 166408 168280 166414 168292
rect 214006 168280 214012 168292
rect 166408 168252 214012 168280
rect 166408 168240 166414 168252
rect 214006 168240 214012 168252
rect 214064 168240 214070 168292
rect 252462 167900 252468 167952
rect 252520 167940 252526 167952
rect 258074 167940 258080 167952
rect 252520 167912 258080 167940
rect 252520 167900 252526 167912
rect 258074 167900 258080 167912
rect 258132 167900 258138 167952
rect 265802 167628 265808 167680
rect 265860 167668 265866 167680
rect 307570 167668 307576 167680
rect 265860 167640 307576 167668
rect 265860 167628 265866 167640
rect 307570 167628 307576 167640
rect 307628 167628 307634 167680
rect 503622 167628 503628 167680
rect 503680 167668 503686 167680
rect 542998 167668 543004 167680
rect 503680 167640 543004 167668
rect 503680 167628 503686 167640
rect 542998 167628 543004 167640
rect 543056 167628 543062 167680
rect 287882 167084 287888 167136
rect 287940 167124 287946 167136
rect 307662 167124 307668 167136
rect 287940 167096 307668 167124
rect 287940 167084 287946 167096
rect 307662 167084 307668 167096
rect 307720 167084 307726 167136
rect 257338 167016 257344 167068
rect 257396 167056 257402 167068
rect 307478 167056 307484 167068
rect 257396 167028 307484 167056
rect 257396 167016 257402 167028
rect 307478 167016 307484 167028
rect 307536 167016 307542 167068
rect 171870 166948 171876 167000
rect 171928 166988 171934 167000
rect 213914 166988 213920 167000
rect 171928 166960 213920 166988
rect 171928 166948 171934 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 324314 166948 324320 167000
rect 324372 166988 324378 167000
rect 335538 166988 335544 167000
rect 324372 166960 335544 166988
rect 324372 166948 324378 166960
rect 335538 166948 335544 166960
rect 335596 166948 335602 167000
rect 496998 166948 497004 167000
rect 497056 166988 497062 167000
rect 505278 166988 505284 167000
rect 497056 166960 505284 166988
rect 497056 166948 497062 166960
rect 505278 166948 505284 166960
rect 505336 166948 505342 167000
rect 252462 166336 252468 166388
rect 252520 166376 252526 166388
rect 258350 166376 258356 166388
rect 252520 166348 258356 166376
rect 252520 166336 252526 166348
rect 258350 166336 258356 166348
rect 258408 166336 258414 166388
rect 269758 166268 269764 166320
rect 269816 166308 269822 166320
rect 307570 166308 307576 166320
rect 269816 166280 307576 166308
rect 269816 166268 269822 166280
rect 307570 166268 307576 166280
rect 307628 166268 307634 166320
rect 505278 166268 505284 166320
rect 505336 166308 505342 166320
rect 544378 166308 544384 166320
rect 505336 166280 544384 166308
rect 505336 166268 505342 166280
rect 544378 166268 544384 166280
rect 544436 166268 544442 166320
rect 252462 166064 252468 166116
rect 252520 166104 252526 166116
rect 259546 166104 259552 166116
rect 252520 166076 259552 166104
rect 252520 166064 252526 166076
rect 259546 166064 259552 166076
rect 259604 166064 259610 166116
rect 258718 165588 258724 165640
rect 258776 165628 258782 165640
rect 306742 165628 306748 165640
rect 258776 165600 306748 165628
rect 258776 165588 258782 165600
rect 306742 165588 306748 165600
rect 306800 165588 306806 165640
rect 546494 165588 546500 165640
rect 546552 165628 546558 165640
rect 580166 165628 580172 165640
rect 546552 165600 580172 165628
rect 546552 165588 546558 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 167914 165520 167920 165572
rect 167972 165560 167978 165572
rect 213914 165560 213920 165572
rect 167972 165532 213920 165560
rect 167972 165520 167978 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 252278 165520 252284 165572
rect 252336 165560 252342 165572
rect 276106 165560 276112 165572
rect 252336 165532 276112 165560
rect 252336 165520 252342 165532
rect 276106 165520 276112 165532
rect 276164 165520 276170 165572
rect 324406 165520 324412 165572
rect 324464 165560 324470 165572
rect 339586 165560 339592 165572
rect 324464 165532 339592 165560
rect 324464 165520 324470 165532
rect 339586 165520 339592 165532
rect 339644 165520 339650 165572
rect 497090 165520 497096 165572
rect 497148 165560 497154 165572
rect 507854 165560 507860 165572
rect 497148 165532 507860 165560
rect 497148 165520 497154 165532
rect 507854 165520 507860 165532
rect 507912 165520 507918 165572
rect 167730 165452 167736 165504
rect 167788 165492 167794 165504
rect 214006 165492 214012 165504
rect 167788 165464 214012 165492
rect 167788 165452 167794 165464
rect 214006 165452 214012 165464
rect 214064 165452 214070 165504
rect 252462 165452 252468 165504
rect 252520 165492 252526 165504
rect 266354 165492 266360 165504
rect 252520 165464 266360 165492
rect 252520 165452 252526 165464
rect 266354 165452 266360 165464
rect 266412 165452 266418 165504
rect 324314 165452 324320 165504
rect 324372 165492 324378 165504
rect 330018 165492 330024 165504
rect 324372 165464 330024 165492
rect 324372 165452 324378 165464
rect 330018 165452 330024 165464
rect 330076 165452 330082 165504
rect 252370 165384 252376 165436
rect 252428 165424 252434 165436
rect 263686 165424 263692 165436
rect 252428 165396 263692 165424
rect 252428 165384 252434 165396
rect 263686 165384 263692 165396
rect 263744 165384 263750 165436
rect 264422 164840 264428 164892
rect 264480 164880 264486 164892
rect 307662 164880 307668 164892
rect 264480 164852 307668 164880
rect 264480 164840 264486 164852
rect 307662 164840 307668 164852
rect 307720 164840 307726 164892
rect 496998 164840 497004 164892
rect 497056 164880 497062 164892
rect 503898 164880 503904 164892
rect 497056 164852 503904 164880
rect 497056 164840 497062 164852
rect 503898 164840 503904 164852
rect 503956 164840 503962 164892
rect 507854 164840 507860 164892
rect 507912 164880 507918 164892
rect 536098 164880 536104 164892
rect 507912 164852 536104 164880
rect 507912 164840 507918 164852
rect 536098 164840 536104 164852
rect 536156 164840 536162 164892
rect 503898 164432 503904 164484
rect 503956 164472 503962 164484
rect 504450 164472 504456 164484
rect 503956 164444 504456 164472
rect 503956 164432 503962 164444
rect 504450 164432 504456 164444
rect 504508 164432 504514 164484
rect 294690 164296 294696 164348
rect 294748 164336 294754 164348
rect 307570 164336 307576 164348
rect 294748 164308 307576 164336
rect 294748 164296 294754 164308
rect 307570 164296 307576 164308
rect 307628 164296 307634 164348
rect 260282 164228 260288 164280
rect 260340 164268 260346 164280
rect 307662 164268 307668 164280
rect 260340 164240 307668 164268
rect 260340 164228 260346 164240
rect 307662 164228 307668 164240
rect 307720 164228 307726 164280
rect 340230 164228 340236 164280
rect 340288 164268 340294 164280
rect 416774 164268 416780 164280
rect 340288 164240 416780 164268
rect 340288 164228 340294 164240
rect 416774 164228 416780 164240
rect 416832 164228 416838 164280
rect 166258 164160 166264 164212
rect 166316 164200 166322 164212
rect 213914 164200 213920 164212
rect 166316 164172 213920 164200
rect 166316 164160 166322 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 252370 164160 252376 164212
rect 252428 164200 252434 164212
rect 273254 164200 273260 164212
rect 252428 164172 273260 164200
rect 252428 164160 252434 164172
rect 273254 164160 273260 164172
rect 273312 164160 273318 164212
rect 324406 164160 324412 164212
rect 324464 164200 324470 164212
rect 338206 164200 338212 164212
rect 324464 164172 338212 164200
rect 324464 164160 324470 164172
rect 338206 164160 338212 164172
rect 338264 164160 338270 164212
rect 496998 164160 497004 164212
rect 497056 164200 497062 164212
rect 517606 164200 517612 164212
rect 497056 164172 517612 164200
rect 497056 164160 497062 164172
rect 517606 164160 517612 164172
rect 517664 164200 517670 164212
rect 546494 164200 546500 164212
rect 517664 164172 546500 164200
rect 517664 164160 517670 164172
rect 546494 164160 546500 164172
rect 546552 164160 546558 164212
rect 252278 164092 252284 164144
rect 252336 164132 252342 164144
rect 270494 164132 270500 164144
rect 252336 164104 270500 164132
rect 252336 164092 252342 164104
rect 270494 164092 270500 164104
rect 270552 164092 270558 164144
rect 324314 164092 324320 164144
rect 324372 164132 324378 164144
rect 331490 164132 331496 164144
rect 324372 164104 331496 164132
rect 324372 164092 324378 164104
rect 331490 164092 331496 164104
rect 331548 164092 331554 164144
rect 252462 164024 252468 164076
rect 252520 164064 252526 164076
rect 269298 164064 269304 164076
rect 252520 164036 269304 164064
rect 252520 164024 252526 164036
rect 269298 164024 269304 164036
rect 269356 164024 269362 164076
rect 253290 163480 253296 163532
rect 253348 163520 253354 163532
rect 267918 163520 267924 163532
rect 253348 163492 267924 163520
rect 253348 163480 253354 163492
rect 267918 163480 267924 163492
rect 267976 163480 267982 163532
rect 268378 163480 268384 163532
rect 268436 163520 268442 163532
rect 307478 163520 307484 163532
rect 268436 163492 307484 163520
rect 268436 163480 268442 163492
rect 307478 163480 307484 163492
rect 307536 163480 307542 163532
rect 304350 163004 304356 163056
rect 304408 163044 304414 163056
rect 307662 163044 307668 163056
rect 304408 163016 307668 163044
rect 304408 163004 304414 163016
rect 307662 163004 307668 163016
rect 307720 163004 307726 163056
rect 298922 162936 298928 162988
rect 298980 162976 298986 162988
rect 307570 162976 307576 162988
rect 298980 162948 307576 162976
rect 298980 162936 298986 162948
rect 307570 162936 307576 162948
rect 307628 162936 307634 162988
rect 261662 162868 261668 162920
rect 261720 162908 261726 162920
rect 307110 162908 307116 162920
rect 261720 162880 307116 162908
rect 261720 162868 261726 162880
rect 307110 162868 307116 162880
rect 307168 162868 307174 162920
rect 169018 162800 169024 162852
rect 169076 162840 169082 162852
rect 213914 162840 213920 162852
rect 169076 162812 213920 162840
rect 169076 162800 169082 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 252370 162800 252376 162852
rect 252428 162840 252434 162852
rect 266446 162840 266452 162852
rect 252428 162812 266452 162840
rect 252428 162800 252434 162812
rect 266446 162800 266452 162812
rect 266504 162800 266510 162852
rect 324314 162800 324320 162852
rect 324372 162840 324378 162852
rect 342438 162840 342444 162852
rect 324372 162812 342444 162840
rect 324372 162800 324378 162812
rect 342438 162800 342444 162812
rect 342496 162800 342502 162852
rect 496998 162800 497004 162852
rect 497056 162840 497062 162852
rect 508498 162840 508504 162852
rect 497056 162812 508504 162840
rect 497056 162800 497062 162812
rect 508498 162800 508504 162812
rect 508556 162800 508562 162852
rect 252462 162732 252468 162784
rect 252520 162772 252526 162784
rect 265066 162772 265072 162784
rect 252520 162744 265072 162772
rect 252520 162732 252526 162744
rect 265066 162732 265072 162744
rect 265124 162732 265130 162784
rect 324406 162732 324412 162784
rect 324464 162772 324470 162784
rect 335446 162772 335452 162784
rect 324464 162744 335452 162772
rect 324464 162732 324470 162744
rect 335446 162732 335452 162744
rect 335504 162732 335510 162784
rect 250438 162188 250444 162240
rect 250496 162228 250502 162240
rect 258258 162228 258264 162240
rect 250496 162200 258264 162228
rect 250496 162188 250502 162200
rect 258258 162188 258264 162200
rect 258316 162188 258322 162240
rect 250530 162120 250536 162172
rect 250588 162160 250594 162172
rect 260926 162160 260932 162172
rect 250588 162132 260932 162160
rect 250588 162120 250594 162132
rect 260926 162120 260932 162132
rect 260984 162120 260990 162172
rect 296070 161576 296076 161628
rect 296128 161616 296134 161628
rect 307570 161616 307576 161628
rect 296128 161588 307576 161616
rect 296128 161576 296134 161588
rect 307570 161576 307576 161588
rect 307628 161576 307634 161628
rect 272702 161508 272708 161560
rect 272760 161548 272766 161560
rect 307662 161548 307668 161560
rect 272760 161520 307668 161548
rect 272760 161508 272766 161520
rect 307662 161508 307668 161520
rect 307720 161508 307726 161560
rect 261478 161440 261484 161492
rect 261536 161480 261542 161492
rect 307294 161480 307300 161492
rect 261536 161452 307300 161480
rect 261536 161440 261542 161452
rect 307294 161440 307300 161452
rect 307352 161440 307358 161492
rect 342898 161440 342904 161492
rect 342956 161480 342962 161492
rect 416774 161480 416780 161492
rect 342956 161452 416780 161480
rect 342956 161440 342962 161452
rect 416774 161440 416780 161452
rect 416832 161440 416838 161492
rect 169202 161372 169208 161424
rect 169260 161412 169266 161424
rect 213914 161412 213920 161424
rect 169260 161384 213920 161412
rect 169260 161372 169266 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 252462 161372 252468 161424
rect 252520 161412 252526 161424
rect 271966 161412 271972 161424
rect 252520 161384 271972 161412
rect 252520 161372 252526 161384
rect 271966 161372 271972 161384
rect 272024 161372 272030 161424
rect 324314 161372 324320 161424
rect 324372 161412 324378 161424
rect 340874 161412 340880 161424
rect 324372 161384 340880 161412
rect 324372 161372 324378 161384
rect 340874 161372 340880 161384
rect 340932 161372 340938 161424
rect 496998 161372 497004 161424
rect 497056 161412 497062 161424
rect 515398 161412 515404 161424
rect 497056 161384 515404 161412
rect 497056 161372 497062 161384
rect 515398 161372 515404 161384
rect 515456 161372 515462 161424
rect 283742 160692 283748 160744
rect 283800 160732 283806 160744
rect 307386 160732 307392 160744
rect 283800 160704 307392 160732
rect 283800 160692 283806 160704
rect 307386 160692 307392 160704
rect 307444 160692 307450 160744
rect 263042 160148 263048 160200
rect 263100 160188 263106 160200
rect 307570 160188 307576 160200
rect 263100 160160 307576 160188
rect 263100 160148 263106 160160
rect 307570 160148 307576 160160
rect 307628 160148 307634 160200
rect 258994 160080 259000 160132
rect 259052 160120 259058 160132
rect 307662 160120 307668 160132
rect 259052 160092 307668 160120
rect 259052 160080 259058 160092
rect 307662 160080 307668 160092
rect 307720 160080 307726 160132
rect 169294 160012 169300 160064
rect 169352 160052 169358 160064
rect 214006 160052 214012 160064
rect 169352 160024 214012 160052
rect 169352 160012 169358 160024
rect 214006 160012 214012 160024
rect 214064 160012 214070 160064
rect 252462 160012 252468 160064
rect 252520 160052 252526 160064
rect 269206 160052 269212 160064
rect 252520 160024 269212 160052
rect 252520 160012 252526 160024
rect 269206 160012 269212 160024
rect 269264 160012 269270 160064
rect 324314 160012 324320 160064
rect 324372 160052 324378 160064
rect 334158 160052 334164 160064
rect 324372 160024 334164 160052
rect 324372 160012 324378 160024
rect 334158 160012 334164 160024
rect 334216 160012 334222 160064
rect 496998 160012 497004 160064
rect 497056 160052 497062 160064
rect 511994 160052 512000 160064
rect 497056 160024 512000 160052
rect 497056 160012 497062 160024
rect 511994 160012 512000 160024
rect 512052 160012 512058 160064
rect 195330 159944 195336 159996
rect 195388 159984 195394 159996
rect 213914 159984 213920 159996
rect 195388 159956 213920 159984
rect 195388 159944 195394 159956
rect 213914 159944 213920 159956
rect 213972 159944 213978 159996
rect 251726 159944 251732 159996
rect 251784 159984 251790 159996
rect 254118 159984 254124 159996
rect 251784 159956 254124 159984
rect 251784 159944 251790 159956
rect 254118 159944 254124 159956
rect 254176 159944 254182 159996
rect 497090 159944 497096 159996
rect 497148 159984 497154 159996
rect 504358 159984 504364 159996
rect 497148 159956 504364 159984
rect 497148 159944 497154 159956
rect 504358 159944 504364 159956
rect 504416 159944 504422 159996
rect 250622 159400 250628 159452
rect 250680 159440 250686 159452
rect 259730 159440 259736 159452
rect 250680 159412 259736 159440
rect 250680 159400 250686 159412
rect 259730 159400 259736 159412
rect 259788 159400 259794 159452
rect 253474 159332 253480 159384
rect 253532 159372 253538 159384
rect 258166 159372 258172 159384
rect 253532 159344 258172 159372
rect 253532 159332 253538 159344
rect 258166 159332 258172 159344
rect 258224 159332 258230 159384
rect 292022 158856 292028 158908
rect 292080 158896 292086 158908
rect 307110 158896 307116 158908
rect 292080 158868 307116 158896
rect 292080 158856 292086 158868
rect 307110 158856 307116 158868
rect 307168 158856 307174 158908
rect 265710 158788 265716 158840
rect 265768 158828 265774 158840
rect 307662 158828 307668 158840
rect 265768 158800 307668 158828
rect 265768 158788 265774 158800
rect 307662 158788 307668 158800
rect 307720 158788 307726 158840
rect 260190 158720 260196 158772
rect 260248 158760 260254 158772
rect 306742 158760 306748 158772
rect 260248 158732 306748 158760
rect 260248 158720 260254 158732
rect 306742 158720 306748 158732
rect 306800 158720 306806 158772
rect 335998 158720 336004 158772
rect 336056 158760 336062 158772
rect 416774 158760 416780 158772
rect 336056 158732 416780 158760
rect 336056 158720 336062 158732
rect 416774 158720 416780 158732
rect 416832 158720 416838 158772
rect 169110 158652 169116 158704
rect 169168 158692 169174 158704
rect 213914 158692 213920 158704
rect 169168 158664 213920 158692
rect 169168 158652 169174 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 252462 158652 252468 158704
rect 252520 158692 252526 158704
rect 261018 158692 261024 158704
rect 252520 158664 261024 158692
rect 252520 158652 252526 158664
rect 261018 158652 261024 158664
rect 261076 158652 261082 158704
rect 324406 158652 324412 158704
rect 324464 158692 324470 158704
rect 343818 158692 343824 158704
rect 324464 158664 343824 158692
rect 324464 158652 324470 158664
rect 343818 158652 343824 158664
rect 343876 158652 343882 158704
rect 496998 158652 497004 158704
rect 497056 158692 497062 158704
rect 519538 158692 519544 158704
rect 497056 158664 519544 158692
rect 497056 158652 497062 158664
rect 519538 158652 519544 158664
rect 519596 158652 519602 158704
rect 324314 158584 324320 158636
rect 324372 158624 324378 158636
rect 331398 158624 331404 158636
rect 324372 158596 331404 158624
rect 324372 158584 324378 158596
rect 331398 158584 331404 158596
rect 331456 158584 331462 158636
rect 251818 158040 251824 158092
rect 251876 158080 251882 158092
rect 259454 158080 259460 158092
rect 251876 158052 259460 158080
rect 251876 158040 251882 158052
rect 259454 158040 259460 158052
rect 259512 158040 259518 158092
rect 300210 157496 300216 157548
rect 300268 157536 300274 157548
rect 306558 157536 306564 157548
rect 300268 157508 306564 157536
rect 300268 157496 300274 157508
rect 306558 157496 306564 157508
rect 306616 157496 306622 157548
rect 276750 157428 276756 157480
rect 276808 157468 276814 157480
rect 307662 157468 307668 157480
rect 276808 157440 307668 157468
rect 276808 157428 276814 157440
rect 307662 157428 307668 157440
rect 307720 157428 307726 157480
rect 258810 157360 258816 157412
rect 258868 157400 258874 157412
rect 307570 157400 307576 157412
rect 258868 157372 307576 157400
rect 258868 157360 258874 157372
rect 307570 157360 307576 157372
rect 307628 157360 307634 157412
rect 341518 157360 341524 157412
rect 341576 157400 341582 157412
rect 416774 157400 416780 157412
rect 341576 157372 416780 157400
rect 341576 157360 341582 157372
rect 416774 157360 416780 157372
rect 416832 157360 416838 157412
rect 170490 157292 170496 157344
rect 170548 157332 170554 157344
rect 214006 157332 214012 157344
rect 170548 157304 214012 157332
rect 170548 157292 170554 157304
rect 214006 157292 214012 157304
rect 214064 157292 214070 157344
rect 252462 157292 252468 157344
rect 252520 157332 252526 157344
rect 262398 157332 262404 157344
rect 252520 157304 262404 157332
rect 252520 157292 252526 157304
rect 262398 157292 262404 157304
rect 262456 157292 262462 157344
rect 324314 157292 324320 157344
rect 324372 157332 324378 157344
rect 336826 157332 336832 157344
rect 324372 157304 336832 157332
rect 324372 157292 324378 157304
rect 336826 157292 336832 157304
rect 336884 157292 336890 157344
rect 496998 157292 497004 157344
rect 497056 157332 497062 157344
rect 582374 157332 582380 157344
rect 497056 157304 582380 157332
rect 497056 157292 497062 157304
rect 582374 157292 582380 157304
rect 582432 157292 582438 157344
rect 173158 157224 173164 157276
rect 173216 157264 173222 157276
rect 213914 157264 213920 157276
rect 173216 157236 213920 157264
rect 173216 157224 173222 157236
rect 213914 157224 213920 157236
rect 213972 157224 213978 157276
rect 324314 156816 324320 156868
rect 324372 156856 324378 156868
rect 327350 156856 327356 156868
rect 324372 156828 327356 156856
rect 324372 156816 324378 156828
rect 327350 156816 327356 156828
rect 327408 156816 327414 156868
rect 285214 156068 285220 156120
rect 285272 156108 285278 156120
rect 307662 156108 307668 156120
rect 285272 156080 307668 156108
rect 285272 156068 285278 156080
rect 307662 156068 307668 156080
rect 307720 156068 307726 156120
rect 271230 156000 271236 156052
rect 271288 156040 271294 156052
rect 307478 156040 307484 156052
rect 271288 156012 307484 156040
rect 271288 156000 271294 156012
rect 307478 156000 307484 156012
rect 307536 156000 307542 156052
rect 261570 155932 261576 155984
rect 261628 155972 261634 155984
rect 307570 155972 307576 155984
rect 261628 155944 307576 155972
rect 261628 155932 261634 155944
rect 307570 155932 307576 155944
rect 307628 155932 307634 155984
rect 352558 155932 352564 155984
rect 352616 155972 352622 155984
rect 416774 155972 416780 155984
rect 352616 155944 416780 155972
rect 352616 155932 352622 155944
rect 416774 155932 416780 155944
rect 416832 155932 416838 155984
rect 170582 155864 170588 155916
rect 170640 155904 170646 155916
rect 213914 155904 213920 155916
rect 170640 155876 213920 155904
rect 170640 155864 170646 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 252370 155864 252376 155916
rect 252428 155904 252434 155916
rect 270678 155904 270684 155916
rect 252428 155876 270684 155904
rect 252428 155864 252434 155876
rect 270678 155864 270684 155876
rect 270736 155864 270742 155916
rect 324406 155864 324412 155916
rect 324464 155904 324470 155916
rect 345290 155904 345296 155916
rect 324464 155876 345296 155904
rect 324464 155864 324470 155876
rect 345290 155864 345296 155876
rect 345348 155864 345354 155916
rect 496998 155864 497004 155916
rect 497056 155904 497062 155916
rect 511258 155904 511264 155916
rect 497056 155876 511264 155904
rect 497056 155864 497062 155876
rect 511258 155864 511264 155876
rect 511316 155864 511322 155916
rect 252462 155796 252468 155848
rect 252520 155836 252526 155848
rect 264974 155836 264980 155848
rect 252520 155808 264980 155836
rect 252520 155796 252526 155808
rect 264974 155796 264980 155808
rect 265032 155796 265038 155848
rect 324314 155796 324320 155848
rect 324372 155836 324378 155848
rect 339678 155836 339684 155848
rect 324372 155808 339684 155836
rect 324372 155796 324378 155808
rect 339678 155796 339684 155808
rect 339736 155796 339742 155848
rect 253934 155184 253940 155236
rect 253992 155224 253998 155236
rect 268010 155224 268016 155236
rect 253992 155196 268016 155224
rect 253992 155184 253998 155196
rect 268010 155184 268016 155196
rect 268068 155184 268074 155236
rect 274082 155184 274088 155236
rect 274140 155224 274146 155236
rect 307386 155224 307392 155236
rect 274140 155196 307392 155224
rect 274140 155184 274146 155196
rect 307386 155184 307392 155196
rect 307444 155184 307450 155236
rect 286594 154640 286600 154692
rect 286652 154680 286658 154692
rect 307662 154680 307668 154692
rect 286652 154652 307668 154680
rect 286652 154640 286658 154652
rect 307662 154640 307668 154652
rect 307720 154640 307726 154692
rect 264330 154572 264336 154624
rect 264388 154612 264394 154624
rect 306558 154612 306564 154624
rect 264388 154584 306564 154612
rect 264388 154572 264394 154584
rect 306558 154572 306564 154584
rect 306616 154572 306622 154624
rect 356790 154572 356796 154624
rect 356848 154612 356854 154624
rect 416774 154612 416780 154624
rect 356848 154584 416780 154612
rect 356848 154572 356854 154584
rect 416774 154572 416780 154584
rect 416832 154572 416838 154624
rect 252462 154504 252468 154556
rect 252520 154544 252526 154556
rect 273346 154544 273352 154556
rect 252520 154516 273352 154544
rect 252520 154504 252526 154516
rect 273346 154504 273352 154516
rect 273404 154504 273410 154556
rect 496998 154504 497004 154556
rect 497056 154544 497062 154556
rect 502518 154544 502524 154556
rect 497056 154516 502524 154544
rect 497056 154504 497062 154516
rect 502518 154504 502524 154516
rect 502576 154504 502582 154556
rect 252094 154436 252100 154488
rect 252152 154476 252158 154488
rect 255406 154476 255412 154488
rect 252152 154448 255412 154476
rect 252152 154436 252158 154448
rect 255406 154436 255412 154448
rect 255464 154436 255470 154488
rect 324406 154436 324412 154488
rect 324464 154476 324470 154488
rect 328638 154476 328644 154488
rect 324464 154448 328644 154476
rect 324464 154436 324470 154448
rect 328638 154436 328644 154448
rect 328696 154436 328702 154488
rect 497090 154436 497096 154488
rect 497148 154476 497154 154488
rect 502610 154476 502616 154488
rect 497148 154448 502616 154476
rect 497148 154436 497154 154448
rect 502610 154436 502616 154448
rect 502668 154436 502674 154488
rect 324314 154300 324320 154352
rect 324372 154340 324378 154352
rect 325970 154340 325976 154352
rect 324372 154312 325976 154340
rect 324372 154300 324378 154312
rect 325970 154300 325976 154312
rect 326028 154300 326034 154352
rect 256234 153824 256240 153876
rect 256292 153864 256298 153876
rect 307294 153864 307300 153876
rect 256292 153836 307300 153864
rect 256292 153824 256298 153836
rect 307294 153824 307300 153836
rect 307352 153824 307358 153876
rect 191282 153280 191288 153332
rect 191340 153320 191346 153332
rect 213914 153320 213920 153332
rect 191340 153292 213920 153320
rect 191340 153280 191346 153292
rect 213914 153280 213920 153292
rect 213972 153280 213978 153332
rect 301590 153280 301596 153332
rect 301648 153320 301654 153332
rect 307662 153320 307668 153332
rect 301648 153292 307668 153320
rect 301648 153280 301654 153292
rect 307662 153280 307668 153292
rect 307720 153280 307726 153332
rect 178862 153212 178868 153264
rect 178920 153252 178926 153264
rect 214006 153252 214012 153264
rect 178920 153224 214012 153252
rect 178920 153212 178926 153224
rect 214006 153212 214012 153224
rect 214064 153212 214070 153264
rect 268470 153212 268476 153264
rect 268528 153252 268534 153264
rect 306926 153252 306932 153264
rect 268528 153224 306932 153252
rect 268528 153212 268534 153224
rect 306926 153212 306932 153224
rect 306984 153212 306990 153264
rect 359458 153212 359464 153264
rect 359516 153252 359522 153264
rect 416774 153252 416780 153264
rect 359516 153224 416780 153252
rect 359516 153212 359522 153224
rect 416774 153212 416780 153224
rect 416832 153212 416838 153264
rect 252278 153144 252284 153196
rect 252336 153184 252342 153196
rect 253934 153184 253940 153196
rect 252336 153156 253940 153184
rect 252336 153144 252342 153156
rect 253934 153144 253940 153156
rect 253992 153144 253998 153196
rect 324314 153144 324320 153196
rect 324372 153184 324378 153196
rect 341150 153184 341156 153196
rect 324372 153156 341156 153184
rect 324372 153144 324378 153156
rect 341150 153144 341156 153156
rect 341208 153144 341214 153196
rect 496998 153144 497004 153196
rect 497056 153184 497062 153196
rect 505186 153184 505192 153196
rect 497056 153156 505192 153184
rect 497056 153144 497062 153156
rect 505186 153144 505192 153156
rect 505244 153144 505250 153196
rect 574738 153144 574744 153196
rect 574796 153184 574802 153196
rect 579798 153184 579804 153196
rect 574796 153156 579804 153184
rect 574796 153144 574802 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 252370 153076 252376 153128
rect 252428 153116 252434 153128
rect 274726 153116 274732 153128
rect 252428 153088 274732 153116
rect 252428 153076 252434 153088
rect 274726 153076 274732 153088
rect 274784 153076 274790 153128
rect 252462 153008 252468 153060
rect 252520 153048 252526 153060
rect 276198 153048 276204 153060
rect 252520 153020 276204 153048
rect 252520 153008 252526 153020
rect 276198 153008 276204 153020
rect 276256 153008 276262 153060
rect 299106 152532 299112 152584
rect 299164 152572 299170 152584
rect 307662 152572 307668 152584
rect 299164 152544 307668 152572
rect 299164 152532 299170 152544
rect 307662 152532 307668 152544
rect 307720 152532 307726 152584
rect 253198 152464 253204 152516
rect 253256 152504 253262 152516
rect 307478 152504 307484 152516
rect 253256 152476 307484 152504
rect 253256 152464 253262 152476
rect 307478 152464 307484 152476
rect 307536 152464 307542 152516
rect 173158 151920 173164 151972
rect 173216 151960 173222 151972
rect 214006 151960 214012 151972
rect 173216 151932 214012 151960
rect 173216 151920 173222 151932
rect 214006 151920 214012 151932
rect 214064 151920 214070 151972
rect 189718 151852 189724 151904
rect 189776 151892 189782 151904
rect 213914 151892 213920 151904
rect 189776 151864 213920 151892
rect 189776 151852 189782 151864
rect 213914 151852 213920 151864
rect 213972 151852 213978 151904
rect 257430 151784 257436 151836
rect 257488 151824 257494 151836
rect 307110 151824 307116 151836
rect 257488 151796 307116 151824
rect 257488 151784 257494 151796
rect 307110 151784 307116 151796
rect 307168 151784 307174 151836
rect 252462 151716 252468 151768
rect 252520 151756 252526 151768
rect 254026 151756 254032 151768
rect 252520 151728 254032 151756
rect 252520 151716 252526 151728
rect 254026 151716 254032 151728
rect 254084 151716 254090 151768
rect 324314 151716 324320 151768
rect 324372 151756 324378 151768
rect 338298 151756 338304 151768
rect 324372 151728 338304 151756
rect 324372 151716 324378 151728
rect 338298 151716 338304 151728
rect 338356 151716 338362 151768
rect 496998 151716 497004 151768
rect 497056 151756 497062 151768
rect 508038 151756 508044 151768
rect 497056 151728 508044 151756
rect 497056 151716 497062 151728
rect 508038 151716 508044 151728
rect 508096 151716 508102 151768
rect 324406 151648 324412 151700
rect 324464 151688 324470 151700
rect 332594 151688 332600 151700
rect 324464 151660 332600 151688
rect 324464 151648 324470 151660
rect 332594 151648 332600 151660
rect 332652 151648 332658 151700
rect 252462 151444 252468 151496
rect 252520 151484 252526 151496
rect 255590 151484 255596 151496
rect 252520 151456 255596 151484
rect 252520 151444 252526 151456
rect 255590 151444 255596 151456
rect 255648 151444 255654 151496
rect 252278 151240 252284 151292
rect 252336 151280 252342 151292
rect 255498 151280 255504 151292
rect 252336 151252 255504 151280
rect 252336 151240 252342 151252
rect 255498 151240 255504 151252
rect 255556 151240 255562 151292
rect 167638 151036 167644 151088
rect 167696 151076 167702 151088
rect 184566 151076 184572 151088
rect 167696 151048 184572 151076
rect 167696 151036 167702 151048
rect 184566 151036 184572 151048
rect 184624 151036 184630 151088
rect 293402 150560 293408 150612
rect 293460 150600 293466 150612
rect 307662 150600 307668 150612
rect 293460 150572 307668 150600
rect 293460 150560 293466 150572
rect 307662 150560 307668 150572
rect 307720 150560 307726 150612
rect 255958 150492 255964 150544
rect 256016 150532 256022 150544
rect 307478 150532 307484 150544
rect 256016 150504 307484 150532
rect 256016 150492 256022 150504
rect 307478 150492 307484 150504
rect 307536 150492 307542 150544
rect 176010 150424 176016 150476
rect 176068 150464 176074 150476
rect 213914 150464 213920 150476
rect 176068 150436 213920 150464
rect 176068 150424 176074 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 254670 150424 254676 150476
rect 254728 150464 254734 150476
rect 307570 150464 307576 150476
rect 254728 150436 307576 150464
rect 254728 150424 254734 150436
rect 307570 150424 307576 150436
rect 307628 150424 307634 150476
rect 331858 150424 331864 150476
rect 331916 150464 331922 150476
rect 416774 150464 416780 150476
rect 331916 150436 416780 150464
rect 331916 150424 331922 150436
rect 416774 150424 416780 150436
rect 416832 150424 416838 150476
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 22738 150396 22744 150408
rect 3476 150368 22744 150396
rect 3476 150356 3482 150368
rect 22738 150356 22744 150368
rect 22796 150356 22802 150408
rect 184566 150356 184572 150408
rect 184624 150396 184630 150408
rect 214006 150396 214012 150408
rect 184624 150368 214012 150396
rect 184624 150356 184630 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 252370 150356 252376 150408
rect 252428 150396 252434 150408
rect 284294 150396 284300 150408
rect 252428 150368 284300 150396
rect 252428 150356 252434 150368
rect 284294 150356 284300 150368
rect 284352 150356 284358 150408
rect 324314 150356 324320 150408
rect 324372 150396 324378 150408
rect 336734 150396 336740 150408
rect 324372 150368 336740 150396
rect 324372 150356 324378 150368
rect 336734 150356 336740 150368
rect 336792 150356 336798 150408
rect 496998 150356 497004 150408
rect 497056 150396 497062 150408
rect 501230 150396 501236 150408
rect 497056 150368 501236 150396
rect 497056 150356 497062 150368
rect 501230 150356 501236 150368
rect 501288 150356 501294 150408
rect 209130 150288 209136 150340
rect 209188 150328 209194 150340
rect 213914 150328 213920 150340
rect 209188 150300 213920 150328
rect 209188 150288 209194 150300
rect 213914 150288 213920 150300
rect 213972 150288 213978 150340
rect 252462 150288 252468 150340
rect 252520 150328 252526 150340
rect 280154 150328 280160 150340
rect 252520 150300 280160 150328
rect 252520 150288 252526 150300
rect 280154 150288 280160 150300
rect 280212 150288 280218 150340
rect 252278 150220 252284 150272
rect 252336 150260 252342 150272
rect 256786 150260 256792 150272
rect 252336 150232 256792 150260
rect 252336 150220 252342 150232
rect 256786 150220 256792 150232
rect 256844 150220 256850 150272
rect 324314 149744 324320 149796
rect 324372 149784 324378 149796
rect 327258 149784 327264 149796
rect 324372 149756 327264 149784
rect 324372 149744 324378 149756
rect 327258 149744 327264 149756
rect 327316 149744 327322 149796
rect 281074 149676 281080 149728
rect 281132 149716 281138 149728
rect 306650 149716 306656 149728
rect 281132 149688 306656 149716
rect 281132 149676 281138 149688
rect 306650 149676 306656 149688
rect 306708 149676 306714 149728
rect 275554 149132 275560 149184
rect 275612 149172 275618 149184
rect 307570 149172 307576 149184
rect 275612 149144 307576 149172
rect 275612 149132 275618 149144
rect 307570 149132 307576 149144
rect 307628 149132 307634 149184
rect 267274 149064 267280 149116
rect 267332 149104 267338 149116
rect 307662 149104 307668 149116
rect 267332 149076 307668 149104
rect 267332 149064 267338 149076
rect 307662 149064 307668 149076
rect 307720 149064 307726 149116
rect 363598 149064 363604 149116
rect 363656 149104 363662 149116
rect 416774 149104 416780 149116
rect 363656 149076 416780 149104
rect 363656 149064 363662 149076
rect 416774 149064 416780 149076
rect 416832 149064 416838 149116
rect 211890 148996 211896 149048
rect 211948 149036 211954 149048
rect 213914 149036 213920 149048
rect 211948 149008 213920 149036
rect 211948 148996 211954 149008
rect 213914 148996 213920 149008
rect 213972 148996 213978 149048
rect 252462 148996 252468 149048
rect 252520 149036 252526 149048
rect 281534 149036 281540 149048
rect 252520 149008 281540 149036
rect 252520 148996 252526 149008
rect 281534 148996 281540 149008
rect 281592 148996 281598 149048
rect 324314 148996 324320 149048
rect 324372 149036 324378 149048
rect 349246 149036 349252 149048
rect 324372 149008 349252 149036
rect 324372 148996 324378 149008
rect 349246 148996 349252 149008
rect 349304 148996 349310 149048
rect 496998 148996 497004 149048
rect 497056 149036 497062 149048
rect 509326 149036 509332 149048
rect 497056 149008 509332 149036
rect 497056 148996 497062 149008
rect 509326 148996 509332 149008
rect 509384 148996 509390 149048
rect 252370 148928 252376 148980
rect 252428 148968 252434 148980
rect 256694 148968 256700 148980
rect 252428 148940 256700 148968
rect 252428 148928 252434 148940
rect 256694 148928 256700 148940
rect 256752 148928 256758 148980
rect 256142 148316 256148 148368
rect 256200 148356 256206 148368
rect 306742 148356 306748 148368
rect 256200 148328 306748 148356
rect 256200 148316 256206 148328
rect 306742 148316 306748 148328
rect 306800 148316 306806 148368
rect 182910 147636 182916 147688
rect 182968 147676 182974 147688
rect 213914 147676 213920 147688
rect 182968 147648 213920 147676
rect 182968 147636 182974 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 256050 147636 256056 147688
rect 256108 147676 256114 147688
rect 307110 147676 307116 147688
rect 256108 147648 307116 147676
rect 256108 147636 256114 147648
rect 307110 147636 307116 147648
rect 307168 147636 307174 147688
rect 374638 147636 374644 147688
rect 374696 147676 374702 147688
rect 416774 147676 416780 147688
rect 374696 147648 416780 147676
rect 374696 147636 374702 147648
rect 416774 147636 416780 147648
rect 416832 147636 416838 147688
rect 252370 147568 252376 147620
rect 252428 147608 252434 147620
rect 278774 147608 278780 147620
rect 252428 147580 278780 147608
rect 252428 147568 252434 147580
rect 278774 147568 278780 147580
rect 278832 147568 278838 147620
rect 324314 147568 324320 147620
rect 324372 147608 324378 147620
rect 350534 147608 350540 147620
rect 324372 147580 350540 147608
rect 324372 147568 324378 147580
rect 350534 147568 350540 147580
rect 350592 147568 350598 147620
rect 496998 147568 497004 147620
rect 497056 147608 497062 147620
rect 505094 147608 505100 147620
rect 497056 147580 505100 147608
rect 497056 147568 497062 147580
rect 505094 147568 505100 147580
rect 505152 147568 505158 147620
rect 252462 147500 252468 147552
rect 252520 147540 252526 147552
rect 274634 147540 274640 147552
rect 252520 147512 274640 147540
rect 252520 147500 252526 147512
rect 274634 147500 274640 147512
rect 274692 147500 274698 147552
rect 251450 147432 251456 147484
rect 251508 147472 251514 147484
rect 254210 147472 254216 147484
rect 251508 147444 254216 147472
rect 251508 147432 251514 147444
rect 254210 147432 254216 147444
rect 254268 147432 254274 147484
rect 325786 147024 325792 147076
rect 325844 147024 325850 147076
rect 325694 146820 325700 146872
rect 325752 146860 325758 146872
rect 325804 146860 325832 147024
rect 325752 146832 325832 146860
rect 325752 146820 325758 146832
rect 254854 146480 254860 146532
rect 254912 146520 254918 146532
rect 307662 146520 307668 146532
rect 254912 146492 307668 146520
rect 254912 146480 254918 146492
rect 307662 146480 307668 146492
rect 307720 146480 307726 146532
rect 276842 146412 276848 146464
rect 276900 146452 276906 146464
rect 307570 146452 307576 146464
rect 276900 146424 307576 146452
rect 276900 146412 276906 146424
rect 307570 146412 307576 146424
rect 307628 146412 307634 146464
rect 185578 146344 185584 146396
rect 185636 146384 185642 146396
rect 214006 146384 214012 146396
rect 185636 146356 214012 146384
rect 185636 146344 185642 146356
rect 214006 146344 214012 146356
rect 214064 146344 214070 146396
rect 257522 146344 257528 146396
rect 257580 146384 257586 146396
rect 307662 146384 307668 146396
rect 257580 146356 307668 146384
rect 257580 146344 257586 146356
rect 307662 146344 307668 146356
rect 307720 146344 307726 146396
rect 171778 146276 171784 146328
rect 171836 146316 171842 146328
rect 213914 146316 213920 146328
rect 171836 146288 213920 146316
rect 171836 146276 171842 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 303614 146276 303620 146328
rect 303672 146316 303678 146328
rect 307478 146316 307484 146328
rect 303672 146288 307484 146316
rect 303672 146276 303678 146288
rect 307478 146276 307484 146288
rect 307536 146276 307542 146328
rect 334710 146276 334716 146328
rect 334768 146316 334774 146328
rect 416774 146316 416780 146328
rect 334768 146288 416780 146316
rect 334768 146276 334774 146288
rect 416774 146276 416780 146288
rect 416832 146276 416838 146328
rect 252462 146208 252468 146260
rect 252520 146248 252526 146260
rect 271874 146248 271880 146260
rect 252520 146220 271880 146248
rect 252520 146208 252526 146220
rect 271874 146208 271880 146220
rect 271932 146208 271938 146260
rect 324314 146208 324320 146260
rect 324372 146248 324378 146260
rect 353386 146248 353392 146260
rect 324372 146220 353392 146248
rect 324372 146208 324378 146220
rect 353386 146208 353392 146220
rect 353444 146208 353450 146260
rect 525794 146208 525800 146260
rect 525852 146248 525858 146260
rect 580258 146248 580264 146260
rect 525852 146220 580264 146248
rect 525852 146208 525858 146220
rect 580258 146208 580264 146220
rect 580316 146208 580322 146260
rect 252370 146140 252376 146192
rect 252428 146180 252434 146192
rect 267826 146180 267832 146192
rect 252428 146152 267832 146180
rect 252428 146140 252434 146152
rect 267826 146140 267832 146152
rect 267884 146140 267890 146192
rect 324406 146140 324412 146192
rect 324464 146180 324470 146192
rect 346486 146180 346492 146192
rect 324464 146152 346492 146180
rect 324464 146140 324470 146152
rect 346486 146140 346492 146152
rect 346544 146140 346550 146192
rect 251174 146072 251180 146124
rect 251232 146112 251238 146124
rect 253474 146112 253480 146124
rect 251232 146084 253480 146112
rect 251232 146072 251238 146084
rect 253474 146072 253480 146084
rect 253532 146072 253538 146124
rect 213362 145664 213368 145716
rect 213420 145704 213426 145716
rect 215018 145704 215024 145716
rect 213420 145676 215024 145704
rect 213420 145664 213426 145676
rect 215018 145664 215024 145676
rect 215076 145664 215082 145716
rect 253382 145528 253388 145580
rect 253440 145568 253446 145580
rect 306834 145568 306840 145580
rect 253440 145540 306840 145568
rect 253440 145528 253446 145540
rect 306834 145528 306840 145540
rect 306892 145528 306898 145580
rect 502978 145528 502984 145580
rect 503036 145568 503042 145580
rect 525794 145568 525800 145580
rect 503036 145540 525800 145568
rect 503036 145528 503042 145540
rect 525794 145528 525800 145540
rect 525852 145528 525858 145580
rect 292114 144916 292120 144968
rect 292172 144956 292178 144968
rect 306558 144956 306564 144968
rect 292172 144928 306564 144956
rect 292172 144916 292178 144928
rect 306558 144916 306564 144928
rect 306616 144916 306622 144968
rect 496998 144916 497004 144968
rect 497056 144956 497062 144968
rect 502334 144956 502340 144968
rect 497056 144928 502340 144956
rect 497056 144916 497062 144928
rect 502334 144916 502340 144928
rect 502392 144916 502398 144968
rect 252462 144848 252468 144900
rect 252520 144888 252526 144900
rect 260834 144888 260840 144900
rect 252520 144860 260840 144888
rect 252520 144848 252526 144860
rect 260834 144848 260840 144860
rect 260892 144848 260898 144900
rect 324314 144848 324320 144900
rect 324372 144888 324378 144900
rect 335354 144888 335360 144900
rect 324372 144860 335360 144888
rect 324372 144848 324378 144860
rect 335354 144848 335360 144860
rect 335412 144848 335418 144900
rect 252094 144304 252100 144356
rect 252152 144344 252158 144356
rect 268562 144344 268568 144356
rect 252152 144316 268568 144344
rect 252152 144304 252158 144316
rect 268562 144304 268568 144316
rect 268620 144304 268626 144356
rect 267182 144236 267188 144288
rect 267240 144276 267246 144288
rect 307386 144276 307392 144288
rect 267240 144248 307392 144276
rect 267240 144236 267246 144248
rect 307386 144236 307392 144248
rect 307444 144236 307450 144288
rect 250714 144168 250720 144220
rect 250772 144208 250778 144220
rect 303614 144208 303620 144220
rect 250772 144180 303620 144208
rect 250772 144168 250778 144180
rect 303614 144168 303620 144180
rect 303672 144168 303678 144220
rect 508038 144168 508044 144220
rect 508096 144208 508102 144220
rect 509142 144208 509148 144220
rect 508096 144180 509148 144208
rect 508096 144168 508102 144180
rect 509142 144168 509148 144180
rect 509200 144208 509206 144220
rect 512086 144208 512092 144220
rect 509200 144180 512092 144208
rect 509200 144168 509206 144180
rect 512086 144168 512092 144180
rect 512144 144168 512150 144220
rect 307018 144100 307024 144152
rect 307076 144140 307082 144152
rect 307386 144140 307392 144152
rect 307076 144112 307392 144140
rect 307076 144100 307082 144112
rect 307386 144100 307392 144112
rect 307444 144100 307450 144152
rect 170490 143624 170496 143676
rect 170548 143664 170554 143676
rect 213914 143664 213920 143676
rect 170548 143636 213920 143664
rect 170548 143624 170554 143636
rect 213914 143624 213920 143636
rect 213972 143624 213978 143676
rect 302970 143624 302976 143676
rect 303028 143664 303034 143676
rect 306558 143664 306564 143676
rect 303028 143636 306564 143664
rect 303028 143624 303034 143636
rect 306558 143624 306564 143636
rect 306616 143624 306622 143676
rect 169018 143556 169024 143608
rect 169076 143596 169082 143608
rect 214006 143596 214012 143608
rect 169076 143568 214012 143596
rect 169076 143556 169082 143568
rect 214006 143556 214012 143568
rect 214064 143556 214070 143608
rect 290642 143556 290648 143608
rect 290700 143596 290706 143608
rect 307662 143596 307668 143608
rect 290700 143568 307668 143596
rect 290700 143556 290706 143568
rect 307662 143556 307668 143568
rect 307720 143556 307726 143608
rect 358078 143556 358084 143608
rect 358136 143596 358142 143608
rect 416774 143596 416780 143608
rect 358136 143568 416780 143596
rect 358136 143556 358142 143568
rect 416774 143556 416780 143568
rect 416832 143556 416838 143608
rect 497090 143556 497096 143608
rect 497148 143596 497154 143608
rect 508038 143596 508044 143608
rect 497148 143568 508044 143596
rect 497148 143556 497154 143568
rect 508038 143556 508044 143568
rect 508096 143556 508102 143608
rect 252462 143488 252468 143540
rect 252520 143528 252526 143540
rect 270586 143528 270592 143540
rect 252520 143500 270592 143528
rect 252520 143488 252526 143500
rect 270586 143488 270592 143500
rect 270644 143488 270650 143540
rect 496998 143488 497004 143540
rect 497056 143528 497062 143540
rect 513374 143528 513380 143540
rect 497056 143500 513380 143528
rect 497056 143488 497062 143500
rect 513374 143488 513380 143500
rect 513432 143488 513438 143540
rect 252370 143420 252376 143472
rect 252428 143460 252434 143472
rect 269114 143460 269120 143472
rect 252428 143432 269120 143460
rect 252428 143420 252434 143432
rect 269114 143420 269120 143432
rect 269172 143420 269178 143472
rect 324314 143420 324320 143472
rect 324372 143460 324378 143472
rect 343726 143460 343732 143472
rect 324372 143432 343732 143460
rect 324372 143420 324378 143432
rect 343726 143420 343732 143432
rect 343784 143420 343790 143472
rect 513374 143352 513380 143404
rect 513432 143392 513438 143404
rect 515398 143392 515404 143404
rect 513432 143364 515404 143392
rect 513432 143352 513438 143364
rect 515398 143352 515404 143364
rect 515456 143352 515462 143404
rect 167638 142808 167644 142860
rect 167696 142848 167702 142860
rect 213454 142848 213460 142860
rect 167696 142820 213460 142848
rect 167696 142808 167702 142820
rect 213454 142808 213460 142820
rect 213512 142808 213518 142860
rect 274174 142808 274180 142860
rect 274232 142848 274238 142860
rect 307478 142848 307484 142860
rect 274232 142820 307484 142848
rect 274232 142808 274238 142820
rect 307478 142808 307484 142820
rect 307536 142808 307542 142860
rect 289354 142196 289360 142248
rect 289412 142236 289418 142248
rect 307662 142236 307668 142248
rect 289412 142208 307668 142236
rect 289412 142196 289418 142208
rect 307662 142196 307668 142208
rect 307720 142196 307726 142248
rect 181530 142128 181536 142180
rect 181588 142168 181594 142180
rect 213914 142168 213920 142180
rect 181588 142140 213920 142168
rect 181588 142128 181594 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 254762 142128 254768 142180
rect 254820 142168 254826 142180
rect 307570 142168 307576 142180
rect 254820 142140 307576 142168
rect 254820 142128 254826 142140
rect 307570 142128 307576 142140
rect 307628 142128 307634 142180
rect 345658 142128 345664 142180
rect 345716 142168 345722 142180
rect 416774 142168 416780 142180
rect 345716 142140 416780 142168
rect 345716 142128 345722 142140
rect 416774 142128 416780 142140
rect 416832 142128 416838 142180
rect 252462 142060 252468 142112
rect 252520 142100 252526 142112
rect 262490 142100 262496 142112
rect 252520 142072 262496 142100
rect 252520 142060 252526 142072
rect 262490 142060 262496 142072
rect 262548 142060 262554 142112
rect 324314 142060 324320 142112
rect 324372 142100 324378 142112
rect 356054 142100 356060 142112
rect 324372 142072 356060 142100
rect 324372 142060 324378 142072
rect 356054 142060 356060 142072
rect 356112 142060 356118 142112
rect 496998 142060 497004 142112
rect 497056 142100 497062 142112
rect 507946 142100 507952 142112
rect 497056 142072 507952 142100
rect 497056 142060 497062 142072
rect 507946 142060 507952 142072
rect 508004 142060 508010 142112
rect 251174 141516 251180 141568
rect 251232 141556 251238 141568
rect 253290 141556 253296 141568
rect 251232 141528 253296 141556
rect 251232 141516 251238 141528
rect 253290 141516 253296 141528
rect 253348 141516 253354 141568
rect 287974 141448 287980 141500
rect 288032 141488 288038 141500
rect 306558 141488 306564 141500
rect 288032 141460 306564 141488
rect 288032 141448 288038 141460
rect 306558 141448 306564 141460
rect 306616 141448 306622 141500
rect 252002 141380 252008 141432
rect 252060 141420 252066 141432
rect 294690 141420 294696 141432
rect 252060 141392 294696 141420
rect 252060 141380 252066 141392
rect 294690 141380 294696 141392
rect 294748 141380 294754 141432
rect 496814 141380 496820 141432
rect 496872 141420 496878 141432
rect 503254 141420 503260 141432
rect 496872 141392 503260 141420
rect 496872 141380 496878 141392
rect 503254 141380 503260 141392
rect 503312 141380 503318 141432
rect 301866 140904 301872 140956
rect 301924 140944 301930 140956
rect 306926 140944 306932 140956
rect 301924 140916 306932 140944
rect 301924 140904 301930 140916
rect 306926 140904 306932 140916
rect 306984 140904 306990 140956
rect 209130 140836 209136 140888
rect 209188 140876 209194 140888
rect 214006 140876 214012 140888
rect 209188 140848 214012 140876
rect 209188 140836 209194 140848
rect 214006 140836 214012 140848
rect 214064 140836 214070 140888
rect 303246 140836 303252 140888
rect 303304 140876 303310 140888
rect 307570 140876 307576 140888
rect 303304 140848 307576 140876
rect 303304 140836 303310 140848
rect 307570 140836 307576 140848
rect 307628 140836 307634 140888
rect 174538 140768 174544 140820
rect 174596 140808 174602 140820
rect 213914 140808 213920 140820
rect 174596 140780 213920 140808
rect 174596 140768 174602 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 262950 140768 262956 140820
rect 263008 140808 263014 140820
rect 307662 140808 307668 140820
rect 263008 140780 307668 140808
rect 263008 140768 263014 140780
rect 307662 140768 307668 140780
rect 307720 140768 307726 140820
rect 333422 140768 333428 140820
rect 333480 140808 333486 140820
rect 416774 140808 416780 140820
rect 333480 140780 416780 140808
rect 333480 140768 333486 140780
rect 416774 140768 416780 140780
rect 416832 140768 416838 140820
rect 507946 140768 507952 140820
rect 508004 140808 508010 140820
rect 511258 140808 511264 140820
rect 508004 140780 511264 140808
rect 508004 140768 508010 140780
rect 511258 140768 511264 140780
rect 511316 140768 511322 140820
rect 252462 140700 252468 140752
rect 252520 140740 252526 140752
rect 277486 140740 277492 140752
rect 252520 140712 277492 140740
rect 252520 140700 252526 140712
rect 277486 140700 277492 140712
rect 277544 140700 277550 140752
rect 324314 140700 324320 140752
rect 324372 140740 324378 140752
rect 328454 140740 328460 140752
rect 324372 140712 328460 140740
rect 324372 140700 324378 140712
rect 328454 140700 328460 140712
rect 328512 140700 328518 140752
rect 496814 140700 496820 140752
rect 496872 140740 496878 140752
rect 502978 140740 502984 140752
rect 496872 140712 502984 140740
rect 496872 140700 496878 140712
rect 502978 140700 502984 140712
rect 503036 140700 503042 140752
rect 252370 140632 252376 140684
rect 252428 140672 252434 140684
rect 276014 140672 276020 140684
rect 252428 140644 276020 140672
rect 252428 140632 252434 140644
rect 276014 140632 276020 140644
rect 276072 140632 276078 140684
rect 177390 140020 177396 140072
rect 177448 140060 177454 140072
rect 214650 140060 214656 140072
rect 177448 140032 214656 140060
rect 177448 140020 177454 140032
rect 214650 140020 214656 140032
rect 214708 140020 214714 140072
rect 503254 140020 503260 140072
rect 503312 140060 503318 140072
rect 580166 140060 580172 140072
rect 503312 140032 580172 140060
rect 503312 140020 503318 140032
rect 580166 140020 580172 140032
rect 580224 140020 580230 140072
rect 251910 139952 251916 140004
rect 251968 139992 251974 140004
rect 258994 139992 259000 140004
rect 251968 139964 259000 139992
rect 251968 139952 251974 139964
rect 258994 139952 259000 139964
rect 259052 139952 259058 140004
rect 271414 139476 271420 139528
rect 271472 139516 271478 139528
rect 306558 139516 306564 139528
rect 271472 139488 306564 139516
rect 271472 139476 271478 139488
rect 306558 139476 306564 139488
rect 306616 139476 306622 139528
rect 184382 139408 184388 139460
rect 184440 139448 184446 139460
rect 213914 139448 213920 139460
rect 184440 139420 213920 139448
rect 184440 139408 184446 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 254578 139408 254584 139460
rect 254636 139448 254642 139460
rect 307662 139448 307668 139460
rect 254636 139420 307668 139448
rect 254636 139408 254642 139420
rect 307662 139408 307668 139420
rect 307720 139408 307726 139460
rect 411898 139408 411904 139460
rect 411956 139448 411962 139460
rect 416774 139448 416780 139460
rect 411956 139420 416780 139448
rect 411956 139408 411962 139420
rect 416774 139408 416780 139420
rect 416832 139408 416838 139460
rect 252462 139340 252468 139392
rect 252520 139380 252526 139392
rect 263594 139380 263600 139392
rect 252520 139352 263600 139380
rect 252520 139340 252526 139352
rect 263594 139340 263600 139352
rect 263652 139340 263658 139392
rect 324406 139340 324412 139392
rect 324464 139380 324470 139392
rect 339494 139380 339500 139392
rect 324464 139352 339500 139380
rect 324464 139340 324470 139352
rect 339494 139340 339500 139352
rect 339552 139340 339558 139392
rect 496814 139340 496820 139392
rect 496872 139380 496878 139392
rect 520918 139380 520924 139392
rect 496872 139352 520924 139380
rect 496872 139340 496878 139352
rect 520918 139340 520924 139352
rect 520976 139340 520982 139392
rect 324314 139272 324320 139324
rect 324372 139312 324378 139324
rect 334066 139312 334072 139324
rect 324372 139284 334072 139312
rect 324372 139272 324378 139284
rect 334066 139272 334072 139284
rect 334124 139272 334130 139324
rect 294874 138116 294880 138168
rect 294932 138156 294938 138168
rect 306926 138156 306932 138168
rect 294932 138128 306932 138156
rect 294932 138116 294938 138128
rect 306926 138116 306932 138128
rect 306984 138116 306990 138168
rect 195330 138048 195336 138100
rect 195388 138088 195394 138100
rect 213914 138088 213920 138100
rect 195388 138060 213920 138088
rect 195388 138048 195394 138060
rect 213914 138048 213920 138060
rect 213972 138048 213978 138100
rect 253290 138048 253296 138100
rect 253348 138088 253354 138100
rect 307662 138088 307668 138100
rect 253348 138060 307668 138088
rect 253348 138048 253354 138060
rect 307662 138048 307668 138060
rect 307720 138048 307726 138100
rect 174630 137980 174636 138032
rect 174688 138020 174694 138032
rect 214006 138020 214012 138032
rect 174688 137992 214012 138020
rect 174688 137980 174694 137992
rect 214006 137980 214012 137992
rect 214064 137980 214070 138032
rect 249058 137980 249064 138032
rect 249116 138020 249122 138032
rect 306558 138020 306564 138032
rect 249116 137992 306564 138020
rect 249116 137980 249122 137992
rect 306558 137980 306564 137992
rect 306616 137980 306622 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 15838 137952 15844 137964
rect 3292 137924 15844 137952
rect 3292 137912 3298 137924
rect 15838 137912 15844 137924
rect 15896 137912 15902 137964
rect 252462 137912 252468 137964
rect 252520 137952 252526 137964
rect 277394 137952 277400 137964
rect 252520 137924 277400 137952
rect 252520 137912 252526 137924
rect 277394 137912 277400 137924
rect 277452 137912 277458 137964
rect 324314 137912 324320 137964
rect 324372 137952 324378 137964
rect 332686 137952 332692 137964
rect 324372 137924 332692 137952
rect 324372 137912 324378 137924
rect 332686 137912 332692 137924
rect 332744 137912 332750 137964
rect 496814 137912 496820 137964
rect 496872 137952 496878 137964
rect 547874 137952 547880 137964
rect 496872 137924 547880 137952
rect 496872 137912 496878 137924
rect 547874 137912 547880 137924
rect 547932 137912 547938 137964
rect 252186 137232 252192 137284
rect 252244 137272 252250 137284
rect 260282 137272 260288 137284
rect 252244 137244 260288 137272
rect 252244 137232 252250 137244
rect 260282 137232 260288 137244
rect 260340 137232 260346 137284
rect 210418 136688 210424 136740
rect 210476 136728 210482 136740
rect 214006 136728 214012 136740
rect 210476 136700 214012 136728
rect 210476 136688 210482 136700
rect 214006 136688 214012 136700
rect 214064 136688 214070 136740
rect 260098 136688 260104 136740
rect 260156 136728 260162 136740
rect 307110 136728 307116 136740
rect 260156 136700 307116 136728
rect 260156 136688 260162 136700
rect 307110 136688 307116 136700
rect 307168 136688 307174 136740
rect 166258 136620 166264 136672
rect 166316 136660 166322 136672
rect 213914 136660 213920 136672
rect 166316 136632 213920 136660
rect 166316 136620 166322 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 250622 136620 250628 136672
rect 250680 136660 250686 136672
rect 307662 136660 307668 136672
rect 250680 136632 307668 136660
rect 250680 136620 250686 136632
rect 307662 136620 307668 136632
rect 307720 136620 307726 136672
rect 376018 136620 376024 136672
rect 376076 136660 376082 136672
rect 416774 136660 416780 136672
rect 376076 136632 416780 136660
rect 376076 136620 376082 136632
rect 416774 136620 416780 136632
rect 416832 136620 416838 136672
rect 252278 136552 252284 136604
rect 252336 136592 252342 136604
rect 302878 136592 302884 136604
rect 252336 136564 302884 136592
rect 252336 136552 252342 136564
rect 302878 136552 302884 136564
rect 302936 136552 302942 136604
rect 324314 136552 324320 136604
rect 324372 136592 324378 136604
rect 329926 136592 329932 136604
rect 324372 136564 329932 136592
rect 324372 136552 324378 136564
rect 329926 136552 329932 136564
rect 329984 136552 329990 136604
rect 496814 136552 496820 136604
rect 496872 136592 496878 136604
rect 538214 136592 538220 136604
rect 496872 136564 538220 136592
rect 496872 136552 496878 136564
rect 538214 136552 538220 136564
rect 538272 136552 538278 136604
rect 252462 136484 252468 136536
rect 252520 136524 252526 136536
rect 297450 136524 297456 136536
rect 252520 136496 297456 136524
rect 252520 136484 252526 136496
rect 297450 136484 297456 136496
rect 297508 136484 297514 136536
rect 496998 136484 497004 136536
rect 497056 136524 497062 136536
rect 506474 136524 506480 136536
rect 497056 136496 506480 136524
rect 497056 136484 497062 136496
rect 506474 136484 506480 136496
rect 506532 136484 506538 136536
rect 252370 136416 252376 136468
rect 252428 136456 252434 136468
rect 266998 136456 267004 136468
rect 252428 136428 267004 136456
rect 252428 136416 252434 136428
rect 266998 136416 267004 136428
rect 267056 136416 267062 136468
rect 268562 135872 268568 135924
rect 268620 135912 268626 135924
rect 307018 135912 307024 135924
rect 268620 135884 307024 135912
rect 268620 135872 268626 135884
rect 307018 135872 307024 135884
rect 307076 135872 307082 135924
rect 304258 135396 304264 135448
rect 304316 135436 304322 135448
rect 307478 135436 307484 135448
rect 304316 135408 307484 135436
rect 304316 135396 304322 135408
rect 307478 135396 307484 135408
rect 307536 135396 307542 135448
rect 206462 135328 206468 135380
rect 206520 135368 206526 135380
rect 213914 135368 213920 135380
rect 206520 135340 213920 135368
rect 206520 135328 206526 135340
rect 213914 135328 213920 135340
rect 213972 135328 213978 135380
rect 298830 135328 298836 135380
rect 298888 135368 298894 135380
rect 307662 135368 307668 135380
rect 298888 135340 307668 135368
rect 298888 135328 298894 135340
rect 307662 135328 307668 135340
rect 307720 135328 307726 135380
rect 171962 135260 171968 135312
rect 172020 135300 172026 135312
rect 214006 135300 214012 135312
rect 172020 135272 214012 135300
rect 172020 135260 172026 135272
rect 214006 135260 214012 135272
rect 214064 135260 214070 135312
rect 250438 135260 250444 135312
rect 250496 135300 250502 135312
rect 306558 135300 306564 135312
rect 250496 135272 306564 135300
rect 250496 135260 250502 135272
rect 306558 135260 306564 135272
rect 306616 135260 306622 135312
rect 403618 135260 403624 135312
rect 403676 135300 403682 135312
rect 416774 135300 416780 135312
rect 403676 135272 416780 135300
rect 403676 135260 403682 135272
rect 416774 135260 416780 135272
rect 416832 135260 416838 135312
rect 252462 135192 252468 135244
rect 252520 135232 252526 135244
rect 285030 135232 285036 135244
rect 252520 135204 285036 135232
rect 252520 135192 252526 135204
rect 285030 135192 285036 135204
rect 285088 135192 285094 135244
rect 336090 135192 336096 135244
rect 336148 135232 336154 135244
rect 417326 135232 417332 135244
rect 336148 135204 417332 135232
rect 336148 135192 336154 135204
rect 417326 135192 417332 135204
rect 417384 135192 417390 135244
rect 496814 135192 496820 135244
rect 496872 135232 496878 135244
rect 525058 135232 525064 135244
rect 496872 135204 525064 135232
rect 496872 135192 496878 135204
rect 525058 135192 525064 135204
rect 525116 135192 525122 135244
rect 252370 135124 252376 135176
rect 252428 135164 252434 135176
rect 271138 135164 271144 135176
rect 252428 135136 271144 135164
rect 252428 135124 252434 135136
rect 271138 135124 271144 135136
rect 271196 135124 271202 135176
rect 297450 134512 297456 134564
rect 297508 134552 297514 134564
rect 307202 134552 307208 134564
rect 297508 134524 307208 134552
rect 297508 134512 297514 134524
rect 307202 134512 307208 134524
rect 307260 134512 307266 134564
rect 282454 133968 282460 134020
rect 282512 134008 282518 134020
rect 307570 134008 307576 134020
rect 282512 133980 307576 134008
rect 282512 133968 282518 133980
rect 307570 133968 307576 133980
rect 307628 133968 307634 134020
rect 175918 133900 175924 133952
rect 175976 133940 175982 133952
rect 213914 133940 213920 133952
rect 175976 133912 213920 133940
rect 175976 133900 175982 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 275370 133900 275376 133952
rect 275428 133940 275434 133952
rect 307662 133940 307668 133952
rect 275428 133912 307668 133940
rect 275428 133900 275434 133912
rect 307662 133900 307668 133912
rect 307720 133900 307726 133952
rect 252278 133832 252284 133884
rect 252336 133872 252342 133884
rect 304442 133872 304448 133884
rect 252336 133844 304448 133872
rect 252336 133832 252342 133844
rect 304442 133832 304448 133844
rect 304500 133832 304506 133884
rect 324314 133832 324320 133884
rect 324372 133872 324378 133884
rect 346394 133872 346400 133884
rect 324372 133844 346400 133872
rect 324372 133832 324378 133844
rect 346394 133832 346400 133844
rect 346452 133832 346458 133884
rect 378778 133832 378784 133884
rect 378836 133872 378842 133884
rect 419350 133872 419356 133884
rect 378836 133844 419356 133872
rect 378836 133832 378842 133844
rect 419350 133832 419356 133844
rect 419408 133832 419414 133884
rect 252370 133764 252376 133816
rect 252428 133804 252434 133816
rect 286410 133804 286416 133816
rect 252428 133776 286416 133804
rect 252428 133764 252434 133776
rect 286410 133764 286416 133776
rect 286468 133764 286474 133816
rect 252462 133696 252468 133748
rect 252520 133736 252526 133748
rect 264238 133736 264244 133748
rect 252520 133708 264244 133736
rect 252520 133696 252526 133708
rect 264238 133696 264244 133708
rect 264296 133696 264302 133748
rect 258994 133152 259000 133204
rect 259052 133192 259058 133204
rect 307386 133192 307392 133204
rect 259052 133164 307392 133192
rect 259052 133152 259058 133164
rect 307386 133152 307392 133164
rect 307444 133152 307450 133204
rect 286502 132540 286508 132592
rect 286560 132580 286566 132592
rect 306926 132580 306932 132592
rect 286560 132552 306932 132580
rect 286560 132540 286566 132552
rect 306926 132540 306932 132552
rect 306984 132540 306990 132592
rect 187142 132472 187148 132524
rect 187200 132512 187206 132524
rect 213914 132512 213920 132524
rect 187200 132484 213920 132512
rect 187200 132472 187206 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 285122 132472 285128 132524
rect 285180 132512 285186 132524
rect 306558 132512 306564 132524
rect 285180 132484 306564 132512
rect 285180 132472 285186 132484
rect 306558 132472 306564 132484
rect 306616 132472 306622 132524
rect 324958 132472 324964 132524
rect 325016 132512 325022 132524
rect 327074 132512 327080 132524
rect 325016 132484 327080 132512
rect 325016 132472 325022 132484
rect 327074 132472 327080 132484
rect 327132 132472 327138 132524
rect 252370 132404 252376 132456
rect 252428 132444 252434 132456
rect 289262 132444 289268 132456
rect 252428 132416 289268 132444
rect 252428 132404 252434 132416
rect 289262 132404 289268 132416
rect 289320 132404 289326 132456
rect 324406 132404 324412 132456
rect 324464 132444 324470 132456
rect 357526 132444 357532 132456
rect 324464 132416 357532 132444
rect 324464 132404 324470 132416
rect 357526 132404 357532 132416
rect 357584 132404 357590 132456
rect 410518 132404 410524 132456
rect 410576 132444 410582 132456
rect 417602 132444 417608 132456
rect 410576 132416 417608 132444
rect 410576 132404 410582 132416
rect 417602 132404 417608 132416
rect 417660 132404 417666 132456
rect 252462 132336 252468 132388
rect 252520 132376 252526 132388
rect 273990 132376 273996 132388
rect 252520 132348 273996 132376
rect 252520 132336 252526 132348
rect 273990 132336 273996 132348
rect 274048 132336 274054 132388
rect 324314 132336 324320 132388
rect 324372 132376 324378 132388
rect 342346 132376 342352 132388
rect 324372 132348 342352 132376
rect 324372 132336 324378 132348
rect 342346 132336 342352 132348
rect 342404 132336 342410 132388
rect 294690 131248 294696 131300
rect 294748 131288 294754 131300
rect 307478 131288 307484 131300
rect 294748 131260 307484 131288
rect 294748 131248 294754 131260
rect 307478 131248 307484 131260
rect 307536 131248 307542 131300
rect 289078 131180 289084 131232
rect 289136 131220 289142 131232
rect 307570 131220 307576 131232
rect 289136 131192 307576 131220
rect 289136 131180 289142 131192
rect 307570 131180 307576 131192
rect 307628 131180 307634 131232
rect 173250 131112 173256 131164
rect 173308 131152 173314 131164
rect 213914 131152 213920 131164
rect 173308 131124 213920 131152
rect 173308 131112 173314 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 278130 131112 278136 131164
rect 278188 131152 278194 131164
rect 307662 131152 307668 131164
rect 278188 131124 307668 131152
rect 278188 131112 278194 131124
rect 307662 131112 307668 131124
rect 307720 131112 307726 131164
rect 252370 131044 252376 131096
rect 252428 131084 252434 131096
rect 290550 131084 290556 131096
rect 252428 131056 290556 131084
rect 252428 131044 252434 131056
rect 290550 131044 290556 131056
rect 290608 131044 290614 131096
rect 324314 131044 324320 131096
rect 324372 131084 324378 131096
rect 349154 131084 349160 131096
rect 324372 131056 349160 131084
rect 324372 131044 324378 131056
rect 349154 131044 349160 131056
rect 349212 131044 349218 131096
rect 252278 130976 252284 131028
rect 252336 131016 252342 131028
rect 267090 131016 267096 131028
rect 252336 130988 267096 131016
rect 252336 130976 252342 130988
rect 267090 130976 267096 130988
rect 267148 130976 267154 131028
rect 324406 130976 324412 131028
rect 324464 131016 324470 131028
rect 328730 131016 328736 131028
rect 324464 130988 328736 131016
rect 324464 130976 324470 130988
rect 328730 130976 328736 130988
rect 328788 130976 328794 131028
rect 252462 130908 252468 130960
rect 252520 130948 252526 130960
rect 262858 130948 262864 130960
rect 252520 130920 262864 130948
rect 252520 130908 252526 130920
rect 262858 130908 262864 130920
rect 262916 130908 262922 130960
rect 202230 130364 202236 130416
rect 202288 130404 202294 130416
rect 214742 130404 214748 130416
rect 202288 130376 214748 130404
rect 202288 130364 202294 130376
rect 214742 130364 214748 130376
rect 214800 130364 214806 130416
rect 267366 130364 267372 130416
rect 267424 130404 267430 130416
rect 305730 130404 305736 130416
rect 267424 130376 305736 130404
rect 267424 130364 267430 130376
rect 305730 130364 305736 130376
rect 305788 130364 305794 130416
rect 291930 129888 291936 129940
rect 291988 129928 291994 129940
rect 307662 129928 307668 129940
rect 291988 129900 307668 129928
rect 291988 129888 291994 129900
rect 307662 129888 307668 129900
rect 307720 129888 307726 129940
rect 290458 129820 290464 129872
rect 290516 129860 290522 129872
rect 307478 129860 307484 129872
rect 290516 129832 307484 129860
rect 290516 129820 290522 129832
rect 307478 129820 307484 129832
rect 307536 129820 307542 129872
rect 171870 129752 171876 129804
rect 171928 129792 171934 129804
rect 213914 129792 213920 129804
rect 171928 129764 213920 129792
rect 171928 129752 171934 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 273990 129752 273996 129804
rect 274048 129792 274054 129804
rect 307570 129792 307576 129804
rect 274048 129764 307576 129792
rect 274048 129752 274054 129764
rect 307570 129752 307576 129764
rect 307628 129752 307634 129804
rect 252462 129684 252468 129736
rect 252520 129724 252526 129736
rect 278222 129724 278228 129736
rect 252520 129696 278228 129724
rect 252520 129684 252526 129696
rect 278222 129684 278228 129696
rect 278280 129684 278286 129736
rect 324314 129684 324320 129736
rect 324372 129724 324378 129736
rect 352006 129724 352012 129736
rect 324372 129696 352012 129724
rect 324372 129684 324378 129696
rect 352006 129684 352012 129696
rect 352064 129684 352070 129736
rect 408402 129684 408408 129736
rect 408460 129724 408466 129736
rect 416774 129724 416780 129736
rect 408460 129696 416780 129724
rect 408460 129684 408466 129696
rect 416774 129684 416780 129696
rect 416832 129684 416838 129736
rect 496814 129684 496820 129736
rect 496872 129724 496878 129736
rect 510614 129724 510620 129736
rect 496872 129696 510620 129724
rect 496872 129684 496878 129696
rect 510614 129684 510620 129696
rect 510672 129684 510678 129736
rect 252370 129616 252376 129668
rect 252428 129656 252434 129668
rect 265802 129656 265808 129668
rect 252428 129628 265808 129656
rect 252428 129616 252434 129628
rect 265802 129616 265808 129628
rect 265860 129616 265866 129668
rect 324406 129616 324412 129668
rect 324464 129656 324470 129668
rect 331214 129656 331220 129668
rect 324464 129628 331220 129656
rect 324464 129616 324470 129628
rect 331214 129616 331220 129628
rect 331272 129616 331278 129668
rect 496906 129616 496912 129668
rect 496964 129656 496970 129668
rect 506658 129656 506664 129668
rect 496964 129628 506664 129656
rect 496964 129616 496970 129628
rect 506658 129616 506664 129628
rect 506716 129616 506722 129668
rect 252278 129548 252284 129600
rect 252336 129588 252342 129600
rect 257338 129588 257344 129600
rect 252336 129560 257344 129588
rect 252336 129548 252342 129560
rect 257338 129548 257344 129560
rect 257396 129548 257402 129600
rect 276750 128392 276756 128444
rect 276808 128432 276814 128444
rect 306926 128432 306932 128444
rect 276808 128404 306932 128432
rect 276808 128392 276814 128404
rect 306926 128392 306932 128404
rect 306984 128392 306990 128444
rect 188522 128324 188528 128376
rect 188580 128364 188586 128376
rect 213914 128364 213920 128376
rect 188580 128336 213920 128364
rect 188580 128324 188586 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 264238 128324 264244 128376
rect 264296 128364 264302 128376
rect 307662 128364 307668 128376
rect 264296 128336 307668 128364
rect 264296 128324 264302 128336
rect 307662 128324 307668 128336
rect 307720 128324 307726 128376
rect 252462 128256 252468 128308
rect 252520 128296 252526 128308
rect 287882 128296 287888 128308
rect 252520 128268 287888 128296
rect 252520 128256 252526 128268
rect 287882 128256 287888 128268
rect 287940 128256 287946 128308
rect 324314 128256 324320 128308
rect 324372 128296 324378 128308
rect 331306 128296 331312 128308
rect 324372 128268 331312 128296
rect 324372 128256 324378 128268
rect 331306 128256 331312 128268
rect 331364 128256 331370 128308
rect 377398 128256 377404 128308
rect 377456 128296 377462 128308
rect 419626 128296 419632 128308
rect 377456 128268 419632 128296
rect 377456 128256 377462 128268
rect 419626 128256 419632 128268
rect 419684 128296 419690 128308
rect 419810 128296 419816 128308
rect 419684 128268 419816 128296
rect 419684 128256 419690 128268
rect 419810 128256 419816 128268
rect 419868 128256 419874 128308
rect 252278 128188 252284 128240
rect 252336 128228 252342 128240
rect 269758 128228 269764 128240
rect 252336 128200 269764 128228
rect 252336 128188 252342 128200
rect 269758 128188 269764 128200
rect 269816 128188 269822 128240
rect 324406 128188 324412 128240
rect 324464 128228 324470 128240
rect 330110 128228 330116 128240
rect 324464 128200 330116 128228
rect 324464 128188 324470 128200
rect 330110 128188 330116 128200
rect 330168 128188 330174 128240
rect 252370 128120 252376 128172
rect 252428 128160 252434 128172
rect 258718 128160 258724 128172
rect 252428 128132 258724 128160
rect 252428 128120 252434 128132
rect 258718 128120 258724 128132
rect 258776 128120 258782 128172
rect 536098 127576 536104 127628
rect 536156 127616 536162 127628
rect 580166 127616 580172 127628
rect 536156 127588 580172 127616
rect 536156 127576 536162 127588
rect 580166 127576 580172 127588
rect 580224 127576 580230 127628
rect 287790 127100 287796 127152
rect 287848 127140 287854 127152
rect 307662 127140 307668 127152
rect 287848 127112 307668 127140
rect 287848 127100 287854 127112
rect 307662 127100 307668 127112
rect 307720 127100 307726 127152
rect 285030 127032 285036 127084
rect 285088 127072 285094 127084
rect 307478 127072 307484 127084
rect 285088 127044 307484 127072
rect 285088 127032 285094 127044
rect 307478 127032 307484 127044
rect 307536 127032 307542 127084
rect 59262 126964 59268 127016
rect 59320 127004 59326 127016
rect 65518 127004 65524 127016
rect 59320 126976 65524 127004
rect 59320 126964 59326 126976
rect 65518 126964 65524 126976
rect 65576 126964 65582 127016
rect 180150 126964 180156 127016
rect 180208 127004 180214 127016
rect 213914 127004 213920 127016
rect 180208 126976 213920 127004
rect 180208 126964 180214 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 269850 126964 269856 127016
rect 269908 127004 269914 127016
rect 307570 127004 307576 127016
rect 269908 126976 307576 127004
rect 269908 126964 269914 126976
rect 307570 126964 307576 126976
rect 307628 126964 307634 127016
rect 496906 126964 496912 127016
rect 496964 127004 496970 127016
rect 498286 127004 498292 127016
rect 496964 126976 498292 127004
rect 496964 126964 496970 126976
rect 498286 126964 498292 126976
rect 498344 126964 498350 127016
rect 252278 126896 252284 126948
rect 252336 126936 252342 126948
rect 283742 126936 283748 126948
rect 252336 126908 283748 126936
rect 252336 126896 252342 126908
rect 283742 126896 283748 126908
rect 283800 126896 283806 126948
rect 406378 126896 406384 126948
rect 406436 126936 406442 126948
rect 418522 126936 418528 126948
rect 406436 126908 418528 126936
rect 406436 126896 406442 126908
rect 418522 126896 418528 126908
rect 418580 126936 418586 126948
rect 419258 126936 419264 126948
rect 418580 126908 419264 126936
rect 418580 126896 418586 126908
rect 419258 126896 419264 126908
rect 419316 126896 419322 126948
rect 496814 126896 496820 126948
rect 496872 126936 496878 126948
rect 514754 126936 514760 126948
rect 496872 126908 514760 126936
rect 496872 126896 496878 126908
rect 514754 126896 514760 126908
rect 514812 126896 514818 126948
rect 252462 126828 252468 126880
rect 252520 126868 252526 126880
rect 268378 126868 268384 126880
rect 252520 126840 268384 126868
rect 252520 126828 252526 126840
rect 268378 126828 268384 126840
rect 268436 126828 268442 126880
rect 252370 126760 252376 126812
rect 252428 126800 252434 126812
rect 264422 126800 264428 126812
rect 252428 126772 264428 126800
rect 252428 126760 252434 126772
rect 264422 126760 264428 126772
rect 264480 126760 264486 126812
rect 202322 125672 202328 125724
rect 202380 125712 202386 125724
rect 213914 125712 213920 125724
rect 202380 125684 213920 125712
rect 202380 125672 202386 125684
rect 213914 125672 213920 125684
rect 213972 125672 213978 125724
rect 283650 125672 283656 125724
rect 283708 125712 283714 125724
rect 307570 125712 307576 125724
rect 283708 125684 307576 125712
rect 283708 125672 283714 125684
rect 307570 125672 307576 125684
rect 307628 125672 307634 125724
rect 169110 125604 169116 125656
rect 169168 125644 169174 125656
rect 214006 125644 214012 125656
rect 169168 125616 214012 125644
rect 169168 125604 169174 125616
rect 214006 125604 214012 125616
rect 214064 125604 214070 125656
rect 276934 125604 276940 125656
rect 276992 125644 276998 125656
rect 307662 125644 307668 125656
rect 276992 125616 307668 125644
rect 276992 125604 276998 125616
rect 307662 125604 307668 125616
rect 307720 125604 307726 125656
rect 252462 125536 252468 125588
rect 252520 125576 252526 125588
rect 297450 125576 297456 125588
rect 252520 125548 297456 125576
rect 252520 125536 252526 125548
rect 297450 125536 297456 125548
rect 297508 125536 297514 125588
rect 324314 125536 324320 125588
rect 324372 125576 324378 125588
rect 328546 125576 328552 125588
rect 324372 125548 328552 125576
rect 324372 125536 324378 125548
rect 328546 125536 328552 125548
rect 328604 125536 328610 125588
rect 342990 125536 342996 125588
rect 343048 125576 343054 125588
rect 418522 125576 418528 125588
rect 343048 125548 418528 125576
rect 343048 125536 343054 125548
rect 418522 125536 418528 125548
rect 418580 125576 418586 125588
rect 419442 125576 419448 125588
rect 418580 125548 419448 125576
rect 418580 125536 418586 125548
rect 419442 125536 419448 125548
rect 419500 125536 419506 125588
rect 496814 125536 496820 125588
rect 496872 125576 496878 125588
rect 521654 125576 521660 125588
rect 496872 125548 521660 125576
rect 496872 125536 496878 125548
rect 521654 125536 521660 125548
rect 521712 125536 521718 125588
rect 324406 125468 324412 125520
rect 324464 125508 324470 125520
rect 345106 125508 345112 125520
rect 324464 125480 345112 125508
rect 324464 125468 324470 125480
rect 345106 125468 345112 125480
rect 345164 125468 345170 125520
rect 252094 124924 252100 124976
rect 252152 124964 252158 124976
rect 263042 124964 263048 124976
rect 252152 124936 263048 124964
rect 252152 124924 252158 124936
rect 263042 124924 263048 124936
rect 263100 124924 263106 124976
rect 251818 124856 251824 124908
rect 251876 124896 251882 124908
rect 302970 124896 302976 124908
rect 251876 124868 302976 124896
rect 251876 124856 251882 124868
rect 302970 124856 302976 124868
rect 303028 124856 303034 124908
rect 303062 124380 303068 124432
rect 303120 124420 303126 124432
rect 307662 124420 307668 124432
rect 303120 124392 307668 124420
rect 303120 124380 303126 124392
rect 307662 124380 307668 124392
rect 307720 124380 307726 124432
rect 297542 124312 297548 124364
rect 297600 124352 297606 124364
rect 307570 124352 307576 124364
rect 297600 124324 307576 124352
rect 297600 124312 297606 124324
rect 307570 124312 307576 124324
rect 307628 124312 307634 124364
rect 199470 124244 199476 124296
rect 199528 124284 199534 124296
rect 213914 124284 213920 124296
rect 199528 124256 213920 124284
rect 199528 124244 199534 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 286410 124244 286416 124296
rect 286468 124284 286474 124296
rect 307478 124284 307484 124296
rect 286468 124256 307484 124284
rect 286468 124244 286474 124256
rect 307478 124244 307484 124256
rect 307536 124244 307542 124296
rect 170582 124176 170588 124228
rect 170640 124216 170646 124228
rect 214006 124216 214012 124228
rect 170640 124188 214012 124216
rect 170640 124176 170646 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 278222 124176 278228 124228
rect 278280 124216 278286 124228
rect 307662 124216 307668 124228
rect 278280 124188 307668 124216
rect 278280 124176 278286 124188
rect 307662 124176 307668 124188
rect 307720 124176 307726 124228
rect 252370 124108 252376 124160
rect 252428 124148 252434 124160
rect 304350 124148 304356 124160
rect 252428 124120 304356 124148
rect 252428 124108 252434 124120
rect 304350 124108 304356 124120
rect 304408 124108 304414 124160
rect 324314 124108 324320 124160
rect 324372 124148 324378 124160
rect 353294 124148 353300 124160
rect 324372 124120 353300 124148
rect 324372 124108 324378 124120
rect 353294 124108 353300 124120
rect 353352 124108 353358 124160
rect 496814 124108 496820 124160
rect 496872 124148 496878 124160
rect 499574 124148 499580 124160
rect 496872 124120 499580 124148
rect 496872 124108 496878 124120
rect 499574 124108 499580 124120
rect 499632 124108 499638 124160
rect 252462 124040 252468 124092
rect 252520 124080 252526 124092
rect 298922 124080 298928 124092
rect 252520 124052 298928 124080
rect 252520 124040 252526 124052
rect 298922 124040 298928 124052
rect 298980 124040 298986 124092
rect 252278 123972 252284 124024
rect 252336 124012 252342 124024
rect 261662 124012 261668 124024
rect 252336 123984 261668 124012
rect 252336 123972 252342 123984
rect 261662 123972 261668 123984
rect 261720 123972 261726 124024
rect 178954 122884 178960 122936
rect 179012 122924 179018 122936
rect 213914 122924 213920 122936
rect 179012 122896 213920 122924
rect 179012 122884 179018 122896
rect 213914 122884 213920 122896
rect 213972 122884 213978 122936
rect 298738 122884 298744 122936
rect 298796 122924 298802 122936
rect 307662 122924 307668 122936
rect 298796 122896 307668 122924
rect 298796 122884 298802 122896
rect 307662 122884 307668 122896
rect 307720 122884 307726 122936
rect 167822 122816 167828 122868
rect 167880 122856 167886 122868
rect 214006 122856 214012 122868
rect 167880 122828 214012 122856
rect 167880 122816 167886 122828
rect 214006 122816 214012 122828
rect 214064 122816 214070 122868
rect 297634 122816 297640 122868
rect 297692 122856 297698 122868
rect 307570 122856 307576 122868
rect 297692 122828 307576 122856
rect 297692 122816 297698 122828
rect 307570 122816 307576 122828
rect 307628 122816 307634 122868
rect 252462 122748 252468 122800
rect 252520 122788 252526 122800
rect 296070 122788 296076 122800
rect 252520 122760 296076 122788
rect 252520 122748 252526 122760
rect 296070 122748 296076 122760
rect 296128 122748 296134 122800
rect 324314 122748 324320 122800
rect 324372 122788 324378 122800
rect 342254 122788 342260 122800
rect 324372 122760 342260 122788
rect 324372 122748 324378 122760
rect 342254 122748 342260 122760
rect 342312 122748 342318 122800
rect 399478 122748 399484 122800
rect 399536 122788 399542 122800
rect 419534 122788 419540 122800
rect 399536 122760 419540 122788
rect 399536 122748 399542 122760
rect 419534 122748 419540 122760
rect 419592 122748 419598 122800
rect 252370 122680 252376 122732
rect 252428 122720 252434 122732
rect 272702 122720 272708 122732
rect 252428 122692 272708 122720
rect 252428 122680 252434 122692
rect 272702 122680 272708 122692
rect 272760 122680 272766 122732
rect 252278 122612 252284 122664
rect 252336 122652 252342 122664
rect 261478 122652 261484 122664
rect 252336 122624 261484 122652
rect 252336 122612 252342 122624
rect 261478 122612 261484 122624
rect 261536 122612 261542 122664
rect 170398 122068 170404 122120
rect 170456 122108 170462 122120
rect 196710 122108 196716 122120
rect 170456 122080 196716 122108
rect 170456 122068 170462 122080
rect 196710 122068 196716 122080
rect 196768 122068 196774 122120
rect 300394 121592 300400 121644
rect 300452 121632 300458 121644
rect 307570 121632 307576 121644
rect 300452 121604 307576 121632
rect 300452 121592 300458 121604
rect 307570 121592 307576 121604
rect 307628 121592 307634 121644
rect 198182 121524 198188 121576
rect 198240 121564 198246 121576
rect 214006 121564 214012 121576
rect 198240 121536 214012 121564
rect 198240 121524 198246 121536
rect 214006 121524 214012 121536
rect 214064 121524 214070 121576
rect 296254 121524 296260 121576
rect 296312 121564 296318 121576
rect 307662 121564 307668 121576
rect 296312 121536 307668 121564
rect 296312 121524 296318 121536
rect 307662 121524 307668 121536
rect 307720 121524 307726 121576
rect 180242 121456 180248 121508
rect 180300 121496 180306 121508
rect 213914 121496 213920 121508
rect 180300 121468 213920 121496
rect 180300 121456 180306 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 272610 121456 272616 121508
rect 272668 121496 272674 121508
rect 306742 121496 306748 121508
rect 272668 121468 306748 121496
rect 272668 121456 272674 121468
rect 306742 121456 306748 121468
rect 306800 121456 306806 121508
rect 252462 121388 252468 121440
rect 252520 121428 252526 121440
rect 256234 121428 256240 121440
rect 252520 121400 256240 121428
rect 252520 121388 252526 121400
rect 256234 121388 256240 121400
rect 256292 121388 256298 121440
rect 324314 121388 324320 121440
rect 324372 121428 324378 121440
rect 352098 121428 352104 121440
rect 324372 121400 352104 121428
rect 324372 121388 324378 121400
rect 352098 121388 352104 121400
rect 352156 121388 352162 121440
rect 496814 121388 496820 121440
rect 496872 121428 496878 121440
rect 517514 121428 517520 121440
rect 496872 121400 517520 121428
rect 496872 121388 496878 121400
rect 517514 121388 517520 121400
rect 517572 121388 517578 121440
rect 324406 121320 324412 121372
rect 324464 121360 324470 121372
rect 347774 121360 347780 121372
rect 324464 121332 347780 121360
rect 324464 121320 324470 121332
rect 347774 121320 347780 121332
rect 347832 121320 347838 121372
rect 258718 120232 258724 120284
rect 258776 120272 258782 120284
rect 307294 120272 307300 120284
rect 258776 120244 307300 120272
rect 258776 120232 258782 120244
rect 307294 120232 307300 120244
rect 307352 120232 307358 120284
rect 210510 120164 210516 120216
rect 210568 120204 210574 120216
rect 214006 120204 214012 120216
rect 210568 120176 214012 120204
rect 210568 120164 210574 120176
rect 214006 120164 214012 120176
rect 214064 120164 214070 120216
rect 250530 120164 250536 120216
rect 250588 120204 250594 120216
rect 250588 120176 254992 120204
rect 250588 120164 250594 120176
rect 176102 120096 176108 120148
rect 176160 120136 176166 120148
rect 213914 120136 213920 120148
rect 176160 120108 213920 120136
rect 176160 120096 176166 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 252002 120096 252008 120148
rect 252060 120136 252066 120148
rect 254854 120136 254860 120148
rect 252060 120108 254860 120136
rect 252060 120096 252066 120108
rect 254854 120096 254860 120108
rect 254912 120096 254918 120148
rect 254964 120136 254992 120176
rect 257338 120164 257344 120216
rect 257396 120204 257402 120216
rect 307662 120204 307668 120216
rect 257396 120176 307668 120204
rect 257396 120164 257402 120176
rect 307662 120164 307668 120176
rect 307720 120164 307726 120216
rect 307570 120136 307576 120148
rect 254964 120108 307576 120136
rect 307570 120096 307576 120108
rect 307628 120096 307634 120148
rect 252278 120028 252284 120080
rect 252336 120068 252342 120080
rect 292022 120068 292028 120080
rect 252336 120040 292028 120068
rect 252336 120028 252342 120040
rect 292022 120028 292028 120040
rect 292080 120028 292086 120080
rect 400858 120028 400864 120080
rect 400916 120068 400922 120080
rect 416774 120068 416780 120080
rect 400916 120040 416780 120068
rect 400916 120028 400922 120040
rect 416774 120028 416780 120040
rect 416832 120028 416838 120080
rect 252462 119960 252468 120012
rect 252520 120000 252526 120012
rect 265710 120000 265716 120012
rect 252520 119972 265716 120000
rect 252520 119960 252526 119972
rect 265710 119960 265716 119972
rect 265768 119960 265774 120012
rect 252370 119824 252376 119876
rect 252428 119864 252434 119876
rect 260190 119864 260196 119876
rect 252428 119836 260196 119864
rect 252428 119824 252434 119836
rect 260190 119824 260196 119836
rect 260248 119824 260254 119876
rect 496814 119756 496820 119808
rect 496872 119796 496878 119808
rect 499758 119796 499764 119808
rect 496872 119768 499764 119796
rect 496872 119756 496878 119768
rect 499758 119756 499764 119768
rect 499816 119756 499822 119808
rect 271506 119348 271512 119400
rect 271564 119388 271570 119400
rect 307202 119388 307208 119400
rect 271564 119360 307208 119388
rect 271564 119348 271570 119360
rect 307202 119348 307208 119360
rect 307260 119348 307266 119400
rect 193950 118804 193956 118856
rect 194008 118844 194014 118856
rect 214006 118844 214012 118856
rect 194008 118816 214012 118844
rect 194008 118804 194014 118816
rect 214006 118804 214012 118816
rect 214064 118804 214070 118856
rect 279602 118804 279608 118856
rect 279660 118844 279666 118856
rect 306558 118844 306564 118856
rect 279660 118816 306564 118844
rect 279660 118804 279666 118816
rect 306558 118804 306564 118816
rect 306616 118804 306622 118856
rect 185670 118736 185676 118788
rect 185728 118776 185734 118788
rect 213914 118776 213920 118788
rect 185728 118748 213920 118776
rect 185728 118736 185734 118748
rect 213914 118736 213920 118748
rect 213972 118736 213978 118788
rect 299014 118736 299020 118788
rect 299072 118776 299078 118788
rect 307662 118776 307668 118788
rect 299072 118748 307668 118776
rect 299072 118736 299078 118748
rect 307662 118736 307668 118748
rect 307720 118736 307726 118788
rect 177482 118668 177488 118720
rect 177540 118708 177546 118720
rect 214098 118708 214104 118720
rect 177540 118680 214104 118708
rect 177540 118668 177546 118680
rect 214098 118668 214104 118680
rect 214156 118668 214162 118720
rect 252370 118600 252376 118652
rect 252428 118640 252434 118652
rect 300210 118640 300216 118652
rect 252428 118612 300216 118640
rect 252428 118600 252434 118612
rect 300210 118600 300216 118612
rect 300268 118600 300274 118652
rect 324314 118600 324320 118652
rect 324372 118640 324378 118652
rect 354674 118640 354680 118652
rect 324372 118612 354680 118640
rect 324372 118600 324378 118612
rect 354674 118600 354680 118612
rect 354732 118600 354738 118652
rect 414658 118600 414664 118652
rect 414716 118640 414722 118652
rect 416958 118640 416964 118652
rect 414716 118612 416964 118640
rect 414716 118600 414722 118612
rect 416958 118600 416964 118612
rect 417016 118600 417022 118652
rect 496814 118600 496820 118652
rect 496872 118640 496878 118652
rect 512178 118640 512184 118652
rect 496872 118612 512184 118640
rect 496872 118600 496878 118612
rect 512178 118600 512184 118612
rect 512236 118600 512242 118652
rect 252278 118532 252284 118584
rect 252336 118572 252342 118584
rect 274082 118572 274088 118584
rect 252336 118544 274088 118572
rect 252336 118532 252342 118544
rect 274082 118532 274088 118544
rect 274140 118532 274146 118584
rect 324406 118532 324412 118584
rect 324464 118572 324470 118584
rect 347866 118572 347872 118584
rect 324464 118544 347872 118572
rect 324464 118532 324470 118544
rect 347866 118532 347872 118544
rect 347924 118532 347930 118584
rect 496906 118532 496912 118584
rect 496964 118572 496970 118584
rect 509234 118572 509240 118584
rect 496964 118544 509240 118572
rect 496964 118532 496970 118544
rect 509234 118532 509240 118544
rect 509292 118532 509298 118584
rect 252462 117648 252468 117700
rect 252520 117688 252526 117700
rect 258810 117688 258816 117700
rect 252520 117660 258816 117688
rect 252520 117648 252526 117660
rect 258810 117648 258816 117660
rect 258868 117648 258874 117700
rect 265710 117512 265716 117564
rect 265768 117552 265774 117564
rect 307662 117552 307668 117564
rect 265768 117524 307668 117552
rect 265768 117512 265774 117524
rect 307662 117512 307668 117524
rect 307720 117512 307726 117564
rect 196894 117376 196900 117428
rect 196952 117416 196958 117428
rect 214006 117416 214012 117428
rect 196952 117388 214012 117416
rect 196952 117376 196958 117388
rect 214006 117376 214012 117388
rect 214064 117376 214070 117428
rect 283742 117376 283748 117428
rect 283800 117416 283806 117428
rect 307570 117416 307576 117428
rect 283800 117388 307576 117416
rect 283800 117376 283806 117388
rect 307570 117376 307576 117388
rect 307628 117376 307634 117428
rect 170398 117308 170404 117360
rect 170456 117348 170462 117360
rect 213914 117348 213920 117360
rect 170456 117320 213920 117348
rect 170456 117308 170462 117320
rect 213914 117308 213920 117320
rect 213972 117308 213978 117360
rect 304350 117308 304356 117360
rect 304408 117348 304414 117360
rect 307294 117348 307300 117360
rect 304408 117320 307300 117348
rect 304408 117308 304414 117320
rect 307294 117308 307300 117320
rect 307352 117308 307358 117360
rect 252462 117240 252468 117292
rect 252520 117280 252526 117292
rect 271230 117280 271236 117292
rect 252520 117252 271236 117280
rect 252520 117240 252526 117252
rect 271230 117240 271236 117252
rect 271288 117240 271294 117292
rect 324314 117240 324320 117292
rect 324372 117280 324378 117292
rect 340966 117280 340972 117292
rect 324372 117252 340972 117280
rect 324372 117240 324378 117252
rect 340966 117240 340972 117252
rect 341024 117240 341030 117292
rect 252370 117172 252376 117224
rect 252428 117212 252434 117224
rect 261570 117212 261576 117224
rect 252428 117184 261576 117212
rect 252428 117172 252434 117184
rect 261570 117172 261576 117184
rect 261628 117172 261634 117224
rect 251910 116560 251916 116612
rect 251968 116600 251974 116612
rect 267274 116600 267280 116612
rect 251968 116572 267280 116600
rect 251968 116560 251974 116572
rect 267274 116560 267280 116572
rect 267332 116560 267338 116612
rect 293310 116084 293316 116136
rect 293368 116124 293374 116136
rect 307662 116124 307668 116136
rect 293368 116096 307668 116124
rect 293368 116084 293374 116096
rect 307662 116084 307668 116096
rect 307720 116084 307726 116136
rect 174814 116016 174820 116068
rect 174872 116056 174878 116068
rect 214006 116056 214012 116068
rect 174872 116028 214012 116056
rect 174872 116016 174878 116028
rect 214006 116016 214012 116028
rect 214064 116016 214070 116068
rect 271138 116016 271144 116068
rect 271196 116056 271202 116068
rect 307570 116056 307576 116068
rect 271196 116028 307576 116056
rect 271196 116016 271202 116028
rect 307570 116016 307576 116028
rect 307628 116016 307634 116068
rect 169202 115948 169208 116000
rect 169260 115988 169266 116000
rect 213914 115988 213920 116000
rect 169260 115960 213920 115988
rect 169260 115948 169266 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 266998 115948 267004 116000
rect 267056 115988 267062 116000
rect 307478 115988 307484 116000
rect 267056 115960 307484 115988
rect 267056 115948 267062 115960
rect 307478 115948 307484 115960
rect 307536 115948 307542 116000
rect 252462 115880 252468 115932
rect 252520 115920 252526 115932
rect 285214 115920 285220 115932
rect 252520 115892 285220 115920
rect 252520 115880 252526 115892
rect 285214 115880 285220 115892
rect 285272 115880 285278 115932
rect 324314 115880 324320 115932
rect 324372 115920 324378 115932
rect 350626 115920 350632 115932
rect 324372 115892 350632 115920
rect 324372 115880 324378 115892
rect 350626 115880 350632 115892
rect 350684 115880 350690 115932
rect 496814 115880 496820 115932
rect 496872 115920 496878 115932
rect 503714 115920 503720 115932
rect 496872 115892 503720 115920
rect 496872 115880 496878 115892
rect 503714 115880 503720 115892
rect 503772 115880 503778 115932
rect 252370 115812 252376 115864
rect 252428 115852 252434 115864
rect 264330 115852 264336 115864
rect 252428 115824 264336 115852
rect 252428 115812 252434 115824
rect 264330 115812 264336 115824
rect 264388 115812 264394 115864
rect 324406 115812 324412 115864
rect 324464 115852 324470 115864
rect 343634 115852 343640 115864
rect 324464 115824 343640 115852
rect 324464 115812 324470 115824
rect 343634 115812 343640 115824
rect 343692 115812 343698 115864
rect 252278 115200 252284 115252
rect 252336 115240 252342 115252
rect 268470 115240 268476 115252
rect 252336 115212 268476 115240
rect 252336 115200 252342 115212
rect 268470 115200 268476 115212
rect 268528 115200 268534 115252
rect 296070 114656 296076 114708
rect 296128 114696 296134 114708
rect 307570 114696 307576 114708
rect 296128 114668 307576 114696
rect 296128 114656 296134 114668
rect 307570 114656 307576 114668
rect 307628 114656 307634 114708
rect 211890 114588 211896 114640
rect 211948 114628 211954 114640
rect 214006 114628 214012 114640
rect 211948 114600 214012 114628
rect 211948 114588 211954 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 280982 114588 280988 114640
rect 281040 114628 281046 114640
rect 307662 114628 307668 114640
rect 281040 114600 307668 114628
rect 281040 114588 281046 114600
rect 307662 114588 307668 114600
rect 307720 114588 307726 114640
rect 167730 114520 167736 114572
rect 167788 114560 167794 114572
rect 213914 114560 213920 114572
rect 167788 114532 213920 114560
rect 167788 114520 167794 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 268378 114520 268384 114572
rect 268436 114560 268442 114572
rect 307294 114560 307300 114572
rect 268436 114532 307300 114560
rect 268436 114520 268442 114532
rect 307294 114520 307300 114532
rect 307352 114520 307358 114572
rect 252462 114452 252468 114504
rect 252520 114492 252526 114504
rect 286594 114492 286600 114504
rect 252520 114464 286600 114492
rect 252520 114452 252526 114464
rect 286594 114452 286600 114464
rect 286652 114452 286658 114504
rect 333330 114452 333336 114504
rect 333388 114492 333394 114504
rect 416774 114492 416780 114504
rect 333388 114464 416780 114492
rect 333388 114452 333394 114464
rect 416774 114452 416780 114464
rect 416832 114452 416838 114504
rect 496814 114452 496820 114504
rect 496872 114492 496878 114504
rect 499666 114492 499672 114504
rect 496872 114464 499672 114492
rect 496872 114452 496878 114464
rect 499666 114452 499672 114464
rect 499724 114452 499730 114504
rect 324314 114384 324320 114436
rect 324372 114424 324378 114436
rect 349338 114424 349344 114436
rect 324372 114396 349344 114424
rect 324372 114384 324378 114396
rect 349338 114384 349344 114396
rect 349396 114384 349402 114436
rect 252370 113772 252376 113824
rect 252428 113812 252434 113824
rect 301590 113812 301596 113824
rect 252428 113784 301596 113812
rect 252428 113772 252434 113784
rect 301590 113772 301596 113784
rect 301648 113772 301654 113824
rect 195422 113228 195428 113280
rect 195480 113268 195486 113280
rect 214006 113268 214012 113280
rect 195480 113240 214012 113268
rect 195480 113228 195486 113240
rect 214006 113228 214012 113240
rect 214064 113228 214070 113280
rect 301682 113228 301688 113280
rect 301740 113268 301746 113280
rect 306558 113268 306564 113280
rect 301740 113240 306564 113268
rect 301740 113228 301746 113240
rect 306558 113228 306564 113240
rect 306616 113228 306622 113280
rect 167914 113160 167920 113212
rect 167972 113200 167978 113212
rect 213914 113200 213920 113212
rect 167972 113172 213920 113200
rect 167972 113160 167978 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 290550 113160 290556 113212
rect 290608 113200 290614 113212
rect 307662 113200 307668 113212
rect 290608 113172 307668 113200
rect 290608 113160 290614 113172
rect 307662 113160 307668 113172
rect 307720 113160 307726 113212
rect 252462 113092 252468 113144
rect 252520 113132 252526 113144
rect 299106 113132 299112 113144
rect 252520 113104 299112 113132
rect 252520 113092 252526 113104
rect 299106 113092 299112 113104
rect 299164 113092 299170 113144
rect 324314 113092 324320 113144
rect 324372 113132 324378 113144
rect 338114 113132 338120 113144
rect 324372 113104 338120 113132
rect 324372 113092 324378 113104
rect 338114 113092 338120 113104
rect 338172 113092 338178 113144
rect 496814 113092 496820 113144
rect 496872 113132 496878 113144
rect 501046 113132 501052 113144
rect 496872 113104 501052 113132
rect 496872 113092 496878 113104
rect 501046 113092 501052 113104
rect 501104 113092 501110 113144
rect 252278 113024 252284 113076
rect 252336 113064 252342 113076
rect 256142 113064 256148 113076
rect 252336 113036 256148 113064
rect 252336 113024 252342 113036
rect 256142 113024 256148 113036
rect 256200 113024 256206 113076
rect 337470 113024 337476 113076
rect 337528 113064 337534 113076
rect 416774 113064 416780 113076
rect 337528 113036 416780 113064
rect 337528 113024 337534 113036
rect 416774 113024 416780 113036
rect 416832 113024 416838 113076
rect 252278 112412 252284 112464
rect 252336 112452 252342 112464
rect 276842 112452 276848 112464
rect 252336 112424 276848 112452
rect 252336 112412 252342 112424
rect 276842 112412 276848 112424
rect 276900 112412 276906 112464
rect 298922 111936 298928 111988
rect 298980 111976 298986 111988
rect 307662 111976 307668 111988
rect 298980 111948 307668 111976
rect 298980 111936 298986 111948
rect 307662 111936 307668 111948
rect 307720 111936 307726 111988
rect 297450 111868 297456 111920
rect 297508 111908 297514 111920
rect 307570 111908 307576 111920
rect 297508 111880 307576 111908
rect 297508 111868 297514 111880
rect 307570 111868 307576 111880
rect 307628 111868 307634 111920
rect 166350 111800 166356 111852
rect 166408 111840 166414 111852
rect 213914 111840 213920 111852
rect 166408 111812 213920 111840
rect 166408 111800 166414 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 269758 111800 269764 111852
rect 269816 111840 269822 111852
rect 307478 111840 307484 111852
rect 269816 111812 307484 111840
rect 269816 111800 269822 111812
rect 307478 111800 307484 111812
rect 307536 111800 307542 111852
rect 168006 111732 168012 111784
rect 168064 111772 168070 111784
rect 176010 111772 176016 111784
rect 168064 111744 176016 111772
rect 168064 111732 168070 111744
rect 176010 111732 176016 111744
rect 176068 111732 176074 111784
rect 251174 111732 251180 111784
rect 251232 111772 251238 111784
rect 253382 111772 253388 111784
rect 251232 111744 253388 111772
rect 251232 111732 251238 111744
rect 253382 111732 253388 111744
rect 253440 111732 253446 111784
rect 367738 111732 367744 111784
rect 367796 111772 367802 111784
rect 416774 111772 416780 111784
rect 367796 111744 416780 111772
rect 367796 111732 367802 111744
rect 416774 111732 416780 111744
rect 416832 111732 416838 111784
rect 496906 111732 496912 111784
rect 496964 111772 496970 111784
rect 503806 111772 503812 111784
rect 496964 111744 503812 111772
rect 496964 111732 496970 111744
rect 503806 111732 503812 111744
rect 503864 111732 503870 111784
rect 252370 111664 252376 111716
rect 252428 111704 252434 111716
rect 257430 111704 257436 111716
rect 252428 111676 257436 111704
rect 252428 111664 252434 111676
rect 257430 111664 257436 111676
rect 257488 111664 257494 111716
rect 496814 111664 496820 111716
rect 496872 111704 496878 111716
rect 502426 111704 502432 111716
rect 496872 111676 502432 111704
rect 496872 111664 496878 111676
rect 502426 111664 502432 111676
rect 502484 111664 502490 111716
rect 252462 111596 252468 111648
rect 252520 111636 252526 111648
rect 281074 111636 281080 111648
rect 252520 111608 281080 111636
rect 252520 111596 252526 111608
rect 281074 111596 281080 111608
rect 281132 111596 281138 111648
rect 3694 111052 3700 111104
rect 3752 111092 3758 111104
rect 4062 111092 4068 111104
rect 3752 111064 4068 111092
rect 3752 111052 3758 111064
rect 4062 111052 4068 111064
rect 4120 111092 4126 111104
rect 14458 111092 14464 111104
rect 4120 111064 14464 111092
rect 4120 111052 4126 111064
rect 14458 111052 14464 111064
rect 14516 111052 14522 111104
rect 294782 110576 294788 110628
rect 294840 110616 294846 110628
rect 306742 110616 306748 110628
rect 294840 110588 306748 110616
rect 294840 110576 294846 110588
rect 306742 110576 306748 110588
rect 306800 110576 306806 110628
rect 184474 110508 184480 110560
rect 184532 110548 184538 110560
rect 213914 110548 213920 110560
rect 184532 110520 213920 110548
rect 184532 110508 184538 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 292022 110508 292028 110560
rect 292080 110548 292086 110560
rect 307294 110548 307300 110560
rect 292080 110520 307300 110548
rect 292080 110508 292086 110520
rect 307294 110508 307300 110520
rect 307352 110508 307358 110560
rect 169294 110440 169300 110492
rect 169352 110480 169358 110492
rect 214006 110480 214012 110492
rect 169352 110452 214012 110480
rect 169352 110440 169358 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 279510 110440 279516 110492
rect 279568 110480 279574 110492
rect 307662 110480 307668 110492
rect 279568 110452 307668 110480
rect 279568 110440 279574 110452
rect 307662 110440 307668 110452
rect 307720 110440 307726 110492
rect 168098 110372 168104 110424
rect 168156 110412 168162 110424
rect 213362 110412 213368 110424
rect 168156 110384 213368 110412
rect 168156 110372 168162 110384
rect 213362 110372 213368 110384
rect 213420 110372 213426 110424
rect 251726 110372 251732 110424
rect 251784 110412 251790 110424
rect 254670 110412 254676 110424
rect 251784 110384 254676 110412
rect 251784 110372 251790 110384
rect 254670 110372 254676 110384
rect 254728 110372 254734 110424
rect 324314 110372 324320 110424
rect 324372 110412 324378 110424
rect 341058 110412 341064 110424
rect 324372 110384 341064 110412
rect 324372 110372 324378 110384
rect 341058 110372 341064 110384
rect 341116 110372 341122 110424
rect 496814 110372 496820 110424
rect 496872 110412 496878 110424
rect 506566 110412 506572 110424
rect 496872 110384 506572 110412
rect 496872 110372 496878 110384
rect 506566 110372 506572 110384
rect 506624 110372 506630 110424
rect 252462 110304 252468 110356
rect 252520 110344 252526 110356
rect 255958 110344 255964 110356
rect 252520 110316 255964 110344
rect 252520 110304 252526 110316
rect 255958 110304 255964 110316
rect 256016 110304 256022 110356
rect 302878 109148 302884 109200
rect 302936 109188 302942 109200
rect 307570 109188 307576 109200
rect 302936 109160 307576 109188
rect 302936 109148 302942 109160
rect 307570 109148 307576 109160
rect 307628 109148 307634 109200
rect 257430 109080 257436 109132
rect 257488 109120 257494 109132
rect 306926 109120 306932 109132
rect 257488 109092 306932 109120
rect 257488 109080 257494 109092
rect 306926 109080 306932 109092
rect 306984 109080 306990 109132
rect 172054 109012 172060 109064
rect 172112 109052 172118 109064
rect 213914 109052 213920 109064
rect 172112 109024 213920 109052
rect 172112 109012 172118 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 253198 109012 253204 109064
rect 253256 109052 253262 109064
rect 307662 109052 307668 109064
rect 253256 109024 307668 109052
rect 253256 109012 253262 109024
rect 307662 109012 307668 109024
rect 307720 109012 307726 109064
rect 252370 108944 252376 108996
rect 252428 108984 252434 108996
rect 278314 108984 278320 108996
rect 252428 108956 278320 108984
rect 252428 108944 252434 108956
rect 278314 108944 278320 108956
rect 278372 108944 278378 108996
rect 324314 108944 324320 108996
rect 324372 108984 324378 108996
rect 345198 108984 345204 108996
rect 324372 108956 345204 108984
rect 324372 108944 324378 108956
rect 345198 108944 345204 108956
rect 345256 108944 345262 108996
rect 252462 108876 252468 108928
rect 252520 108916 252526 108928
rect 275554 108916 275560 108928
rect 252520 108888 275560 108916
rect 252520 108876 252526 108888
rect 275554 108876 275560 108888
rect 275612 108876 275618 108928
rect 268470 107856 268476 107908
rect 268528 107896 268534 107908
rect 307478 107896 307484 107908
rect 268528 107868 307484 107896
rect 268528 107856 268534 107868
rect 307478 107856 307484 107868
rect 307536 107856 307542 107908
rect 174722 107720 174728 107772
rect 174780 107760 174786 107772
rect 214006 107760 214012 107772
rect 174780 107732 214012 107760
rect 174780 107720 174786 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 275462 107720 275468 107772
rect 275520 107760 275526 107772
rect 307662 107760 307668 107772
rect 275520 107732 307668 107760
rect 275520 107720 275526 107732
rect 307662 107720 307668 107732
rect 307720 107720 307726 107772
rect 170674 107652 170680 107704
rect 170732 107692 170738 107704
rect 213914 107692 213920 107704
rect 170732 107664 213920 107692
rect 170732 107652 170738 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 300302 107652 300308 107704
rect 300360 107692 300366 107704
rect 307570 107692 307576 107704
rect 300360 107664 307576 107692
rect 300360 107652 300366 107664
rect 307570 107652 307576 107664
rect 307628 107652 307634 107704
rect 252462 107584 252468 107636
rect 252520 107624 252526 107636
rect 267182 107624 267188 107636
rect 252520 107596 267188 107624
rect 252520 107584 252526 107596
rect 267182 107584 267188 107596
rect 267240 107584 267246 107636
rect 413278 107584 413284 107636
rect 413336 107624 413342 107636
rect 416774 107624 416780 107636
rect 413336 107596 416780 107624
rect 413336 107584 413342 107596
rect 416774 107584 416780 107596
rect 416832 107584 416838 107636
rect 252370 107516 252376 107568
rect 252428 107556 252434 107568
rect 256050 107556 256056 107568
rect 252428 107528 256056 107556
rect 252428 107516 252434 107528
rect 256050 107516 256056 107528
rect 256108 107516 256114 107568
rect 252462 106904 252468 106956
rect 252520 106944 252526 106956
rect 258994 106944 259000 106956
rect 252520 106916 259000 106944
rect 252520 106904 252526 106916
rect 258994 106904 259000 106916
rect 259052 106904 259058 106956
rect 301590 106428 301596 106480
rect 301648 106468 301654 106480
rect 307662 106468 307668 106480
rect 301648 106440 307668 106468
rect 301648 106428 301654 106440
rect 307662 106428 307668 106440
rect 307720 106428 307726 106480
rect 176010 106360 176016 106412
rect 176068 106400 176074 106412
rect 213914 106400 213920 106412
rect 176068 106372 213920 106400
rect 176068 106360 176074 106372
rect 213914 106360 213920 106372
rect 213972 106360 213978 106412
rect 264330 106360 264336 106412
rect 264388 106400 264394 106412
rect 307478 106400 307484 106412
rect 264388 106372 307484 106400
rect 264388 106360 264394 106372
rect 307478 106360 307484 106372
rect 307536 106360 307542 106412
rect 167638 106292 167644 106344
rect 167696 106332 167702 106344
rect 214006 106332 214012 106344
rect 167696 106304 214012 106332
rect 167696 106292 167702 106304
rect 214006 106292 214012 106304
rect 214064 106292 214070 106344
rect 256142 106292 256148 106344
rect 256200 106332 256206 106344
rect 306742 106332 306748 106344
rect 256200 106304 306748 106332
rect 256200 106292 256206 106304
rect 306742 106292 306748 106304
rect 306800 106292 306806 106344
rect 371878 106224 371884 106276
rect 371936 106264 371942 106276
rect 416774 106264 416780 106276
rect 371936 106236 416780 106264
rect 371936 106224 371942 106236
rect 416774 106224 416780 106236
rect 416832 106224 416838 106276
rect 324314 105816 324320 105868
rect 324372 105856 324378 105868
rect 327166 105856 327172 105868
rect 324372 105828 327172 105856
rect 324372 105816 324378 105828
rect 327166 105816 327172 105828
rect 327224 105816 327230 105868
rect 251358 105612 251364 105664
rect 251416 105652 251422 105664
rect 262950 105652 262956 105664
rect 251416 105624 262956 105652
rect 251416 105612 251422 105624
rect 262950 105612 262956 105624
rect 263008 105612 263014 105664
rect 252370 105544 252376 105596
rect 252428 105584 252434 105596
rect 292114 105584 292120 105596
rect 252428 105556 292120 105584
rect 252428 105544 252434 105556
rect 292114 105544 292120 105556
rect 292172 105544 292178 105596
rect 203610 105000 203616 105052
rect 203668 105040 203674 105052
rect 213914 105040 213920 105052
rect 203668 105012 213920 105040
rect 203668 105000 203674 105012
rect 213914 105000 213920 105012
rect 213972 105000 213978 105052
rect 303154 105000 303160 105052
rect 303212 105040 303218 105052
rect 307570 105040 307576 105052
rect 303212 105012 307576 105040
rect 303212 105000 303218 105012
rect 307570 105000 307576 105012
rect 307628 105000 307634 105052
rect 188614 104932 188620 104984
rect 188672 104972 188678 104984
rect 214006 104972 214012 104984
rect 188672 104944 214012 104972
rect 188672 104932 188678 104944
rect 214006 104932 214012 104944
rect 214064 104932 214070 104984
rect 282362 104932 282368 104984
rect 282420 104972 282426 104984
rect 307662 104972 307668 104984
rect 282420 104944 307668 104972
rect 282420 104932 282426 104944
rect 307662 104932 307668 104944
rect 307720 104932 307726 104984
rect 173434 104864 173440 104916
rect 173492 104904 173498 104916
rect 214098 104904 214104 104916
rect 173492 104876 214104 104904
rect 173492 104864 173498 104876
rect 214098 104864 214104 104876
rect 214156 104864 214162 104916
rect 261478 104864 261484 104916
rect 261536 104904 261542 104916
rect 306742 104904 306748 104916
rect 261536 104876 306748 104904
rect 261536 104864 261542 104876
rect 306742 104864 306748 104876
rect 306800 104864 306806 104916
rect 252462 104796 252468 104848
rect 252520 104836 252526 104848
rect 271506 104836 271512 104848
rect 252520 104808 271512 104836
rect 252520 104796 252526 104808
rect 271506 104796 271512 104808
rect 271564 104796 271570 104848
rect 395338 104796 395344 104848
rect 395396 104836 395402 104848
rect 416774 104836 416780 104848
rect 395396 104808 416780 104836
rect 395396 104796 395402 104808
rect 416774 104796 416780 104808
rect 416832 104796 416838 104848
rect 252278 104728 252284 104780
rect 252336 104768 252342 104780
rect 257522 104768 257528 104780
rect 252336 104740 257528 104768
rect 252336 104728 252342 104740
rect 257522 104728 257528 104740
rect 257580 104728 257586 104780
rect 330478 104116 330484 104168
rect 330536 104156 330542 104168
rect 403618 104156 403624 104168
rect 330536 104128 403624 104156
rect 330536 104116 330542 104128
rect 403618 104116 403624 104128
rect 403676 104116 403682 104168
rect 286594 103640 286600 103692
rect 286652 103680 286658 103692
rect 307478 103680 307484 103692
rect 286652 103652 307484 103680
rect 286652 103640 286658 103652
rect 307478 103640 307484 103652
rect 307536 103640 307542 103692
rect 271322 103572 271328 103624
rect 271380 103612 271386 103624
rect 306926 103612 306932 103624
rect 271380 103584 306932 103612
rect 271380 103572 271386 103584
rect 306926 103572 306932 103584
rect 306984 103572 306990 103624
rect 206554 103504 206560 103556
rect 206612 103544 206618 103556
rect 213914 103544 213920 103556
rect 206612 103516 213920 103544
rect 206612 103504 206618 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 255958 103504 255964 103556
rect 256016 103544 256022 103556
rect 306742 103544 306748 103556
rect 256016 103516 306748 103544
rect 256016 103504 256022 103516
rect 306742 103504 306748 103516
rect 306800 103504 306806 103556
rect 252370 103436 252376 103488
rect 252428 103476 252434 103488
rect 274174 103476 274180 103488
rect 252428 103448 274180 103476
rect 252428 103436 252434 103448
rect 274174 103436 274180 103448
rect 274232 103436 274238 103488
rect 354030 103436 354036 103488
rect 354088 103476 354094 103488
rect 416774 103476 416780 103488
rect 354088 103448 416780 103476
rect 354088 103436 354094 103448
rect 416774 103436 416780 103448
rect 416832 103436 416838 103488
rect 251726 102824 251732 102876
rect 251784 102864 251790 102876
rect 254762 102864 254768 102876
rect 251784 102836 254768 102864
rect 251784 102824 251790 102836
rect 254762 102824 254768 102836
rect 254820 102824 254826 102876
rect 495434 102824 495440 102876
rect 495492 102864 495498 102876
rect 495618 102864 495624 102876
rect 495492 102836 495624 102864
rect 495492 102824 495498 102836
rect 495618 102824 495624 102836
rect 495676 102824 495682 102876
rect 173342 102756 173348 102808
rect 173400 102796 173406 102808
rect 214650 102796 214656 102808
rect 173400 102768 214656 102796
rect 173400 102756 173406 102768
rect 214650 102756 214656 102768
rect 214708 102756 214714 102808
rect 252462 102552 252468 102604
rect 252520 102592 252526 102604
rect 258902 102592 258908 102604
rect 252520 102564 258908 102592
rect 252520 102552 252526 102564
rect 258902 102552 258908 102564
rect 258960 102552 258966 102604
rect 289262 102280 289268 102332
rect 289320 102320 289326 102332
rect 306558 102320 306564 102332
rect 289320 102292 306564 102320
rect 289320 102280 289326 102292
rect 306558 102280 306564 102292
rect 306616 102280 306622 102332
rect 274082 102212 274088 102264
rect 274140 102252 274146 102264
rect 307662 102252 307668 102264
rect 274140 102224 307668 102252
rect 274140 102212 274146 102224
rect 307662 102212 307668 102224
rect 307720 102212 307726 102264
rect 209222 102144 209228 102196
rect 209280 102184 209286 102196
rect 213914 102184 213920 102196
rect 209280 102156 213920 102184
rect 209280 102144 209286 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 258810 102144 258816 102196
rect 258868 102184 258874 102196
rect 307570 102184 307576 102196
rect 258868 102156 307576 102184
rect 258868 102144 258874 102156
rect 307570 102144 307576 102156
rect 307628 102144 307634 102196
rect 252462 102076 252468 102128
rect 252520 102116 252526 102128
rect 290642 102116 290648 102128
rect 252520 102088 290648 102116
rect 252520 102076 252526 102088
rect 290642 102076 290648 102088
rect 290700 102076 290706 102128
rect 382918 102076 382924 102128
rect 382976 102116 382982 102128
rect 416774 102116 416780 102128
rect 382976 102088 416780 102116
rect 382976 102076 382982 102088
rect 416774 102076 416780 102088
rect 416832 102076 416838 102128
rect 252370 102008 252376 102060
rect 252428 102048 252434 102060
rect 287974 102048 287980 102060
rect 252428 102020 287980 102048
rect 252428 102008 252434 102020
rect 287974 102008 287980 102020
rect 288032 102008 288038 102060
rect 252186 101396 252192 101448
rect 252244 101436 252250 101448
rect 271414 101436 271420 101448
rect 252244 101408 271420 101436
rect 252244 101396 252250 101408
rect 271414 101396 271420 101408
rect 271472 101396 271478 101448
rect 326338 101396 326344 101448
rect 326396 101436 326402 101448
rect 376018 101436 376024 101448
rect 326396 101408 376024 101436
rect 326396 101396 326402 101408
rect 376018 101396 376024 101408
rect 376076 101396 376082 101448
rect 511258 101396 511264 101448
rect 511316 101436 511322 101448
rect 580166 101436 580172 101448
rect 511316 101408 580172 101436
rect 511316 101396 511322 101408
rect 580166 101396 580172 101408
rect 580224 101396 580230 101448
rect 271230 100920 271236 100972
rect 271288 100960 271294 100972
rect 307662 100960 307668 100972
rect 271288 100932 307668 100960
rect 271288 100920 271294 100932
rect 307662 100920 307668 100932
rect 307720 100920 307726 100972
rect 300210 100852 300216 100904
rect 300268 100892 300274 100904
rect 306558 100892 306564 100904
rect 300268 100864 306564 100892
rect 300268 100852 300274 100864
rect 306558 100852 306564 100864
rect 306616 100852 306622 100904
rect 287882 100784 287888 100836
rect 287940 100824 287946 100836
rect 307570 100824 307576 100836
rect 287940 100796 307576 100824
rect 287940 100784 287946 100796
rect 307570 100784 307576 100796
rect 307628 100784 307634 100836
rect 177574 100716 177580 100768
rect 177632 100756 177638 100768
rect 213914 100756 213920 100768
rect 177632 100728 213920 100756
rect 177632 100716 177638 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 304442 100716 304448 100768
rect 304500 100756 304506 100768
rect 307478 100756 307484 100768
rect 304500 100728 307484 100756
rect 304500 100716 304506 100728
rect 307478 100716 307484 100728
rect 307536 100716 307542 100768
rect 252278 100648 252284 100700
rect 252336 100688 252342 100700
rect 301866 100688 301872 100700
rect 252336 100660 301872 100688
rect 252336 100648 252342 100660
rect 301866 100648 301872 100660
rect 301924 100648 301930 100700
rect 419718 100648 419724 100700
rect 419776 100688 419782 100700
rect 580258 100688 580264 100700
rect 419776 100660 580264 100688
rect 419776 100648 419782 100660
rect 580258 100648 580264 100660
rect 580316 100648 580322 100700
rect 252462 100580 252468 100632
rect 252520 100620 252526 100632
rect 289354 100620 289360 100632
rect 252520 100592 289360 100620
rect 252520 100580 252526 100592
rect 289354 100580 289360 100592
rect 289412 100580 289418 100632
rect 389818 100580 389824 100632
rect 389876 100620 389882 100632
rect 496814 100620 496820 100632
rect 389876 100592 496820 100620
rect 389876 100580 389882 100592
rect 496814 100580 496820 100592
rect 496872 100580 496878 100632
rect 252370 100512 252376 100564
rect 252428 100552 252434 100564
rect 268562 100552 268568 100564
rect 252428 100524 268568 100552
rect 252428 100512 252434 100524
rect 268562 100512 268568 100524
rect 268620 100512 268626 100564
rect 323578 99968 323584 100020
rect 323636 100008 323642 100020
rect 411898 100008 411904 100020
rect 323636 99980 411904 100008
rect 323636 99968 323642 99980
rect 411898 99968 411904 99980
rect 411956 99968 411962 100020
rect 301774 99492 301780 99544
rect 301832 99532 301838 99544
rect 307478 99532 307484 99544
rect 301832 99504 307484 99532
rect 301832 99492 301838 99504
rect 307478 99492 307484 99504
rect 307536 99492 307542 99544
rect 296162 99424 296168 99476
rect 296220 99464 296226 99476
rect 307570 99464 307576 99476
rect 296220 99436 307576 99464
rect 296220 99424 296226 99436
rect 307570 99424 307576 99436
rect 307628 99424 307634 99476
rect 211982 99356 211988 99408
rect 212040 99396 212046 99408
rect 214282 99396 214288 99408
rect 212040 99368 214288 99396
rect 212040 99356 212046 99368
rect 214282 99356 214288 99368
rect 214340 99356 214346 99408
rect 285214 99356 285220 99408
rect 285272 99396 285278 99408
rect 307662 99396 307668 99408
rect 285272 99368 307668 99396
rect 285272 99356 285278 99368
rect 307662 99356 307668 99368
rect 307720 99356 307726 99408
rect 252370 99288 252376 99340
rect 252428 99328 252434 99340
rect 303246 99328 303252 99340
rect 252428 99300 303252 99328
rect 252428 99288 252434 99300
rect 303246 99288 303252 99300
rect 303304 99288 303310 99340
rect 388438 99288 388444 99340
rect 388496 99328 388502 99340
rect 497090 99328 497096 99340
rect 388496 99300 497096 99328
rect 388496 99288 388502 99300
rect 497090 99288 497096 99300
rect 497148 99288 497154 99340
rect 252462 99220 252468 99272
rect 252520 99260 252526 99272
rect 267366 99260 267372 99272
rect 252520 99232 267372 99260
rect 252520 99220 252526 99232
rect 267366 99220 267372 99232
rect 267424 99220 267430 99272
rect 393958 99220 393964 99272
rect 394016 99260 394022 99272
rect 496998 99260 497004 99272
rect 394016 99232 497004 99260
rect 394016 99220 394022 99232
rect 496998 99220 497004 99232
rect 497056 99220 497062 99272
rect 396718 99152 396724 99204
rect 396776 99192 396782 99204
rect 494054 99192 494060 99204
rect 396776 99164 494060 99192
rect 396776 99152 396782 99164
rect 494054 99152 494060 99164
rect 494112 99152 494118 99204
rect 302970 98132 302976 98184
rect 303028 98172 303034 98184
rect 307662 98172 307668 98184
rect 303028 98144 307668 98172
rect 303028 98132 303034 98144
rect 307662 98132 307668 98144
rect 307720 98132 307726 98184
rect 199562 98064 199568 98116
rect 199620 98104 199626 98116
rect 213914 98104 213920 98116
rect 199620 98076 213920 98104
rect 199620 98064 199626 98076
rect 213914 98064 213920 98076
rect 213972 98064 213978 98116
rect 281074 98064 281080 98116
rect 281132 98104 281138 98116
rect 307570 98104 307576 98116
rect 281132 98076 307576 98104
rect 281132 98064 281138 98076
rect 307570 98064 307576 98076
rect 307628 98064 307634 98116
rect 166442 97996 166448 98048
rect 166500 98036 166506 98048
rect 214006 98036 214012 98048
rect 166500 98008 214012 98036
rect 166500 97996 166506 98008
rect 214006 97996 214012 98008
rect 214064 97996 214070 98048
rect 249242 97996 249248 98048
rect 249300 98036 249306 98048
rect 307294 98036 307300 98048
rect 249300 98008 307300 98036
rect 249300 97996 249306 98008
rect 307294 97996 307300 98008
rect 307352 97996 307358 98048
rect 370498 97928 370504 97980
rect 370556 97968 370562 97980
rect 495434 97968 495440 97980
rect 370556 97940 495440 97968
rect 370556 97928 370562 97940
rect 495434 97928 495440 97940
rect 495492 97928 495498 97980
rect 392578 97860 392584 97912
rect 392636 97900 392642 97912
rect 496906 97900 496912 97912
rect 392636 97872 496912 97900
rect 392636 97860 392642 97872
rect 496906 97860 496912 97872
rect 496964 97860 496970 97912
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 421006 97316 421012 97368
rect 421064 97356 421070 97368
rect 426526 97356 426532 97368
rect 421064 97328 426532 97356
rect 421064 97316 421070 97328
rect 426526 97316 426532 97328
rect 426584 97316 426590 97368
rect 421558 97248 421564 97300
rect 421616 97288 421622 97300
rect 456518 97288 456524 97300
rect 421616 97260 456524 97288
rect 421616 97248 421622 97260
rect 456518 97248 456524 97260
rect 456576 97248 456582 97300
rect 461578 97248 461584 97300
rect 461636 97288 461642 97300
rect 474550 97288 474556 97300
rect 461636 97260 474556 97288
rect 461636 97248 461642 97260
rect 474550 97248 474556 97260
rect 474608 97248 474614 97300
rect 475378 97248 475384 97300
rect 475436 97288 475442 97300
rect 492490 97288 492496 97300
rect 475436 97260 492496 97288
rect 475436 97248 475442 97260
rect 492490 97248 492496 97260
rect 492548 97248 492554 97300
rect 414658 96908 414664 96960
rect 414716 96948 414722 96960
rect 420546 96948 420552 96960
rect 414716 96920 420552 96948
rect 414716 96908 414722 96920
rect 420546 96908 420552 96920
rect 420604 96908 420610 96960
rect 439498 96908 439504 96960
rect 439556 96948 439562 96960
rect 440878 96948 440884 96960
rect 439556 96920 440884 96948
rect 439556 96908 439562 96920
rect 440878 96908 440884 96920
rect 440936 96908 440942 96960
rect 454034 96908 454040 96960
rect 454092 96948 454098 96960
rect 455046 96948 455052 96960
rect 454092 96920 455052 96948
rect 454092 96908 454098 96920
rect 455046 96908 455052 96920
rect 455104 96908 455110 96960
rect 481634 96908 481640 96960
rect 481692 96948 481698 96960
rect 482646 96948 482652 96960
rect 481692 96920 482652 96948
rect 481692 96908 481698 96920
rect 482646 96908 482652 96920
rect 482704 96908 482710 96960
rect 486418 96908 486424 96960
rect 486476 96948 486482 96960
rect 487706 96948 487712 96960
rect 486476 96920 487712 96948
rect 486476 96908 486482 96920
rect 487706 96908 487712 96920
rect 487764 96908 487770 96960
rect 457438 96772 457444 96824
rect 457496 96812 457502 96824
rect 460106 96812 460112 96824
rect 457496 96784 460112 96812
rect 457496 96772 457502 96784
rect 460106 96772 460112 96784
rect 460164 96772 460170 96824
rect 278314 96704 278320 96756
rect 278372 96744 278378 96756
rect 307662 96744 307668 96756
rect 278372 96716 307668 96744
rect 278372 96704 278378 96716
rect 307662 96704 307668 96716
rect 307720 96704 307726 96756
rect 267090 96636 267096 96688
rect 267148 96676 267154 96688
rect 307570 96676 307576 96688
rect 267148 96648 307576 96676
rect 267148 96636 267154 96648
rect 307570 96636 307576 96648
rect 307628 96636 307634 96688
rect 191190 96568 191196 96620
rect 191248 96608 191254 96620
rect 323026 96608 323032 96620
rect 191248 96580 323032 96608
rect 191248 96568 191254 96580
rect 323026 96568 323032 96580
rect 323084 96568 323090 96620
rect 381538 96568 381544 96620
rect 381596 96608 381602 96620
rect 495618 96608 495624 96620
rect 381596 96580 495624 96608
rect 381596 96568 381602 96580
rect 495618 96568 495624 96580
rect 495676 96568 495682 96620
rect 300118 96500 300124 96552
rect 300176 96540 300182 96552
rect 321462 96540 321468 96552
rect 300176 96512 321468 96540
rect 300176 96500 300182 96512
rect 321462 96500 321468 96512
rect 321520 96500 321526 96552
rect 351914 96500 351920 96552
rect 351972 96540 351978 96552
rect 421006 96540 421012 96552
rect 351972 96512 421012 96540
rect 351972 96500 351978 96512
rect 421006 96500 421012 96512
rect 421064 96500 421070 96552
rect 166902 95888 166908 95940
rect 166960 95928 166966 95940
rect 214098 95928 214104 95940
rect 166960 95900 214104 95928
rect 166960 95888 166966 95900
rect 214098 95888 214104 95900
rect 214156 95888 214162 95940
rect 324314 95888 324320 95940
rect 324372 95928 324378 95940
rect 351914 95928 351920 95940
rect 324372 95900 351920 95928
rect 324372 95888 324378 95900
rect 351914 95888 351920 95900
rect 351972 95888 351978 95940
rect 419166 95888 419172 95940
rect 419224 95928 419230 95940
rect 580258 95928 580264 95940
rect 419224 95900 580264 95928
rect 419224 95888 419230 95900
rect 580258 95888 580264 95900
rect 580316 95888 580322 95940
rect 164878 95616 164884 95668
rect 164936 95656 164942 95668
rect 165614 95656 165620 95668
rect 164936 95628 165620 95656
rect 164936 95616 164942 95628
rect 165614 95616 165620 95628
rect 165672 95616 165678 95668
rect 251818 95208 251824 95260
rect 251876 95248 251882 95260
rect 307662 95248 307668 95260
rect 251876 95220 307668 95248
rect 251876 95208 251882 95220
rect 307662 95208 307668 95220
rect 307720 95208 307726 95260
rect 178770 95140 178776 95192
rect 178828 95180 178834 95192
rect 321554 95180 321560 95192
rect 178828 95152 321560 95180
rect 178828 95140 178834 95152
rect 321554 95140 321560 95152
rect 321612 95140 321618 95192
rect 337378 95140 337384 95192
rect 337436 95180 337442 95192
rect 498470 95180 498476 95192
rect 337436 95152 498476 95180
rect 337436 95140 337442 95152
rect 498470 95140 498476 95152
rect 498528 95140 498534 95192
rect 181438 95072 181444 95124
rect 181496 95112 181502 95124
rect 321370 95112 321376 95124
rect 181496 95084 321376 95112
rect 181496 95072 181502 95084
rect 321370 95072 321376 95084
rect 321428 95072 321434 95124
rect 193858 95004 193864 95056
rect 193916 95044 193922 95056
rect 322934 95044 322940 95056
rect 193916 95016 322940 95044
rect 193916 95004 193922 95016
rect 322934 95004 322940 95016
rect 322992 95004 322998 95056
rect 199378 94936 199384 94988
rect 199436 94976 199442 94988
rect 321646 94976 321652 94988
rect 199436 94948 321652 94976
rect 199436 94936 199442 94948
rect 321646 94936 321652 94948
rect 321704 94936 321710 94988
rect 206370 94868 206376 94920
rect 206428 94908 206434 94920
rect 321830 94908 321836 94920
rect 206428 94880 321836 94908
rect 206428 94868 206434 94880
rect 321830 94868 321836 94880
rect 321888 94868 321894 94920
rect 336734 94664 336740 94716
rect 336792 94704 336798 94716
rect 337378 94704 337384 94716
rect 336792 94676 337384 94704
rect 336792 94664 336798 94676
rect 337378 94664 337384 94676
rect 337436 94664 337442 94716
rect 320818 94460 320824 94512
rect 320876 94500 320882 94512
rect 427722 94500 427728 94512
rect 320876 94472 427728 94500
rect 320876 94460 320882 94472
rect 427722 94460 427728 94472
rect 427780 94460 427786 94512
rect 152090 94120 152096 94172
rect 152148 94160 152154 94172
rect 189718 94160 189724 94172
rect 152148 94132 189724 94160
rect 152148 94120 152154 94132
rect 189718 94120 189724 94132
rect 189776 94120 189782 94172
rect 126514 94052 126520 94104
rect 126572 94092 126578 94104
rect 169110 94092 169116 94104
rect 126572 94064 169116 94092
rect 126572 94052 126578 94064
rect 169110 94052 169116 94064
rect 169168 94052 169174 94104
rect 126698 93984 126704 94036
rect 126756 94024 126762 94036
rect 181530 94024 181536 94036
rect 126756 93996 181536 94024
rect 126756 93984 126762 93996
rect 181530 93984 181536 93996
rect 181588 93984 181594 94036
rect 112346 93916 112352 93968
rect 112404 93956 112410 93968
rect 185670 93956 185676 93968
rect 112404 93928 185676 93956
rect 112404 93916 112410 93928
rect 185670 93916 185676 93928
rect 185728 93916 185734 93968
rect 96154 93848 96160 93900
rect 96212 93888 96218 93900
rect 172054 93888 172060 93900
rect 96212 93860 172060 93888
rect 96212 93848 96218 93860
rect 172054 93848 172060 93860
rect 172112 93848 172118 93900
rect 133138 93440 133144 93492
rect 133196 93480 133202 93492
rect 171778 93480 171784 93492
rect 133196 93452 171784 93480
rect 133196 93440 133202 93452
rect 171778 93440 171784 93452
rect 171836 93440 171842 93492
rect 151722 93372 151728 93424
rect 151780 93412 151786 93424
rect 191282 93412 191288 93424
rect 151780 93384 191288 93412
rect 151780 93372 151786 93384
rect 191282 93372 191288 93384
rect 191340 93372 191346 93424
rect 121730 93304 121736 93356
rect 121788 93344 121794 93356
rect 167822 93344 167828 93356
rect 121788 93316 167828 93344
rect 121788 93304 121794 93316
rect 167822 93304 167828 93316
rect 167880 93304 167886 93356
rect 116762 93236 116768 93288
rect 116820 93276 116826 93288
rect 166258 93276 166264 93288
rect 116820 93248 166264 93276
rect 116820 93236 116826 93248
rect 166258 93236 166264 93248
rect 166316 93236 166322 93288
rect 109218 93168 109224 93220
rect 109276 93208 109282 93220
rect 174814 93208 174820 93220
rect 109276 93180 174820 93208
rect 109276 93168 109282 93180
rect 174814 93168 174820 93180
rect 174872 93168 174878 93220
rect 100938 93100 100944 93152
rect 100996 93140 101002 93152
rect 188522 93140 188528 93152
rect 100996 93112 188528 93140
rect 100996 93100 101002 93112
rect 188522 93100 188528 93112
rect 188580 93100 188586 93152
rect 232498 93100 232504 93152
rect 232556 93140 232562 93152
rect 278222 93140 278228 93152
rect 232556 93112 278228 93140
rect 232556 93100 232562 93112
rect 278222 93100 278228 93112
rect 278280 93100 278286 93152
rect 88978 92420 88984 92472
rect 89036 92460 89042 92472
rect 166902 92460 166908 92472
rect 89036 92432 166908 92460
rect 89036 92420 89042 92432
rect 166902 92420 166908 92432
rect 166960 92420 166966 92472
rect 187050 92420 187056 92472
rect 187108 92460 187114 92472
rect 321738 92460 321744 92472
rect 187108 92432 321744 92460
rect 187108 92420 187114 92432
rect 321738 92420 321744 92432
rect 321796 92420 321802 92472
rect 118050 92352 118056 92404
rect 118108 92392 118114 92404
rect 195330 92392 195336 92404
rect 118108 92364 195336 92392
rect 118108 92352 118114 92364
rect 195330 92352 195336 92364
rect 195388 92352 195394 92404
rect 196802 92352 196808 92404
rect 196860 92392 196866 92404
rect 321922 92392 321928 92404
rect 196860 92364 321928 92392
rect 196860 92352 196866 92364
rect 321922 92352 321928 92364
rect 321980 92352 321986 92404
rect 115474 92284 115480 92336
rect 115532 92324 115538 92336
rect 210418 92324 210424 92336
rect 115532 92296 210424 92324
rect 115532 92284 115538 92296
rect 210418 92284 210424 92296
rect 210476 92284 210482 92336
rect 114462 92216 114468 92268
rect 114520 92256 114526 92268
rect 202230 92256 202236 92268
rect 114520 92228 202236 92256
rect 114520 92216 114526 92228
rect 202230 92216 202236 92228
rect 202288 92216 202294 92268
rect 103330 92148 103336 92200
rect 103388 92188 103394 92200
rect 173342 92188 173348 92200
rect 103388 92160 173348 92188
rect 103388 92148 103394 92160
rect 173342 92148 173348 92160
rect 173400 92148 173406 92200
rect 132402 92080 132408 92132
rect 132460 92120 132466 92132
rect 177390 92120 177396 92132
rect 132460 92092 177396 92120
rect 132460 92080 132466 92092
rect 177390 92080 177396 92092
rect 177448 92080 177454 92132
rect 238018 91808 238024 91860
rect 238076 91848 238082 91860
rect 251174 91848 251180 91860
rect 238076 91820 251180 91848
rect 238076 91808 238082 91820
rect 251174 91808 251180 91820
rect 251232 91808 251238 91860
rect 200758 91740 200764 91792
rect 200816 91780 200822 91792
rect 253382 91780 253388 91792
rect 200816 91752 253388 91780
rect 200816 91740 200822 91752
rect 253382 91740 253388 91752
rect 253440 91740 253446 91792
rect 277394 91740 277400 91792
rect 277452 91780 277458 91792
rect 481726 91780 481732 91792
rect 277452 91752 481732 91780
rect 277452 91740 277458 91752
rect 481726 91740 481732 91752
rect 481784 91740 481790 91792
rect 74810 91128 74816 91180
rect 74868 91168 74874 91180
rect 88978 91168 88984 91180
rect 74868 91140 88984 91168
rect 74868 91128 74874 91140
rect 88978 91128 88984 91140
rect 89036 91128 89042 91180
rect 97534 91128 97540 91180
rect 97592 91168 97598 91180
rect 116118 91168 116124 91180
rect 97592 91140 116124 91168
rect 97592 91128 97598 91140
rect 116118 91128 116124 91140
rect 116176 91128 116182 91180
rect 85850 91060 85856 91112
rect 85908 91100 85914 91112
rect 122098 91100 122104 91112
rect 85908 91072 122104 91100
rect 85908 91060 85914 91072
rect 122098 91060 122104 91072
rect 122156 91060 122162 91112
rect 88058 90992 88064 91044
rect 88116 91032 88122 91044
rect 211982 91032 211988 91044
rect 88116 91004 211988 91032
rect 88116 90992 88122 91004
rect 211982 90992 211988 91004
rect 212040 90992 212046 91044
rect 252462 90992 252468 91044
rect 252520 91032 252526 91044
rect 420914 91032 420920 91044
rect 252520 91004 420920 91032
rect 252520 90992 252526 91004
rect 420914 90992 420920 91004
rect 420972 90992 420978 91044
rect 98822 90924 98828 90976
rect 98880 90964 98886 90976
rect 184474 90964 184480 90976
rect 98880 90936 184480 90964
rect 98880 90924 98886 90936
rect 184474 90924 184480 90936
rect 184532 90924 184538 90976
rect 114922 90856 114928 90908
rect 114980 90896 114986 90908
rect 193950 90896 193956 90908
rect 114980 90868 193956 90896
rect 114980 90856 114986 90868
rect 193950 90856 193956 90868
rect 194008 90856 194014 90908
rect 103238 90788 103244 90840
rect 103296 90828 103302 90840
rect 167914 90828 167920 90840
rect 103296 90800 167920 90828
rect 103296 90788 103302 90800
rect 167914 90788 167920 90800
rect 167972 90788 167978 90840
rect 151538 90720 151544 90772
rect 151596 90760 151602 90772
rect 178862 90760 178868 90772
rect 151596 90732 178868 90760
rect 151596 90720 151602 90732
rect 178862 90720 178868 90732
rect 178920 90720 178926 90772
rect 151630 90652 151636 90704
rect 151688 90692 151694 90704
rect 173158 90692 173164 90704
rect 151688 90664 173164 90692
rect 151688 90652 151694 90664
rect 173158 90652 173164 90664
rect 173216 90652 173222 90704
rect 311894 90380 311900 90432
rect 311952 90420 311958 90432
rect 358078 90420 358084 90432
rect 311952 90392 358084 90420
rect 311952 90380 311958 90392
rect 358078 90380 358084 90392
rect 358136 90380 358142 90432
rect 352650 90312 352656 90364
rect 352708 90352 352714 90364
rect 456794 90352 456800 90364
rect 352708 90324 456800 90352
rect 352708 90312 352714 90324
rect 456794 90312 456800 90324
rect 456852 90312 456858 90364
rect 251910 89700 251916 89752
rect 251968 89740 251974 89752
rect 252462 89740 252468 89752
rect 251968 89712 252468 89740
rect 251968 89700 251974 89712
rect 252462 89700 252468 89712
rect 252520 89700 252526 89752
rect 67634 89632 67640 89684
rect 67692 89672 67698 89684
rect 214834 89672 214840 89684
rect 67692 89644 214840 89672
rect 67692 89632 67698 89644
rect 214834 89632 214840 89644
rect 214892 89632 214898 89684
rect 348418 89632 348424 89684
rect 348476 89672 348482 89684
rect 501138 89672 501144 89684
rect 348476 89644 501144 89672
rect 348476 89632 348482 89644
rect 501138 89632 501144 89644
rect 501196 89632 501202 89684
rect 110138 89564 110144 89616
rect 110196 89604 110202 89616
rect 170398 89604 170404 89616
rect 110196 89576 170404 89604
rect 110196 89564 110202 89576
rect 170398 89564 170404 89576
rect 170456 89564 170462 89616
rect 182818 89564 182824 89616
rect 182876 89604 182882 89616
rect 324406 89604 324412 89616
rect 182876 89576 324412 89604
rect 182876 89564 182882 89576
rect 324406 89564 324412 89576
rect 324464 89564 324470 89616
rect 90726 89496 90732 89548
rect 90784 89536 90790 89548
rect 188614 89536 188620 89548
rect 90784 89508 188620 89536
rect 90784 89496 90790 89508
rect 188614 89496 188620 89508
rect 188672 89496 188678 89548
rect 122834 89428 122840 89480
rect 122892 89468 122898 89480
rect 199470 89468 199476 89480
rect 122892 89440 199476 89468
rect 122892 89428 122898 89440
rect 199470 89428 199476 89440
rect 199528 89428 199534 89480
rect 119798 89360 119804 89412
rect 119856 89400 119862 89412
rect 174630 89400 174636 89412
rect 119856 89372 174636 89400
rect 119856 89360 119862 89372
rect 174630 89360 174636 89372
rect 174688 89360 174694 89412
rect 136450 89292 136456 89344
rect 136508 89332 136514 89344
rect 182910 89332 182916 89344
rect 136508 89304 182916 89332
rect 136508 89292 136514 89304
rect 182910 89292 182916 89304
rect 182968 89292 182974 89344
rect 347774 89224 347780 89276
rect 347832 89264 347838 89276
rect 348418 89264 348424 89276
rect 347832 89236 348424 89264
rect 347832 89224 347838 89236
rect 348418 89224 348424 89236
rect 348476 89224 348482 89276
rect 295978 88952 295984 89004
rect 296036 88992 296042 89004
rect 315298 88992 315304 89004
rect 296036 88964 315304 88992
rect 296036 88952 296042 88964
rect 315298 88952 315304 88964
rect 315356 88952 315362 89004
rect 316678 88952 316684 89004
rect 316736 88992 316742 89004
rect 345658 88992 345664 89004
rect 316736 88964 345664 88992
rect 316736 88952 316742 88964
rect 345658 88952 345664 88964
rect 345716 88952 345722 89004
rect 67726 88272 67732 88324
rect 67784 88312 67790 88324
rect 214650 88312 214656 88324
rect 67784 88284 214656 88312
rect 67784 88272 67790 88284
rect 214650 88272 214656 88284
rect 214708 88272 214714 88324
rect 116118 88204 116124 88256
rect 116176 88244 116182 88256
rect 214742 88244 214748 88256
rect 116176 88216 214748 88244
rect 116176 88204 116182 88216
rect 214742 88204 214748 88216
rect 214800 88204 214806 88256
rect 104250 88136 104256 88188
rect 104308 88176 104314 88188
rect 195422 88176 195428 88188
rect 104308 88148 195428 88176
rect 104308 88136 104314 88148
rect 195422 88136 195428 88148
rect 195480 88136 195486 88188
rect 120718 88068 120724 88120
rect 120776 88108 120782 88120
rect 178954 88108 178960 88120
rect 120776 88080 178960 88108
rect 120776 88068 120782 88080
rect 178954 88068 178960 88080
rect 179012 88068 179018 88120
rect 129458 88000 129464 88052
rect 129516 88040 129522 88052
rect 169018 88040 169024 88052
rect 129516 88012 169024 88040
rect 129516 88000 129522 88012
rect 169018 88000 169024 88012
rect 169076 88000 169082 88052
rect 308490 87660 308496 87712
rect 308548 87700 308554 87712
rect 324958 87700 324964 87712
rect 308548 87672 324964 87700
rect 308548 87660 308554 87672
rect 324958 87660 324964 87672
rect 325016 87660 325022 87712
rect 213178 87592 213184 87644
rect 213236 87632 213242 87644
rect 276014 87632 276020 87644
rect 213236 87604 276020 87632
rect 213236 87592 213242 87604
rect 276014 87592 276020 87604
rect 276072 87592 276078 87644
rect 278038 87592 278044 87644
rect 278096 87632 278102 87644
rect 331950 87632 331956 87644
rect 278096 87604 331956 87632
rect 278096 87592 278102 87604
rect 331950 87592 331956 87604
rect 332008 87592 332014 87644
rect 342346 87592 342352 87644
rect 342404 87632 342410 87644
rect 458174 87632 458180 87644
rect 342404 87604 458180 87632
rect 342404 87592 342410 87604
rect 458174 87592 458180 87604
rect 458232 87592 458238 87644
rect 276014 86980 276020 87032
rect 276072 87020 276078 87032
rect 276842 87020 276848 87032
rect 276072 86992 276848 87020
rect 276072 86980 276078 86992
rect 276842 86980 276848 86992
rect 276900 87020 276906 87032
rect 277394 87020 277400 87032
rect 276900 86992 277400 87020
rect 276900 86980 276906 86992
rect 277394 86980 277400 86992
rect 277452 86980 277458 87032
rect 88978 86912 88984 86964
rect 89036 86952 89042 86964
rect 214558 86952 214564 86964
rect 89036 86924 214564 86952
rect 89036 86912 89042 86924
rect 214558 86912 214564 86924
rect 214616 86912 214622 86964
rect 339494 86912 339500 86964
rect 339552 86952 339558 86964
rect 340138 86952 340144 86964
rect 339552 86924 340144 86952
rect 339552 86912 339558 86924
rect 340138 86912 340144 86924
rect 340196 86952 340202 86964
rect 457438 86952 457444 86964
rect 340196 86924 457444 86952
rect 340196 86912 340202 86924
rect 457438 86912 457444 86924
rect 457496 86912 457502 86964
rect 504450 86912 504456 86964
rect 504508 86952 504514 86964
rect 580166 86952 580172 86964
rect 504508 86924 580172 86952
rect 504508 86912 504514 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 126514 86844 126520 86896
rect 126572 86884 126578 86896
rect 213270 86884 213276 86896
rect 126572 86856 213276 86884
rect 126572 86844 126578 86856
rect 213270 86844 213276 86856
rect 213328 86844 213334 86896
rect 86770 86776 86776 86828
rect 86828 86816 86834 86828
rect 166442 86816 166448 86828
rect 86828 86788 166448 86816
rect 86828 86776 86834 86788
rect 166442 86776 166448 86788
rect 166500 86776 166506 86828
rect 100570 86708 100576 86760
rect 100628 86748 100634 86760
rect 166350 86748 166356 86760
rect 100628 86720 166356 86748
rect 100628 86708 100634 86720
rect 166350 86708 166356 86720
rect 166408 86708 166414 86760
rect 107930 86640 107936 86692
rect 107988 86680 107994 86692
rect 169202 86680 169208 86692
rect 107988 86652 169208 86680
rect 107988 86640 107994 86652
rect 169202 86640 169208 86652
rect 169260 86640 169266 86692
rect 117130 86572 117136 86624
rect 117188 86612 117194 86624
rect 176102 86612 176108 86624
rect 117188 86584 176108 86612
rect 117188 86572 117194 86584
rect 176102 86572 176108 86584
rect 176160 86572 176166 86624
rect 211798 86232 211804 86284
rect 211856 86272 211862 86284
rect 322198 86272 322204 86284
rect 211856 86244 322204 86272
rect 211856 86232 211862 86244
rect 322198 86232 322204 86244
rect 322256 86232 322262 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 17218 85524 17224 85536
rect 3200 85496 17224 85524
rect 3200 85484 3206 85496
rect 17218 85484 17224 85496
rect 17276 85484 17282 85536
rect 65978 85484 65984 85536
rect 66036 85524 66042 85536
rect 216674 85524 216680 85536
rect 66036 85496 216680 85524
rect 66036 85484 66042 85496
rect 216674 85484 216680 85496
rect 216732 85484 216738 85536
rect 101858 85416 101864 85468
rect 101916 85456 101922 85468
rect 213454 85456 213460 85468
rect 101916 85428 213460 85456
rect 101916 85416 101922 85428
rect 213454 85416 213460 85428
rect 213512 85416 213518 85468
rect 113358 85348 113364 85400
rect 113416 85388 113422 85400
rect 177482 85388 177488 85400
rect 113416 85360 177488 85388
rect 113416 85348 113422 85360
rect 177482 85348 177488 85360
rect 177540 85348 177546 85400
rect 114370 85280 114376 85332
rect 114428 85320 114434 85332
rect 171962 85320 171968 85332
rect 114428 85292 171968 85320
rect 114428 85280 114434 85292
rect 171962 85280 171968 85292
rect 172020 85280 172026 85332
rect 124030 85212 124036 85264
rect 124088 85252 124094 85264
rect 170582 85252 170588 85264
rect 124088 85224 170588 85252
rect 124088 85212 124094 85224
rect 170582 85212 170588 85224
rect 170640 85212 170646 85264
rect 319438 84804 319444 84856
rect 319496 84844 319502 84856
rect 333422 84844 333428 84856
rect 319496 84816 333428 84844
rect 319496 84804 319502 84816
rect 333422 84804 333428 84816
rect 333480 84804 333486 84856
rect 336090 84804 336096 84856
rect 336148 84844 336154 84856
rect 460934 84844 460940 84856
rect 336148 84816 460940 84844
rect 336148 84804 336154 84816
rect 460934 84804 460940 84816
rect 460992 84804 460998 84856
rect 107470 84124 107476 84176
rect 107528 84164 107534 84176
rect 187142 84164 187148 84176
rect 107528 84136 187148 84164
rect 107528 84124 107534 84136
rect 187142 84124 187148 84136
rect 187200 84124 187206 84176
rect 100662 84056 100668 84108
rect 100720 84096 100726 84108
rect 169294 84096 169300 84108
rect 100720 84068 169300 84096
rect 100720 84056 100726 84068
rect 169294 84056 169300 84068
rect 169352 84056 169358 84108
rect 106090 83988 106096 84040
rect 106148 84028 106154 84040
rect 167730 84028 167736 84040
rect 106148 84000 167736 84028
rect 106148 83988 106154 84000
rect 167730 83988 167736 84000
rect 167788 83988 167794 84040
rect 118602 83920 118608 83972
rect 118660 83960 118666 83972
rect 180242 83960 180248 83972
rect 118660 83932 180248 83960
rect 118660 83920 118666 83932
rect 180242 83920 180248 83932
rect 180300 83920 180306 83972
rect 124122 83852 124128 83904
rect 124180 83892 124186 83904
rect 174538 83892 174544 83904
rect 124180 83864 174544 83892
rect 124180 83852 124186 83864
rect 174538 83852 174544 83864
rect 174596 83852 174602 83904
rect 308490 83580 308496 83632
rect 308548 83620 308554 83632
rect 334710 83620 334716 83632
rect 308548 83592 334716 83620
rect 308548 83580 308554 83592
rect 334710 83580 334716 83592
rect 334768 83580 334774 83632
rect 207658 83512 207664 83564
rect 207716 83552 207722 83564
rect 331214 83552 331220 83564
rect 207716 83524 331220 83552
rect 207716 83512 207722 83524
rect 331214 83512 331220 83524
rect 331272 83552 331278 83564
rect 331272 83524 335354 83552
rect 331272 83512 331278 83524
rect 178770 83444 178776 83496
rect 178828 83484 178834 83496
rect 307110 83484 307116 83496
rect 178828 83456 307116 83484
rect 178828 83444 178834 83456
rect 307110 83444 307116 83456
rect 307168 83444 307174 83496
rect 335326 83484 335354 83524
rect 463786 83484 463792 83496
rect 335326 83456 463792 83484
rect 463786 83444 463792 83456
rect 463844 83444 463850 83496
rect 107562 82764 107568 82816
rect 107620 82804 107626 82816
rect 211890 82804 211896 82816
rect 107620 82776 211896 82804
rect 107620 82764 107626 82776
rect 211890 82764 211896 82776
rect 211948 82764 211954 82816
rect 119982 82696 119988 82748
rect 120040 82736 120046 82748
rect 198182 82736 198188 82748
rect 120040 82708 198188 82736
rect 120040 82696 120046 82708
rect 198182 82696 198188 82708
rect 198240 82696 198246 82748
rect 95050 82628 95056 82680
rect 95108 82668 95114 82680
rect 170674 82668 170680 82680
rect 95108 82640 170680 82668
rect 95108 82628 95114 82640
rect 170674 82628 170680 82640
rect 170732 82628 170738 82680
rect 104802 82560 104808 82612
rect 104860 82600 104866 82612
rect 173250 82600 173256 82612
rect 104860 82572 173256 82600
rect 104860 82560 104866 82572
rect 173250 82560 173256 82572
rect 173308 82560 173314 82612
rect 135162 82492 135168 82544
rect 135220 82532 135226 82544
rect 185578 82532 185584 82544
rect 135220 82504 185584 82532
rect 135220 82492 135226 82504
rect 185578 82492 185584 82504
rect 185636 82492 185642 82544
rect 206278 82084 206284 82136
rect 206336 82124 206342 82136
rect 261570 82124 261576 82136
rect 206336 82096 261576 82124
rect 206336 82084 206342 82096
rect 261570 82084 261576 82096
rect 261628 82084 261634 82136
rect 289170 82084 289176 82136
rect 289228 82124 289234 82136
rect 317414 82124 317420 82136
rect 289228 82096 317420 82124
rect 289228 82084 289234 82096
rect 317414 82084 317420 82096
rect 317472 82124 317478 82136
rect 466454 82124 466460 82136
rect 317472 82096 466460 82124
rect 317472 82084 317478 82096
rect 466454 82084 466460 82096
rect 466512 82084 466518 82136
rect 111702 81336 111708 81388
rect 111760 81376 111766 81388
rect 196894 81376 196900 81388
rect 111760 81348 196900 81376
rect 111760 81336 111766 81348
rect 196894 81336 196900 81348
rect 196952 81336 196958 81388
rect 125410 81268 125416 81320
rect 125468 81308 125474 81320
rect 209130 81308 209136 81320
rect 125468 81280 209136 81308
rect 125468 81268 125474 81280
rect 209130 81268 209136 81280
rect 209188 81268 209194 81320
rect 97810 81200 97816 81252
rect 97868 81240 97874 81252
rect 180150 81240 180156 81252
rect 97868 81212 180156 81240
rect 97868 81200 97874 81212
rect 180150 81200 180156 81212
rect 180208 81200 180214 81252
rect 93762 81132 93768 81184
rect 93820 81172 93826 81184
rect 167638 81172 167644 81184
rect 93820 81144 167644 81172
rect 93820 81132 93826 81144
rect 167638 81132 167644 81144
rect 167696 81132 167702 81184
rect 209038 80656 209044 80708
rect 209096 80696 209102 80708
rect 278038 80696 278044 80708
rect 209096 80668 278044 80696
rect 209096 80656 209102 80668
rect 278038 80656 278044 80668
rect 278096 80656 278102 80708
rect 309870 80656 309876 80708
rect 309928 80696 309934 80708
rect 470594 80696 470600 80708
rect 309928 80668 470600 80696
rect 309928 80656 309934 80668
rect 470594 80656 470600 80668
rect 470652 80656 470658 80708
rect 204898 79976 204904 80028
rect 204956 80016 204962 80028
rect 325694 80016 325700 80028
rect 204956 79988 325700 80016
rect 204956 79976 204962 79988
rect 325694 79976 325700 79988
rect 325752 80016 325758 80028
rect 326338 80016 326344 80028
rect 325752 79988 326344 80016
rect 325752 79976 325758 79988
rect 326338 79976 326344 79988
rect 326396 79976 326402 80028
rect 92382 79908 92388 79960
rect 92440 79948 92446 79960
rect 176010 79948 176016 79960
rect 92440 79920 176016 79948
rect 92440 79908 92446 79920
rect 176010 79908 176016 79920
rect 176068 79908 176074 79960
rect 125502 79840 125508 79892
rect 125560 79880 125566 79892
rect 202322 79880 202328 79892
rect 125560 79852 202328 79880
rect 125560 79840 125566 79852
rect 202322 79840 202328 79852
rect 202380 79840 202386 79892
rect 113082 79772 113088 79824
rect 113140 79812 113146 79824
rect 206462 79812 206468 79824
rect 113140 79784 206468 79812
rect 113140 79772 113146 79784
rect 206462 79772 206468 79784
rect 206520 79772 206526 79824
rect 202138 79364 202144 79416
rect 202196 79404 202202 79416
rect 246298 79404 246304 79416
rect 202196 79376 246304 79404
rect 202196 79364 202202 79376
rect 246298 79364 246304 79376
rect 246356 79364 246362 79416
rect 184198 79296 184204 79348
rect 184256 79336 184262 79348
rect 303614 79336 303620 79348
rect 184256 79308 303620 79336
rect 184256 79296 184262 79308
rect 303614 79296 303620 79308
rect 303672 79336 303678 79348
rect 471974 79336 471980 79348
rect 303672 79308 471980 79336
rect 303672 79296 303678 79308
rect 471974 79296 471980 79308
rect 472032 79296 472038 79348
rect 115750 78616 115756 78668
rect 115808 78656 115814 78668
rect 210510 78656 210516 78668
rect 115808 78628 210516 78656
rect 115808 78616 115814 78628
rect 210510 78616 210516 78628
rect 210568 78616 210574 78668
rect 95142 78548 95148 78600
rect 95200 78588 95206 78600
rect 174722 78588 174728 78600
rect 95200 78560 174728 78588
rect 95200 78548 95206 78560
rect 174722 78548 174728 78560
rect 174780 78548 174786 78600
rect 102042 78480 102048 78532
rect 102100 78520 102106 78532
rect 171870 78520 171876 78532
rect 102100 78492 171876 78520
rect 102100 78480 102106 78492
rect 171870 78480 171876 78492
rect 171928 78480 171934 78532
rect 121362 78412 121368 78464
rect 121420 78452 121426 78464
rect 184382 78452 184388 78464
rect 121420 78424 184388 78452
rect 121420 78412 121426 78424
rect 184382 78412 184388 78424
rect 184440 78412 184446 78464
rect 249150 78004 249156 78056
rect 249208 78044 249214 78056
rect 355318 78044 355324 78056
rect 249208 78016 355324 78044
rect 249208 78004 249214 78016
rect 355318 78004 355324 78016
rect 355376 78004 355382 78056
rect 310514 77936 310520 77988
rect 310572 77976 310578 77988
rect 469214 77976 469220 77988
rect 310572 77948 469220 77976
rect 310572 77936 310578 77948
rect 469214 77936 469220 77948
rect 469272 77936 469278 77988
rect 85482 77188 85488 77240
rect 85540 77228 85546 77240
rect 177574 77228 177580 77240
rect 85540 77200 177580 77228
rect 85540 77188 85546 77200
rect 177574 77188 177580 77200
rect 177632 77188 177638 77240
rect 297358 77188 297364 77240
rect 297416 77228 297422 77240
rect 329834 77228 329840 77240
rect 297416 77200 329840 77228
rect 297416 77188 297422 77200
rect 329834 77188 329840 77200
rect 329892 77228 329898 77240
rect 330478 77228 330484 77240
rect 329892 77200 330484 77228
rect 329892 77188 329898 77200
rect 330478 77188 330484 77200
rect 330536 77188 330542 77240
rect 110322 77120 110328 77172
rect 110380 77160 110386 77172
rect 175918 77160 175924 77172
rect 110380 77132 175924 77160
rect 110380 77120 110386 77132
rect 175918 77120 175924 77132
rect 175976 77120 175982 77172
rect 177298 76508 177304 76560
rect 177356 76548 177362 76560
rect 254670 76548 254676 76560
rect 177356 76520 254676 76548
rect 177356 76508 177362 76520
rect 254670 76508 254676 76520
rect 254728 76508 254734 76560
rect 324958 76508 324964 76560
rect 325016 76548 325022 76560
rect 463878 76548 463884 76560
rect 325016 76520 463884 76548
rect 325016 76508 325022 76520
rect 463878 76508 463884 76520
rect 463936 76508 463942 76560
rect 122098 75828 122104 75880
rect 122156 75868 122162 75880
rect 199562 75868 199568 75880
rect 122156 75840 199568 75868
rect 122156 75828 122162 75840
rect 199562 75828 199568 75840
rect 199620 75828 199626 75880
rect 93854 75216 93860 75268
rect 93912 75256 93918 75268
rect 300394 75256 300400 75268
rect 93912 75228 300400 75256
rect 93912 75216 93918 75228
rect 300394 75216 300400 75228
rect 300452 75216 300458 75268
rect 69014 75148 69020 75200
rect 69072 75188 69078 75200
rect 299014 75188 299020 75200
rect 69072 75160 299020 75188
rect 69072 75148 69078 75160
rect 299014 75148 299020 75160
rect 299072 75148 299078 75200
rect 300118 75148 300124 75200
rect 300176 75188 300182 75200
rect 473354 75188 473360 75200
rect 300176 75160 473360 75188
rect 300176 75148 300182 75160
rect 473354 75148 473360 75160
rect 473412 75148 473418 75200
rect 51718 74468 51724 74520
rect 51776 74508 51782 74520
rect 502334 74508 502340 74520
rect 51776 74480 502340 74508
rect 51776 74468 51782 74480
rect 502334 74468 502340 74480
rect 502392 74468 502398 74520
rect 104894 73856 104900 73908
rect 104952 73896 104958 73908
rect 246482 73896 246488 73908
rect 104952 73868 246488 73896
rect 104952 73856 104958 73868
rect 246482 73856 246488 73868
rect 246540 73856 246546 73908
rect 102134 73788 102140 73840
rect 102192 73828 102198 73840
rect 297634 73828 297640 73840
rect 102192 73800 297640 73828
rect 102192 73788 102198 73800
rect 297634 73788 297640 73800
rect 297692 73788 297698 73840
rect 63126 73108 63132 73160
rect 63184 73148 63190 73160
rect 335354 73148 335360 73160
rect 63184 73120 335360 73148
rect 63184 73108 63190 73120
rect 335354 73108 335360 73120
rect 335412 73148 335418 73160
rect 336090 73148 336096 73160
rect 335412 73120 336096 73148
rect 335412 73108 335418 73120
rect 336090 73108 336096 73120
rect 336148 73108 336154 73160
rect 419350 73108 419356 73160
rect 419408 73148 419414 73160
rect 579982 73148 579988 73160
rect 419408 73120 579988 73148
rect 419408 73108 419414 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 338758 73040 338764 73092
rect 338816 73080 338822 73092
rect 422294 73080 422300 73092
rect 338816 73052 422300 73080
rect 338816 73040 338822 73052
rect 422294 73040 422300 73052
rect 422352 73040 422358 73092
rect 33134 72428 33140 72480
rect 33192 72468 33198 72480
rect 304442 72468 304448 72480
rect 33192 72440 304448 72468
rect 33192 72428 33198 72440
rect 304442 72428 304448 72440
rect 304500 72428 304506 72480
rect 338114 71748 338120 71800
rect 338172 71788 338178 71800
rect 338758 71788 338764 71800
rect 338172 71760 338764 71788
rect 338172 71748 338178 71760
rect 338758 71748 338764 71760
rect 338816 71748 338822 71800
rect 3418 71612 3424 71664
rect 3476 71652 3482 71664
rect 7558 71652 7564 71664
rect 3476 71624 7564 71652
rect 3476 71612 3482 71624
rect 7558 71612 7564 71624
rect 7616 71612 7622 71664
rect 297358 71136 297364 71188
rect 297416 71176 297422 71188
rect 461578 71176 461584 71188
rect 297416 71148 461584 71176
rect 297416 71136 297422 71148
rect 461578 71136 461584 71148
rect 461636 71136 461642 71188
rect 115934 71068 115940 71120
rect 115992 71108 115998 71120
rect 297542 71108 297548 71120
rect 115992 71080 297548 71108
rect 115992 71068 115998 71080
rect 297542 71068 297548 71080
rect 297600 71068 297606 71120
rect 89714 71000 89720 71052
rect 89772 71040 89778 71052
rect 305914 71040 305920 71052
rect 89772 71012 305920 71040
rect 89772 71000 89778 71012
rect 305914 71000 305920 71012
rect 305972 71000 305978 71052
rect 293218 69708 293224 69760
rect 293276 69748 293282 69760
rect 474734 69748 474740 69760
rect 293276 69720 474740 69748
rect 293276 69708 293282 69720
rect 474734 69708 474740 69720
rect 474792 69708 474798 69760
rect 86954 69640 86960 69692
rect 87012 69680 87018 69692
rect 296254 69680 296260 69692
rect 87012 69652 296260 69680
rect 87012 69640 87018 69652
rect 296254 69640 296260 69652
rect 296312 69640 296318 69692
rect 122834 68416 122840 68468
rect 122892 68456 122898 68468
rect 276934 68456 276940 68468
rect 122892 68428 276940 68456
rect 122892 68416 122898 68428
rect 276934 68416 276940 68428
rect 276992 68416 276998 68468
rect 75914 68348 75920 68400
rect 75972 68388 75978 68400
rect 256142 68388 256148 68400
rect 75972 68360 256148 68388
rect 75972 68348 75978 68360
rect 256142 68348 256148 68360
rect 256200 68348 256206 68400
rect 291102 68348 291108 68400
rect 291160 68388 291166 68400
rect 476114 68388 476120 68400
rect 291160 68360 476120 68388
rect 291160 68348 291166 68360
rect 476114 68348 476120 68360
rect 476172 68348 476178 68400
rect 88978 68280 88984 68332
rect 89036 68320 89042 68332
rect 307018 68320 307024 68332
rect 89036 68292 307024 68320
rect 89036 68280 89042 68292
rect 307018 68280 307024 68292
rect 307076 68280 307082 68332
rect 203518 67532 203524 67584
rect 203576 67572 203582 67584
rect 289814 67572 289820 67584
rect 203576 67544 289820 67572
rect 203576 67532 203582 67544
rect 289814 67532 289820 67544
rect 289872 67572 289878 67584
rect 291102 67572 291108 67584
rect 289872 67544 291108 67572
rect 289872 67532 289878 67544
rect 291102 67532 291108 67544
rect 291160 67532 291166 67584
rect 22094 66852 22100 66904
rect 22152 66892 22158 66904
rect 290550 66892 290556 66904
rect 22152 66864 290556 66892
rect 22152 66852 22158 66864
rect 290550 66852 290556 66864
rect 290608 66852 290614 66904
rect 14 66172 20 66224
rect 72 66212 78 66224
rect 1302 66212 1308 66224
rect 72 66184 1308 66212
rect 72 66172 78 66184
rect 1302 66172 1308 66184
rect 1360 66212 1366 66224
rect 251910 66212 251916 66224
rect 1360 66184 251916 66212
rect 1360 66172 1366 66184
rect 251910 66172 251916 66184
rect 251968 66172 251974 66224
rect 279418 66172 279424 66224
rect 279476 66212 279482 66224
rect 480254 66212 480260 66224
rect 279476 66184 480260 66212
rect 279476 66172 279482 66184
rect 480254 66172 480260 66184
rect 480312 66172 480318 66224
rect 332594 66104 332600 66156
rect 332652 66144 332658 66156
rect 385678 66144 385684 66156
rect 332652 66116 385684 66144
rect 332652 66104 332658 66116
rect 385678 66104 385684 66116
rect 385736 66104 385742 66156
rect 260098 65668 260104 65680
rect 238726 65640 260104 65668
rect 106274 65560 106280 65612
rect 106332 65600 106338 65612
rect 238726 65600 238754 65640
rect 260098 65628 260104 65640
rect 260156 65628 260162 65680
rect 106332 65572 238754 65600
rect 106332 65560 106338 65572
rect 259546 65560 259552 65612
rect 259604 65600 259610 65612
rect 334618 65600 334624 65612
rect 259604 65572 334624 65600
rect 259604 65560 259610 65572
rect 334618 65560 334624 65572
rect 334676 65560 334682 65612
rect 73154 65492 73160 65544
rect 73212 65532 73218 65544
rect 279602 65532 279608 65544
rect 73212 65504 279608 65532
rect 73212 65492 73218 65504
rect 279602 65492 279608 65504
rect 279660 65492 279666 65544
rect 278774 65424 278780 65476
rect 278832 65464 278838 65476
rect 279418 65464 279424 65476
rect 278832 65436 279424 65464
rect 278832 65424 278838 65436
rect 279418 65424 279424 65436
rect 279476 65424 279482 65476
rect 272518 64812 272524 64864
rect 272576 64852 272582 64864
rect 481634 64852 481640 64864
rect 272576 64824 481640 64852
rect 272576 64812 272582 64824
rect 481634 64812 481640 64824
rect 481692 64812 481698 64864
rect 6914 64132 6920 64184
rect 6972 64172 6978 64184
rect 281074 64172 281080 64184
rect 6972 64144 281080 64172
rect 6972 64132 6978 64144
rect 281074 64132 281080 64144
rect 281132 64132 281138 64184
rect 271874 63520 271880 63572
rect 271932 63560 271938 63572
rect 272518 63560 272524 63572
rect 271932 63532 272524 63560
rect 271932 63520 271938 63532
rect 272518 63520 272524 63532
rect 272576 63520 272582 63572
rect 46934 62840 46940 62892
rect 46992 62880 46998 62892
rect 258810 62880 258816 62892
rect 46992 62852 258816 62880
rect 46992 62840 46998 62852
rect 258810 62840 258816 62852
rect 258868 62840 258874 62892
rect 267734 62840 267740 62892
rect 267792 62880 267798 62892
rect 483014 62880 483020 62892
rect 267792 62852 483020 62880
rect 267792 62840 267798 62852
rect 483014 62840 483020 62852
rect 483072 62840 483078 62892
rect 70394 62772 70400 62824
rect 70452 62812 70458 62824
rect 285122 62812 285128 62824
rect 70452 62784 285128 62812
rect 70452 62772 70458 62784
rect 285122 62772 285128 62784
rect 285180 62772 285186 62824
rect 264974 62024 264980 62076
rect 265032 62064 265038 62076
rect 265618 62064 265624 62076
rect 265032 62036 265624 62064
rect 265032 62024 265038 62036
rect 265618 62024 265624 62036
rect 265676 62064 265682 62076
rect 484394 62064 484400 62076
rect 265676 62036 484400 62064
rect 265676 62024 265682 62036
rect 484394 62024 484400 62036
rect 484452 62024 484458 62076
rect 74534 61412 74540 61464
rect 74592 61452 74598 61464
rect 286502 61452 286508 61464
rect 74592 61424 286508 61452
rect 74592 61412 74598 61424
rect 286502 61412 286508 61424
rect 286560 61412 286566 61464
rect 53834 61344 53840 61396
rect 53892 61384 53898 61396
rect 271322 61384 271328 61396
rect 53892 61356 271328 61384
rect 53892 61344 53898 61356
rect 271322 61344 271328 61356
rect 271380 61344 271386 61396
rect 261570 60664 261576 60716
rect 261628 60704 261634 60716
rect 485774 60704 485780 60716
rect 261628 60676 485780 60704
rect 261628 60664 261634 60676
rect 485774 60664 485780 60676
rect 485832 60664 485838 60716
rect 515398 60664 515404 60716
rect 515456 60704 515462 60716
rect 580166 60704 580172 60716
rect 515456 60676 580172 60704
rect 515456 60664 515462 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 260834 60256 260840 60308
rect 260892 60296 260898 60308
rect 261570 60296 261576 60308
rect 260892 60268 261576 60296
rect 260892 60256 260898 60268
rect 261570 60256 261576 60268
rect 261628 60256 261634 60308
rect 111794 60120 111800 60172
rect 111852 60160 111858 60172
rect 303062 60160 303068 60172
rect 111852 60132 303068 60160
rect 111852 60120 111858 60132
rect 303062 60120 303068 60132
rect 303120 60120 303126 60172
rect 64874 60052 64880 60104
rect 64932 60092 64938 60104
rect 261478 60092 261484 60104
rect 64932 60064 261484 60092
rect 64932 60052 64938 60064
rect 261478 60052 261484 60064
rect 261536 60052 261542 60104
rect 4154 59984 4160 60036
rect 4212 60024 4218 60036
rect 251818 60024 251824 60036
rect 4212 59996 251824 60024
rect 4212 59984 4218 59996
rect 251818 59984 251824 59996
rect 251876 59984 251882 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 21358 59344 21364 59356
rect 3108 59316 21364 59344
rect 3108 59304 3114 59316
rect 21358 59304 21364 59316
rect 21416 59304 21422 59356
rect 85574 58760 85580 58812
rect 85632 58800 85638 58812
rect 282454 58800 282460 58812
rect 85632 58772 282460 58800
rect 85632 58760 85638 58772
rect 282454 58760 282460 58772
rect 282512 58760 282518 58812
rect 259362 58692 259368 58744
rect 259420 58732 259426 58744
rect 488534 58732 488540 58744
rect 259420 58704 488540 58732
rect 259420 58692 259426 58704
rect 488534 58692 488540 58704
rect 488592 58692 488598 58744
rect 69106 58624 69112 58676
rect 69164 58664 69170 58676
rect 303154 58664 303160 58676
rect 69164 58636 303160 58664
rect 69164 58624 69170 58636
rect 303154 58624 303160 58636
rect 303212 58624 303218 58676
rect 254670 57944 254676 57996
rect 254728 57984 254734 57996
rect 259362 57984 259368 57996
rect 254728 57956 259368 57984
rect 254728 57944 254734 57956
rect 259362 57944 259368 57956
rect 259420 57944 259426 57996
rect 71774 57264 71780 57316
rect 71832 57304 71838 57316
rect 264330 57304 264336 57316
rect 71832 57276 264336 57304
rect 71832 57264 71838 57276
rect 264330 57264 264336 57276
rect 264388 57264 264394 57316
rect 246390 57196 246396 57248
rect 246448 57236 246454 57248
rect 251266 57236 251272 57248
rect 246448 57208 251272 57236
rect 246448 57196 246454 57208
rect 251266 57196 251272 57208
rect 251324 57236 251330 57248
rect 489914 57236 489920 57248
rect 251324 57208 489920 57236
rect 251324 57196 251330 57208
rect 489914 57196 489920 57208
rect 489972 57196 489978 57248
rect 93946 55972 93952 56024
rect 94004 56012 94010 56024
rect 268470 56012 268476 56024
rect 94004 55984 268476 56012
rect 94004 55972 94010 55984
rect 268470 55972 268476 55984
rect 268528 55972 268534 56024
rect 263594 55904 263600 55956
rect 263652 55944 263658 55956
rect 491294 55944 491300 55956
rect 263652 55916 491300 55944
rect 263652 55904 263658 55916
rect 491294 55904 491300 55916
rect 491352 55904 491358 55956
rect 18598 55836 18604 55888
rect 18656 55876 18662 55888
rect 307386 55876 307392 55888
rect 18656 55848 307392 55876
rect 18656 55836 18662 55848
rect 307386 55836 307392 55848
rect 307444 55836 307450 55888
rect 110414 54680 110420 54732
rect 110472 54720 110478 54732
rect 250622 54720 250628 54732
rect 110472 54692 250628 54720
rect 110472 54680 110478 54692
rect 250622 54680 250628 54692
rect 250680 54680 250686 54732
rect 82814 54612 82820 54664
rect 82872 54652 82878 54664
rect 275462 54652 275468 54664
rect 82872 54624 275468 54652
rect 82872 54612 82878 54624
rect 275462 54612 275468 54624
rect 275520 54612 275526 54664
rect 243538 54544 243544 54596
rect 243596 54584 243602 54596
rect 475378 54584 475384 54596
rect 243596 54556 475384 54584
rect 243596 54544 243602 54556
rect 475378 54544 475384 54556
rect 475436 54544 475442 54596
rect 15194 54476 15200 54528
rect 15252 54516 15258 54528
rect 307202 54516 307208 54528
rect 15252 54488 307208 54516
rect 15252 54476 15258 54488
rect 307202 54476 307208 54488
rect 307260 54476 307266 54528
rect 117314 53184 117320 53236
rect 117372 53224 117378 53236
rect 294874 53224 294880 53236
rect 117372 53196 294880 53224
rect 117372 53184 117378 53196
rect 294874 53184 294880 53196
rect 294932 53184 294938 53236
rect 35802 53116 35808 53168
rect 35860 53156 35866 53168
rect 132494 53156 132500 53168
rect 35860 53128 132500 53156
rect 35860 53116 35866 53128
rect 132494 53116 132500 53128
rect 132552 53116 132558 53168
rect 240778 53116 240784 53168
rect 240836 53156 240842 53168
rect 492674 53156 492680 53168
rect 240836 53128 492680 53156
rect 240836 53116 240842 53128
rect 492674 53116 492680 53128
rect 492732 53116 492738 53168
rect 11054 53048 11060 53100
rect 11112 53088 11118 53100
rect 267090 53088 267096 53100
rect 11112 53060 267096 53088
rect 11112 53048 11118 53060
rect 267090 53048 267096 53060
rect 267148 53048 267154 53100
rect 349798 52368 349804 52420
rect 349856 52408 349862 52420
rect 495526 52408 495532 52420
rect 349856 52380 495532 52408
rect 349856 52368 349862 52380
rect 495526 52368 495532 52380
rect 495584 52368 495590 52420
rect 204990 51824 204996 51876
rect 205048 51864 205054 51876
rect 241514 51864 241520 51876
rect 205048 51836 241520 51864
rect 205048 51824 205054 51836
rect 241514 51824 241520 51836
rect 241572 51864 241578 51876
rect 360930 51864 360936 51876
rect 241572 51836 360936 51864
rect 241572 51824 241578 51836
rect 360930 51824 360936 51836
rect 360988 51824 360994 51876
rect 120074 51756 120080 51808
rect 120132 51796 120138 51808
rect 249058 51796 249064 51808
rect 120132 51768 249064 51796
rect 120132 51756 120138 51768
rect 249058 51756 249064 51768
rect 249116 51756 249122 51808
rect 114554 51688 114560 51740
rect 114612 51728 114618 51740
rect 292022 51728 292028 51740
rect 114612 51700 292028 51728
rect 114612 51688 114618 51700
rect 292022 51688 292028 51700
rect 292080 51688 292086 51740
rect 349154 51076 349160 51128
rect 349212 51116 349218 51128
rect 349798 51116 349804 51128
rect 349212 51088 349804 51116
rect 349212 51076 349218 51088
rect 349798 51076 349804 51088
rect 349856 51076 349862 51128
rect 244274 50532 244280 50584
rect 244332 50572 244338 50584
rect 356698 50572 356704 50584
rect 244332 50544 356704 50572
rect 244332 50532 244338 50544
rect 356698 50532 356704 50544
rect 356756 50532 356762 50584
rect 113174 50464 113180 50516
rect 113232 50504 113238 50516
rect 253290 50504 253296 50516
rect 113232 50476 253296 50504
rect 113232 50464 113238 50476
rect 253290 50464 253296 50476
rect 253348 50464 253354 50516
rect 85666 50396 85672 50448
rect 85724 50436 85730 50448
rect 300302 50436 300308 50448
rect 85724 50408 300308 50436
rect 85724 50396 85730 50408
rect 300302 50396 300308 50408
rect 300360 50396 300366 50448
rect 19334 50328 19340 50380
rect 19392 50368 19398 50380
rect 249242 50368 249248 50380
rect 19392 50340 249248 50368
rect 19392 50328 19398 50340
rect 249242 50328 249248 50340
rect 249300 50328 249306 50380
rect 192478 49648 192484 49700
rect 192536 49688 192542 49700
rect 244274 49688 244280 49700
rect 192536 49660 244280 49688
rect 192536 49648 192542 49660
rect 244274 49648 244280 49660
rect 244332 49648 244338 49700
rect 358814 49648 358820 49700
rect 358872 49688 358878 49700
rect 359274 49688 359280 49700
rect 358872 49660 359280 49688
rect 358872 49648 358878 49660
rect 359274 49648 359280 49660
rect 359332 49688 359338 49700
rect 494146 49688 494152 49700
rect 359332 49660 494152 49688
rect 359332 49648 359338 49660
rect 494146 49648 494152 49660
rect 494204 49648 494210 49700
rect 99374 49036 99380 49088
rect 99432 49076 99438 49088
rect 304258 49076 304264 49088
rect 99432 49048 304264 49076
rect 99432 49036 99438 49048
rect 304258 49036 304264 49048
rect 304316 49036 304322 49088
rect 340874 49036 340880 49088
rect 340932 49076 340938 49088
rect 359274 49076 359280 49088
rect 340932 49048 359280 49076
rect 340932 49036 340938 49048
rect 359274 49036 359280 49048
rect 359332 49036 359338 49088
rect 11146 48968 11152 49020
rect 11204 49008 11210 49020
rect 11204 48980 277394 49008
rect 11204 48968 11210 48980
rect 277366 48940 277394 48980
rect 284386 48968 284392 49020
rect 284444 49008 284450 49020
rect 341518 49008 341524 49020
rect 284444 48980 341524 49008
rect 284444 48968 284450 48980
rect 341518 48968 341524 48980
rect 341576 48968 341582 49020
rect 285214 48940 285220 48952
rect 277366 48912 285220 48940
rect 285214 48900 285220 48912
rect 285272 48900 285278 48952
rect 343634 48220 343640 48272
rect 343692 48260 343698 48272
rect 344278 48260 344284 48272
rect 343692 48232 344284 48260
rect 343692 48220 343698 48232
rect 344278 48220 344284 48232
rect 344336 48260 344342 48272
rect 498194 48260 498200 48272
rect 344336 48232 498200 48260
rect 344336 48220 344342 48232
rect 498194 48220 498200 48232
rect 498252 48220 498258 48272
rect 118694 47608 118700 47660
rect 118752 47648 118758 47660
rect 298922 47648 298928 47660
rect 118752 47620 298928 47648
rect 118752 47608 118758 47620
rect 298922 47608 298928 47620
rect 298980 47608 298986 47660
rect 23474 47540 23480 47592
rect 23532 47580 23538 47592
rect 269850 47580 269856 47592
rect 23532 47552 269856 47580
rect 23532 47540 23538 47552
rect 269850 47540 269856 47552
rect 269908 47540 269914 47592
rect 340230 47580 340236 47592
rect 277366 47552 340236 47580
rect 269114 47472 269120 47524
rect 269172 47512 269178 47524
rect 277366 47512 277394 47552
rect 340230 47540 340236 47552
rect 340288 47540 340294 47592
rect 269172 47484 277394 47512
rect 269172 47472 269178 47484
rect 544378 46860 544384 46912
rect 544436 46900 544442 46912
rect 580166 46900 580172 46912
rect 544436 46872 580172 46900
rect 544436 46860 544442 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 284938 46248 284944 46300
rect 284996 46288 285002 46300
rect 352558 46288 352564 46300
rect 284996 46260 352564 46288
rect 284996 46248 285002 46260
rect 352558 46248 352564 46260
rect 352616 46248 352622 46300
rect 26234 46180 26240 46232
rect 26292 46220 26298 46232
rect 271230 46220 271236 46232
rect 26292 46192 271236 46220
rect 26292 46180 26298 46192
rect 271230 46180 271236 46192
rect 271288 46180 271294 46232
rect 334066 46180 334072 46232
rect 334124 46220 334130 46232
rect 494422 46220 494428 46232
rect 334124 46192 494428 46220
rect 334124 46180 334130 46192
rect 494422 46180 494428 46192
rect 494480 46180 494486 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 29638 45540 29644 45552
rect 3476 45512 29644 45540
rect 3476 45500 3482 45512
rect 29638 45500 29644 45512
rect 29696 45500 29702 45552
rect 280890 45500 280896 45552
rect 280948 45540 280954 45552
rect 335998 45540 336004 45552
rect 280948 45512 336004 45540
rect 280948 45500 280954 45512
rect 335998 45500 336004 45512
rect 336056 45500 336062 45552
rect 95234 44956 95240 45008
rect 95292 44996 95298 45008
rect 250438 44996 250444 45008
rect 95292 44968 250444 44996
rect 95292 44956 95298 44968
rect 250438 44956 250444 44968
rect 250496 44956 250502 45008
rect 121454 44888 121460 44940
rect 121512 44928 121518 44940
rect 297450 44928 297456 44940
rect 121512 44900 297456 44928
rect 121512 44888 121518 44900
rect 297450 44888 297456 44900
rect 297508 44888 297514 44940
rect 27614 44820 27620 44872
rect 27672 44860 27678 44872
rect 285030 44860 285036 44872
rect 27672 44832 285036 44860
rect 27672 44820 27678 44832
rect 285030 44820 285036 44832
rect 285088 44820 285094 44872
rect 316770 44820 316776 44872
rect 316828 44860 316834 44872
rect 427814 44860 427820 44872
rect 316828 44832 427820 44860
rect 316828 44820 316834 44832
rect 427814 44820 427820 44832
rect 427872 44820 427878 44872
rect 280154 44140 280160 44192
rect 280212 44180 280218 44192
rect 280890 44180 280896 44192
rect 280212 44152 280896 44180
rect 280212 44140 280218 44152
rect 280890 44140 280896 44152
rect 280948 44140 280954 44192
rect 92474 43460 92480 43512
rect 92532 43500 92538 43512
rect 298830 43500 298836 43512
rect 92532 43472 298836 43500
rect 92532 43460 92538 43472
rect 298830 43460 298836 43472
rect 298888 43460 298894 43512
rect 320082 43460 320088 43512
rect 320140 43500 320146 43512
rect 429194 43500 429200 43512
rect 320140 43472 429200 43500
rect 320140 43460 320146 43472
rect 429194 43460 429200 43472
rect 429252 43460 429258 43512
rect 57974 43392 57980 43444
rect 58032 43432 58038 43444
rect 286594 43432 286600 43444
rect 58032 43404 286600 43432
rect 58032 43392 58038 43404
rect 286594 43392 286600 43404
rect 286652 43392 286658 43444
rect 298186 43392 298192 43444
rect 298244 43432 298250 43444
rect 331858 43432 331864 43444
rect 298244 43404 331864 43432
rect 298244 43392 298250 43404
rect 331858 43392 331864 43404
rect 331916 43392 331922 43444
rect 342990 43392 342996 43444
rect 343048 43432 343054 43444
rect 462314 43432 462320 43444
rect 343048 43404 462320 43432
rect 343048 43392 343054 43404
rect 462314 43392 462320 43404
rect 462372 43392 462378 43444
rect 322198 42712 322204 42764
rect 322256 42752 322262 42764
rect 465074 42752 465080 42764
rect 322256 42724 465080 42752
rect 322256 42712 322262 42724
rect 465074 42712 465080 42724
rect 465132 42712 465138 42764
rect 276014 42644 276020 42696
rect 276072 42684 276078 42696
rect 276658 42684 276664 42696
rect 276072 42656 276664 42684
rect 276072 42644 276078 42656
rect 276658 42644 276664 42656
rect 276716 42684 276722 42696
rect 342898 42684 342904 42696
rect 276716 42656 342904 42684
rect 276716 42644 276722 42656
rect 342898 42644 342904 42656
rect 342956 42644 342962 42696
rect 38654 42100 38660 42152
rect 38712 42140 38718 42152
rect 264238 42140 264244 42152
rect 38712 42112 264244 42140
rect 38712 42100 38718 42112
rect 264238 42100 264244 42112
rect 264296 42100 264302 42152
rect 20714 42032 20720 42084
rect 20772 42072 20778 42084
rect 301774 42072 301780 42084
rect 20772 42044 301780 42072
rect 20772 42032 20778 42044
rect 301774 42032 301780 42044
rect 301832 42032 301838 42084
rect 321554 41420 321560 41472
rect 321612 41460 321618 41472
rect 322198 41460 322204 41472
rect 321612 41432 322204 41460
rect 321612 41420 321618 41432
rect 322198 41420 322204 41432
rect 322256 41420 322262 41472
rect 45554 40740 45560 40792
rect 45612 40780 45618 40792
rect 273990 40780 273996 40792
rect 45612 40752 273996 40780
rect 45612 40740 45618 40752
rect 273990 40740 273996 40752
rect 274048 40740 274054 40792
rect 35894 40672 35900 40724
rect 35952 40712 35958 40724
rect 300210 40712 300216 40724
rect 35952 40684 300216 40712
rect 35952 40672 35958 40684
rect 300210 40672 300216 40684
rect 300268 40672 300274 40724
rect 302234 40672 302240 40724
rect 302292 40712 302298 40724
rect 433334 40712 433340 40724
rect 302292 40684 433340 40712
rect 302292 40672 302298 40684
rect 433334 40672 433340 40684
rect 433392 40672 433398 40724
rect 280798 39992 280804 40044
rect 280856 40032 280862 40044
rect 296714 40032 296720 40044
rect 280856 40004 296720 40032
rect 280856 39992 280862 40004
rect 296714 39992 296720 40004
rect 296772 40032 296778 40044
rect 297358 40032 297364 40044
rect 296772 40004 297364 40032
rect 296772 39992 296778 40004
rect 297358 39992 297364 40004
rect 297416 39992 297422 40044
rect 59354 39380 59360 39432
rect 59412 39420 59418 39432
rect 304350 39420 304356 39432
rect 59412 39392 304356 39420
rect 59412 39380 59418 39392
rect 304350 39380 304356 39392
rect 304408 39380 304414 39432
rect 2774 39312 2780 39364
rect 2832 39352 2838 39364
rect 278314 39352 278320 39364
rect 2832 39324 278320 39352
rect 2832 39312 2838 39324
rect 278314 39312 278320 39324
rect 278372 39312 278378 39364
rect 299658 39312 299664 39364
rect 299716 39352 299722 39364
rect 434714 39352 434720 39364
rect 299716 39324 434720 39352
rect 299716 39312 299722 39324
rect 434714 39312 434720 39324
rect 434772 39312 434778 39364
rect 196618 38020 196624 38072
rect 196676 38060 196682 38072
rect 295334 38060 295340 38072
rect 196676 38032 295340 38060
rect 196676 38020 196682 38032
rect 295334 38020 295340 38032
rect 295392 38060 295398 38072
rect 295392 38032 296714 38060
rect 295392 38020 295398 38032
rect 91094 37952 91100 38004
rect 91152 37992 91158 38004
rect 272610 37992 272616 38004
rect 91152 37964 272616 37992
rect 91152 37952 91158 37964
rect 272610 37952 272616 37964
rect 272668 37952 272674 38004
rect 296686 37992 296714 38032
rect 436186 37992 436192 38004
rect 296686 37964 436192 37992
rect 436186 37952 436192 37964
rect 436244 37952 436250 38004
rect 16574 37884 16580 37936
rect 16632 37924 16638 37936
rect 296162 37924 296168 37936
rect 16632 37896 296168 37924
rect 16632 37884 16638 37896
rect 296162 37884 296168 37896
rect 296220 37884 296226 37936
rect 64690 37204 64696 37256
rect 64748 37244 64754 37256
rect 307754 37244 307760 37256
rect 64748 37216 307760 37244
rect 64748 37204 64754 37216
rect 307754 37204 307760 37216
rect 307812 37244 307818 37256
rect 308490 37244 308496 37256
rect 307812 37216 308496 37244
rect 307812 37204 307818 37216
rect 308490 37204 308496 37216
rect 308548 37204 308554 37256
rect 195238 36592 195244 36644
rect 195296 36632 195302 36644
rect 292574 36632 292580 36644
rect 195296 36604 292580 36632
rect 195296 36592 195302 36604
rect 292574 36592 292580 36604
rect 292632 36632 292638 36644
rect 436278 36632 436284 36644
rect 292632 36604 436284 36632
rect 292632 36592 292638 36604
rect 436278 36592 436284 36604
rect 436336 36592 436342 36644
rect 41414 36524 41420 36576
rect 41472 36564 41478 36576
rect 293310 36564 293316 36576
rect 41472 36536 293316 36564
rect 41472 36524 41478 36536
rect 293310 36524 293316 36536
rect 293368 36524 293374 36576
rect 37182 35232 37188 35284
rect 37240 35272 37246 35284
rect 135254 35272 135260 35284
rect 37240 35244 135260 35272
rect 37240 35232 37246 35244
rect 135254 35232 135260 35244
rect 135312 35232 135318 35284
rect 178678 35232 178684 35284
rect 178736 35272 178742 35284
rect 256050 35272 256056 35284
rect 178736 35244 256056 35272
rect 178736 35232 178742 35244
rect 256050 35232 256056 35244
rect 256108 35232 256114 35284
rect 28994 35164 29000 35216
rect 29052 35204 29058 35216
rect 287882 35204 287888 35216
rect 29052 35176 287888 35204
rect 29052 35164 29058 35176
rect 287882 35164 287888 35176
rect 287940 35164 287946 35216
rect 289722 35164 289728 35216
rect 289780 35204 289786 35216
rect 437474 35204 437480 35216
rect 289780 35176 437480 35204
rect 289780 35164 289786 35176
rect 437474 35164 437480 35176
rect 437532 35164 437538 35216
rect 184290 34416 184296 34468
rect 184348 34456 184354 34468
rect 288434 34456 288440 34468
rect 184348 34428 288440 34456
rect 184348 34416 184354 34428
rect 288434 34416 288440 34428
rect 288492 34456 288498 34468
rect 289722 34456 289728 34468
rect 288492 34428 289728 34456
rect 288492 34416 288498 34428
rect 289722 34416 289728 34428
rect 289780 34416 289786 34468
rect 60734 33736 60740 33788
rect 60792 33776 60798 33788
rect 289078 33776 289084 33788
rect 60792 33748 289084 33776
rect 60792 33736 60798 33748
rect 289078 33736 289084 33748
rect 289136 33736 289142 33788
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 51718 33096 51724 33108
rect 3568 33068 51724 33096
rect 3568 33056 3574 33068
rect 51718 33056 51724 33068
rect 51776 33056 51782 33108
rect 180058 33056 180064 33108
rect 180116 33096 180122 33108
rect 316126 33096 316132 33108
rect 180116 33068 316132 33096
rect 180116 33056 180122 33068
rect 316126 33056 316132 33068
rect 316184 33096 316190 33108
rect 316770 33096 316776 33108
rect 316184 33068 316776 33096
rect 316184 33056 316190 33068
rect 316770 33056 316776 33068
rect 316828 33056 316834 33108
rect 357434 33056 357440 33108
rect 357492 33096 357498 33108
rect 425054 33096 425060 33108
rect 357492 33068 425060 33096
rect 357492 33056 357498 33068
rect 425054 33056 425060 33068
rect 425112 33056 425118 33108
rect 291838 32988 291844 33040
rect 291896 33028 291902 33040
rect 356790 33028 356796 33040
rect 291896 33000 356796 33028
rect 291896 32988 291902 33000
rect 356790 32988 356796 33000
rect 356848 32988 356854 33040
rect 80054 32444 80060 32496
rect 80112 32484 80118 32496
rect 250530 32484 250536 32496
rect 80112 32456 250536 32484
rect 80112 32444 80118 32456
rect 250530 32444 250536 32456
rect 250588 32444 250594 32496
rect 62114 32376 62120 32428
rect 62172 32416 62178 32428
rect 283742 32416 283748 32428
rect 62172 32388 283748 32416
rect 62172 32376 62178 32388
rect 283742 32376 283748 32388
rect 283800 32376 283806 32428
rect 327074 32376 327080 32428
rect 327132 32416 327138 32428
rect 357434 32416 357440 32428
rect 327132 32388 357440 32416
rect 327132 32376 327138 32388
rect 357434 32376 357440 32388
rect 357492 32376 357498 32428
rect 291194 31764 291200 31816
rect 291252 31804 291258 31816
rect 291838 31804 291844 31816
rect 291252 31776 291844 31804
rect 291252 31764 291258 31776
rect 291838 31764 291844 31776
rect 291896 31764 291902 31816
rect 44174 31084 44180 31136
rect 44232 31124 44238 31136
rect 274082 31124 274088 31136
rect 44232 31096 274088 31124
rect 44232 31084 44238 31096
rect 274082 31084 274088 31096
rect 274140 31084 274146 31136
rect 282178 31084 282184 31136
rect 282236 31124 282242 31136
rect 438854 31124 438860 31136
rect 282236 31096 438860 31124
rect 282236 31084 282242 31096
rect 438854 31084 438860 31096
rect 438912 31084 438918 31136
rect 24854 31016 24860 31068
rect 24912 31056 24918 31068
rect 302970 31056 302976 31068
rect 24912 31028 302976 31056
rect 24912 31016 24918 31028
rect 302970 31016 302976 31028
rect 303028 31016 303034 31068
rect 277394 30268 277400 30320
rect 277452 30308 277458 30320
rect 278038 30308 278044 30320
rect 277452 30280 278044 30308
rect 277452 30268 277458 30280
rect 278038 30268 278044 30280
rect 278096 30308 278102 30320
rect 441614 30308 441620 30320
rect 278096 30280 441620 30308
rect 278096 30268 278102 30280
rect 441614 30268 441620 30280
rect 441672 30268 441678 30320
rect 52454 29656 52460 29708
rect 52512 29696 52518 29708
rect 265710 29696 265716 29708
rect 52512 29668 265716 29696
rect 52512 29656 52518 29668
rect 265710 29656 265716 29668
rect 265768 29656 265774 29708
rect 64782 29588 64788 29640
rect 64840 29628 64846 29640
rect 309962 29628 309968 29640
rect 64840 29600 309968 29628
rect 64840 29588 64846 29600
rect 309962 29588 309968 29600
rect 310020 29588 310026 29640
rect 81434 28228 81440 28280
rect 81492 28268 81498 28280
rect 275370 28268 275376 28280
rect 81492 28240 275376 28268
rect 81492 28228 81498 28240
rect 275370 28228 275376 28240
rect 275428 28228 275434 28280
rect 280798 28228 280804 28280
rect 280856 28268 280862 28280
rect 442994 28268 443000 28280
rect 280856 28240 443000 28268
rect 280856 28228 280862 28240
rect 442994 28228 443000 28240
rect 443052 28228 443058 28280
rect 51074 26868 51080 26920
rect 51132 26908 51138 26920
rect 255958 26908 255964 26920
rect 51132 26880 255964 26908
rect 51132 26868 51138 26880
rect 255958 26868 255964 26880
rect 256016 26868 256022 26920
rect 270586 26868 270592 26920
rect 270644 26908 270650 26920
rect 444374 26908 444380 26920
rect 270644 26880 444380 26908
rect 270644 26868 270650 26880
rect 444374 26868 444380 26880
rect 444432 26868 444438 26920
rect 196710 25644 196716 25696
rect 196768 25684 196774 25696
rect 274634 25684 274640 25696
rect 196768 25656 274640 25684
rect 196768 25644 196774 25656
rect 274634 25644 274640 25656
rect 274692 25684 274698 25696
rect 445846 25684 445852 25696
rect 274692 25656 445852 25684
rect 274692 25644 274698 25656
rect 445846 25644 445852 25656
rect 445904 25644 445910 25696
rect 35986 25576 35992 25628
rect 36044 25616 36050 25628
rect 276750 25616 276756 25628
rect 36044 25588 276756 25616
rect 36044 25576 36050 25588
rect 276750 25576 276756 25588
rect 276808 25576 276814 25628
rect 40034 25508 40040 25560
rect 40092 25548 40098 25560
rect 289262 25548 289268 25560
rect 40092 25520 289268 25548
rect 40092 25508 40098 25520
rect 289262 25508 289268 25520
rect 289320 25508 289326 25560
rect 118786 24216 118792 24268
rect 118844 24256 118850 24268
rect 286410 24256 286416 24268
rect 118844 24228 286416 24256
rect 118844 24216 118850 24228
rect 286410 24216 286416 24228
rect 286468 24216 286474 24268
rect 263686 24148 263692 24200
rect 263744 24188 263750 24200
rect 445938 24188 445944 24200
rect 263744 24160 445944 24188
rect 263744 24148 263750 24160
rect 445938 24148 445944 24160
rect 445996 24148 446002 24200
rect 48314 24080 48320 24132
rect 48372 24120 48378 24132
rect 266998 24120 267004 24132
rect 48372 24092 267004 24120
rect 48372 24080 48378 24092
rect 266998 24080 267004 24092
rect 267056 24080 267062 24132
rect 43438 23400 43444 23452
rect 43496 23440 43502 23452
rect 44082 23440 44088 23452
rect 43496 23412 44088 23440
rect 43496 23400 43502 23412
rect 44082 23400 44088 23412
rect 44140 23440 44146 23452
rect 249794 23440 249800 23452
rect 44140 23412 249800 23440
rect 44140 23400 44146 23412
rect 249794 23400 249800 23412
rect 249852 23400 249858 23452
rect 186958 22788 186964 22840
rect 187016 22828 187022 22840
rect 259454 22828 259460 22840
rect 187016 22800 259460 22828
rect 187016 22788 187022 22800
rect 259454 22788 259460 22800
rect 259512 22828 259518 22840
rect 447134 22828 447140 22840
rect 259512 22800 447140 22828
rect 259512 22788 259518 22800
rect 447134 22788 447140 22800
rect 447192 22788 447198 22840
rect 52546 22720 52552 22772
rect 52604 22760 52610 22772
rect 290458 22760 290464 22772
rect 52604 22732 290464 22760
rect 52604 22720 52610 22732
rect 290458 22720 290464 22732
rect 290516 22720 290522 22772
rect 253382 22040 253388 22092
rect 253440 22080 253446 22092
rect 449894 22080 449900 22092
rect 253440 22052 449900 22080
rect 253440 22040 253446 22052
rect 449894 22040 449900 22052
rect 449952 22040 449958 22092
rect 252554 21564 252560 21616
rect 252612 21604 252618 21616
rect 253382 21604 253388 21616
rect 252612 21576 253388 21604
rect 252612 21564 252618 21576
rect 253382 21564 253388 21576
rect 253440 21564 253446 21616
rect 30374 21360 30380 21412
rect 30432 21400 30438 21412
rect 280982 21400 280988 21412
rect 30432 21372 280988 21400
rect 30432 21360 30438 21372
rect 280982 21360 280988 21372
rect 281040 21360 281046 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 57238 20652 57244 20664
rect 3476 20624 57244 20652
rect 3476 20612 3482 20624
rect 57238 20612 57244 20624
rect 57296 20612 57302 20664
rect 64598 20612 64604 20664
rect 64656 20652 64662 20664
rect 64656 20624 238754 20652
rect 64656 20612 64662 20624
rect 238726 20584 238754 20624
rect 246298 20612 246304 20664
rect 246356 20652 246362 20664
rect 249794 20652 249800 20664
rect 246356 20624 249800 20652
rect 246356 20612 246362 20624
rect 249794 20612 249800 20624
rect 249852 20652 249858 20664
rect 250806 20652 250812 20664
rect 249852 20624 250812 20652
rect 249852 20612 249858 20624
rect 250806 20612 250812 20624
rect 250864 20612 250870 20664
rect 509142 20612 509148 20664
rect 509200 20652 509206 20664
rect 579982 20652 579988 20664
rect 509200 20624 579988 20652
rect 509200 20612 509206 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 248414 20584 248420 20596
rect 238726 20556 248420 20584
rect 248414 20544 248420 20556
rect 248472 20584 248478 20596
rect 249150 20584 249156 20596
rect 248472 20556 249156 20584
rect 248472 20544 248478 20556
rect 249150 20544 249156 20556
rect 249208 20544 249214 20596
rect 250806 20000 250812 20052
rect 250864 20040 250870 20052
rect 451274 20040 451280 20052
rect 250864 20012 451280 20040
rect 250864 20000 250870 20012
rect 451274 20000 451280 20012
rect 451332 20000 451338 20052
rect 56594 19932 56600 19984
rect 56652 19972 56658 19984
rect 278130 19972 278136 19984
rect 56652 19944 278136 19972
rect 56652 19932 56658 19944
rect 278130 19932 278136 19944
rect 278188 19932 278194 19984
rect 100754 18708 100760 18760
rect 100812 18748 100818 18760
rect 257430 18748 257436 18760
rect 100812 18720 257436 18748
rect 100812 18708 100818 18720
rect 257430 18708 257436 18720
rect 257488 18708 257494 18760
rect 246298 18640 246304 18692
rect 246356 18680 246362 18692
rect 452654 18680 452660 18692
rect 246356 18652 452660 18680
rect 246356 18640 246362 18652
rect 452654 18640 452660 18652
rect 452712 18640 452718 18692
rect 27706 18572 27712 18624
rect 27764 18612 27770 18624
rect 301682 18612 301688 18624
rect 27764 18584 301688 18612
rect 27764 18572 27770 18584
rect 301682 18572 301688 18584
rect 301740 18572 301746 18624
rect 103514 17280 103520 17332
rect 103572 17320 103578 17332
rect 302878 17320 302884 17332
rect 103572 17292 302884 17320
rect 103572 17280 103578 17292
rect 302878 17280 302884 17292
rect 302936 17280 302942 17332
rect 37274 17212 37280 17264
rect 37332 17252 37338 17264
rect 268378 17252 268384 17264
rect 37332 17224 268384 17252
rect 37332 17212 37338 17224
rect 268378 17212 268384 17224
rect 268436 17212 268442 17264
rect 271230 17212 271236 17264
rect 271288 17252 271294 17264
rect 454126 17252 454132 17264
rect 271288 17224 454132 17252
rect 271288 17212 271294 17224
rect 454126 17212 454132 17224
rect 454184 17212 454190 17264
rect 301498 16532 301504 16584
rect 301556 16572 301562 16584
rect 363598 16572 363604 16584
rect 301556 16544 363604 16572
rect 301556 16532 301562 16544
rect 363598 16532 363604 16544
rect 363656 16532 363662 16584
rect 108114 15920 108120 15972
rect 108172 15960 108178 15972
rect 279510 15960 279516 15972
rect 108172 15932 279516 15960
rect 108172 15920 108178 15932
rect 279510 15920 279516 15932
rect 279568 15920 279574 15972
rect 286410 15920 286416 15972
rect 286468 15960 286474 15972
rect 454034 15960 454040 15972
rect 286468 15932 454040 15960
rect 286468 15920 286474 15932
rect 454034 15920 454040 15932
rect 454092 15920 454098 15972
rect 19426 15852 19432 15904
rect 19484 15892 19490 15904
rect 287790 15892 287796 15904
rect 19484 15864 287796 15892
rect 19484 15852 19490 15864
rect 287790 15852 287796 15864
rect 287848 15852 287854 15904
rect 84194 14560 84200 14612
rect 84252 14600 84258 14612
rect 258718 14600 258724 14612
rect 84252 14572 258724 14600
rect 84252 14560 84258 14572
rect 258718 14560 258724 14572
rect 258776 14560 258782 14612
rect 66714 14492 66720 14544
rect 66772 14532 66778 14544
rect 305730 14532 305736 14544
rect 66772 14504 305736 14532
rect 66772 14492 66778 14504
rect 305730 14492 305736 14504
rect 305788 14492 305794 14544
rect 164418 14424 164424 14476
rect 164476 14464 164482 14476
rect 414658 14464 414664 14476
rect 164476 14436 414664 14464
rect 164476 14424 164482 14436
rect 414658 14424 414664 14436
rect 414716 14424 414722 14476
rect 314654 13744 314660 13796
rect 314712 13784 314718 13796
rect 315298 13784 315304 13796
rect 314712 13756 315304 13784
rect 314712 13744 314718 13756
rect 315298 13744 315304 13756
rect 315356 13784 315362 13796
rect 467834 13784 467840 13796
rect 315356 13756 467840 13784
rect 315356 13744 315362 13756
rect 467834 13744 467840 13756
rect 467892 13744 467898 13796
rect 255866 13676 255872 13728
rect 255924 13716 255930 13728
rect 256050 13716 256056 13728
rect 255924 13688 256056 13716
rect 255924 13676 255930 13688
rect 256050 13676 256056 13688
rect 256108 13716 256114 13728
rect 353938 13716 353944 13728
rect 256108 13688 353944 13716
rect 256108 13676 256114 13688
rect 353938 13676 353944 13688
rect 353996 13676 354002 13728
rect 191098 13200 191104 13252
rect 191156 13240 191162 13252
rect 257430 13240 257436 13252
rect 191156 13212 257436 13240
rect 191156 13200 191162 13212
rect 257430 13200 257436 13212
rect 257488 13200 257494 13252
rect 97442 13132 97448 13184
rect 97500 13172 97506 13184
rect 253198 13172 253204 13184
rect 97500 13144 253204 13172
rect 97500 13132 97506 13144
rect 253198 13132 253204 13144
rect 253256 13132 253262 13184
rect 56042 13064 56048 13116
rect 56100 13104 56106 13116
rect 305822 13104 305828 13116
rect 56100 13076 305828 13104
rect 56100 13064 56106 13076
rect 305822 13064 305828 13076
rect 305880 13064 305886 13116
rect 283098 12384 283104 12436
rect 283156 12424 283162 12436
rect 283558 12424 283564 12436
rect 283156 12396 283564 12424
rect 283156 12384 283162 12396
rect 283558 12384 283564 12396
rect 283616 12424 283622 12436
rect 478874 12424 478880 12436
rect 283616 12396 478880 12424
rect 283616 12384 283622 12396
rect 478874 12384 478880 12396
rect 478932 12384 478938 12436
rect 77386 11772 77392 11824
rect 77444 11812 77450 11824
rect 257338 11812 257344 11824
rect 77444 11784 257344 11812
rect 77444 11772 77450 11784
rect 257338 11772 257344 11784
rect 257396 11772 257402 11824
rect 98178 11704 98184 11756
rect 98236 11744 98242 11756
rect 298738 11744 298744 11756
rect 98236 11716 298744 11744
rect 98236 11704 98242 11716
rect 298738 11704 298744 11716
rect 298796 11704 298802 11756
rect 360838 10956 360844 11008
rect 360896 10996 360902 11008
rect 421558 10996 421564 11008
rect 360896 10968 421564 10996
rect 360896 10956 360902 10968
rect 421558 10956 421564 10968
rect 421616 10956 421622 11008
rect 258442 10888 258448 10940
rect 258500 10928 258506 10940
rect 259362 10928 259368 10940
rect 258500 10900 259368 10928
rect 258500 10888 258506 10900
rect 259362 10888 259368 10900
rect 259420 10888 259426 10940
rect 124674 10276 124680 10328
rect 124732 10316 124738 10328
rect 254578 10316 254584 10328
rect 124732 10288 254584 10316
rect 124732 10276 124738 10288
rect 254578 10276 254584 10288
rect 254636 10276 254642 10328
rect 259362 10276 259368 10328
rect 259420 10316 259426 10328
rect 486418 10316 486424 10328
rect 259420 10288 486424 10316
rect 259420 10276 259426 10288
rect 486418 10276 486424 10288
rect 486476 10276 486482 10328
rect 284938 9596 284944 9648
rect 284996 9636 285002 9648
rect 287790 9636 287796 9648
rect 284996 9608 287796 9636
rect 284996 9596 285002 9608
rect 287790 9596 287796 9608
rect 287848 9596 287854 9648
rect 305638 9596 305644 9648
rect 305696 9636 305702 9648
rect 374638 9636 374644 9648
rect 305696 9608 374644 9636
rect 305696 9596 305702 9608
rect 374638 9596 374644 9608
rect 374696 9596 374702 9648
rect 3418 8984 3424 9036
rect 3476 9024 3482 9036
rect 35158 9024 35164 9036
rect 3476 8996 35164 9024
rect 3476 8984 3482 8996
rect 35158 8984 35164 8996
rect 35216 8984 35222 9036
rect 62022 8984 62028 9036
rect 62080 9024 62086 9036
rect 282362 9024 282368 9036
rect 62080 8996 282368 9024
rect 62080 8984 62086 8996
rect 282362 8984 282368 8996
rect 282420 8984 282426 9036
rect 34790 8916 34796 8968
rect 34848 8956 34854 8968
rect 296070 8956 296076 8968
rect 34848 8928 296076 8956
rect 34848 8916 34854 8928
rect 296070 8916 296076 8928
rect 296128 8916 296134 8968
rect 339862 8916 339868 8968
rect 339920 8956 339926 8968
rect 423674 8956 423680 8968
rect 339920 8928 423680 8956
rect 339920 8916 339926 8928
rect 423674 8916 423680 8928
rect 423732 8916 423738 8968
rect 188338 7692 188344 7744
rect 188396 7732 188402 7744
rect 188396 7704 296714 7732
rect 188396 7692 188402 7704
rect 109310 7624 109316 7676
rect 109368 7664 109374 7676
rect 232498 7664 232504 7676
rect 109368 7636 232504 7664
rect 109368 7624 109374 7636
rect 232498 7624 232504 7636
rect 232556 7624 232562 7676
rect 1670 7556 1676 7608
rect 1728 7596 1734 7608
rect 43438 7596 43444 7608
rect 1728 7568 43444 7596
rect 1728 7556 1734 7568
rect 43438 7556 43444 7568
rect 43496 7556 43502 7608
rect 45462 7556 45468 7608
rect 45520 7596 45526 7608
rect 271138 7596 271144 7608
rect 45520 7568 271144 7596
rect 45520 7556 45526 7568
rect 271138 7556 271144 7568
rect 271196 7556 271202 7608
rect 296686 7596 296714 7704
rect 306742 7596 306748 7608
rect 296686 7568 306748 7596
rect 306742 7556 306748 7568
rect 306800 7596 306806 7608
rect 431954 7596 431960 7608
rect 306800 7568 431960 7596
rect 306800 7556 306806 7568
rect 431954 7556 431960 7568
rect 432012 7556 432018 7608
rect 282270 6808 282276 6860
rect 282328 6848 282334 6860
rect 439498 6848 439504 6860
rect 282328 6820 439504 6848
rect 282328 6808 282334 6820
rect 439498 6808 439504 6820
rect 439556 6808 439562 6860
rect 542998 6808 543004 6860
rect 543056 6848 543062 6860
rect 580166 6848 580172 6860
rect 543056 6820 580172 6848
rect 543056 6808 543062 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 308582 6740 308588 6792
rect 308640 6780 308646 6792
rect 309870 6780 309876 6792
rect 308640 6752 309876 6780
rect 308640 6740 308646 6752
rect 309870 6740 309876 6752
rect 309928 6740 309934 6792
rect 309962 6740 309968 6792
rect 310020 6780 310026 6792
rect 430574 6780 430580 6792
rect 310020 6752 430580 6780
rect 310020 6740 310026 6752
rect 430574 6740 430580 6752
rect 430632 6740 430638 6792
rect 79686 6196 79692 6248
rect 79744 6236 79750 6248
rect 301590 6236 301596 6248
rect 79744 6208 301596 6236
rect 79744 6196 79750 6208
rect 301590 6196 301596 6208
rect 301648 6196 301654 6248
rect 14734 6128 14740 6180
rect 14792 6168 14798 6180
rect 283650 6168 283656 6180
rect 14792 6140 283656 6168
rect 14792 6128 14798 6140
rect 283650 6128 283656 6140
rect 283708 6128 283714 6180
rect 257062 5448 257068 5500
rect 257120 5488 257126 5500
rect 257430 5488 257436 5500
rect 257120 5460 257436 5488
rect 257120 5448 257126 5460
rect 257430 5448 257436 5460
rect 257488 5488 257494 5500
rect 448514 5488 448520 5500
rect 257488 5460 448520 5488
rect 257488 5448 257494 5460
rect 448514 5448 448520 5460
rect 448572 5448 448578 5500
rect 43070 4836 43076 4888
rect 43128 4876 43134 4888
rect 291930 4876 291936 4888
rect 43128 4848 291936 4876
rect 43128 4836 43134 4848
rect 291930 4836 291936 4848
rect 291988 4836 291994 4888
rect 8754 4768 8760 4820
rect 8812 4808 8818 4820
rect 269758 4808 269764 4820
rect 8812 4780 269764 4808
rect 8812 4768 8818 4780
rect 269758 4768 269764 4780
rect 269816 4768 269822 4820
rect 293954 4768 293960 4820
rect 294012 4808 294018 4820
rect 294874 4808 294880 4820
rect 294012 4780 294880 4808
rect 294012 4768 294018 4780
rect 294874 4768 294880 4780
rect 294932 4808 294938 4820
rect 359458 4808 359464 4820
rect 294932 4780 359464 4808
rect 294932 4768 294938 4780
rect 359458 4768 359464 4780
rect 359516 4768 359522 4820
rect 197998 4088 198004 4140
rect 198056 4128 198062 4140
rect 246390 4128 246396 4140
rect 198056 4100 246396 4128
rect 198056 4088 198062 4100
rect 246390 4088 246396 4100
rect 246448 4088 246454 4140
rect 332686 4088 332692 4140
rect 332744 4128 332750 4140
rect 333238 4128 333244 4140
rect 332744 4100 333244 4128
rect 332744 4088 332750 4100
rect 333238 4088 333244 4100
rect 333296 4128 333302 4140
rect 342990 4128 342996 4140
rect 333296 4100 342996 4128
rect 333296 4088 333302 4100
rect 342990 4088 342996 4100
rect 343048 4088 343054 4140
rect 351178 4088 351184 4140
rect 351236 4128 351242 4140
rect 351638 4128 351644 4140
rect 351236 4100 351644 4128
rect 351236 4088 351242 4100
rect 351638 4088 351644 4100
rect 351696 4128 351702 4140
rect 373994 4128 374000 4140
rect 351696 4100 374000 4128
rect 351696 4088 351702 4100
rect 373994 4088 374000 4100
rect 374052 4088 374058 4140
rect 216030 4020 216036 4072
rect 216088 4060 216094 4072
rect 240502 4060 240508 4072
rect 216088 4032 240508 4060
rect 216088 4020 216094 4032
rect 240502 4020 240508 4032
rect 240560 4060 240566 4072
rect 240778 4060 240784 4072
rect 240560 4032 240784 4060
rect 240560 4020 240566 4032
rect 240778 4020 240784 4032
rect 240836 4020 240842 4072
rect 294598 4020 294604 4072
rect 294656 4060 294662 4072
rect 323302 4060 323308 4072
rect 294656 4032 323308 4060
rect 294656 4020 294662 4032
rect 323302 4020 323308 4032
rect 323360 4020 323366 4072
rect 331582 4020 331588 4072
rect 331640 4060 331646 4072
rect 339862 4060 339868 4072
rect 331640 4032 339868 4060
rect 331640 4020 331646 4032
rect 339862 4020 339868 4032
rect 339920 4020 339926 4072
rect 346946 4020 346952 4072
rect 347004 4060 347010 4072
rect 352650 4060 352656 4072
rect 347004 4032 352656 4060
rect 347004 4020 347010 4032
rect 352650 4020 352656 4032
rect 352708 4020 352714 4072
rect 274818 3952 274824 4004
rect 274876 3992 274882 4004
rect 275278 3992 275284 4004
rect 274876 3964 275284 3992
rect 274876 3952 274882 3964
rect 275278 3952 275284 3964
rect 275336 3992 275342 4004
rect 280798 3992 280804 4004
rect 275336 3964 280804 3992
rect 275336 3952 275342 3964
rect 280798 3952 280804 3964
rect 280856 3952 280862 4004
rect 309778 3952 309784 4004
rect 309836 3992 309842 4004
rect 320910 3992 320916 4004
rect 309836 3964 320916 3992
rect 309836 3952 309842 3964
rect 320910 3952 320916 3964
rect 320968 3952 320974 4004
rect 273898 3884 273904 3936
rect 273956 3924 273962 3936
rect 293954 3924 293960 3936
rect 273956 3896 293960 3924
rect 273956 3884 273962 3896
rect 293954 3884 293960 3896
rect 294012 3884 294018 3936
rect 308398 3884 308404 3936
rect 308456 3924 308462 3936
rect 319714 3924 319720 3936
rect 308456 3896 319720 3924
rect 308456 3884 308462 3896
rect 319714 3884 319720 3896
rect 319772 3884 319778 3936
rect 287698 3816 287704 3868
rect 287756 3856 287762 3868
rect 316218 3856 316224 3868
rect 287756 3828 316224 3856
rect 287756 3816 287762 3828
rect 316218 3816 316224 3828
rect 316276 3856 316282 3868
rect 316678 3856 316684 3868
rect 316276 3828 316684 3856
rect 316276 3816 316282 3828
rect 316678 3816 316684 3828
rect 316736 3816 316742 3868
rect 125870 3612 125876 3664
rect 125928 3652 125934 3664
rect 164878 3652 164884 3664
rect 125928 3624 164884 3652
rect 125928 3612 125934 3624
rect 164878 3612 164884 3624
rect 164936 3612 164942 3664
rect 251174 3612 251180 3664
rect 251232 3652 251238 3664
rect 252370 3652 252376 3664
rect 251232 3624 252376 3652
rect 251232 3612 251238 3624
rect 252370 3612 252376 3624
rect 252428 3612 252434 3664
rect 263594 3652 263600 3664
rect 258046 3624 263600 3652
rect 78582 3544 78588 3596
rect 78640 3584 78646 3596
rect 88978 3584 88984 3596
rect 78640 3556 88984 3584
rect 78640 3544 78646 3556
rect 88978 3544 88984 3556
rect 89036 3544 89042 3596
rect 93854 3544 93860 3596
rect 93912 3584 93918 3596
rect 94774 3584 94780 3596
rect 93912 3556 94780 3584
rect 93912 3544 93918 3556
rect 94774 3544 94780 3556
rect 94832 3544 94838 3596
rect 103330 3544 103336 3596
rect 103388 3584 103394 3596
rect 170398 3584 170404 3596
rect 103388 3556 170404 3584
rect 103388 3544 103394 3556
rect 170398 3544 170404 3556
rect 170456 3544 170462 3596
rect 242986 3584 242992 3596
rect 238726 3556 242992 3584
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 18598 3516 18604 3528
rect 6512 3488 18604 3516
rect 6512 3476 6518 3488
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 20254 3516 20260 3528
rect 19392 3488 20260 3516
rect 19392 3476 19398 3488
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 27614 3476 27620 3528
rect 27672 3516 27678 3528
rect 28534 3516 28540 3528
rect 27672 3488 28540 3516
rect 27672 3476 27678 3488
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 35894 3476 35900 3528
rect 35952 3516 35958 3528
rect 36814 3516 36820 3528
rect 35952 3488 36820 3516
rect 35952 3476 35958 3488
rect 36814 3476 36820 3488
rect 36872 3476 36878 3528
rect 69014 3476 69020 3528
rect 69072 3516 69078 3528
rect 69934 3516 69940 3528
rect 69072 3488 69940 3516
rect 69072 3476 69078 3488
rect 69934 3476 69940 3488
rect 69992 3476 69998 3528
rect 89162 3476 89168 3528
rect 89220 3516 89226 3528
rect 178770 3516 178776 3528
rect 89220 3488 178776 3516
rect 89220 3476 89226 3488
rect 178770 3476 178776 3488
rect 178828 3476 178834 3528
rect 217318 3476 217324 3528
rect 217376 3516 217382 3528
rect 238726 3516 238754 3556
rect 242986 3544 242992 3556
rect 243044 3584 243050 3596
rect 243044 3556 244228 3584
rect 243044 3544 243050 3556
rect 217376 3488 238754 3516
rect 217376 3476 217382 3488
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 244090 3516 244096 3528
rect 242952 3488 244096 3516
rect 242952 3476 242958 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 244200 3516 244228 3556
rect 247586 3544 247592 3596
rect 247644 3584 247650 3596
rect 258046 3584 258074 3624
rect 263594 3612 263600 3624
rect 263652 3612 263658 3664
rect 247644 3556 258074 3584
rect 247644 3544 247650 3556
rect 259454 3544 259460 3596
rect 259512 3584 259518 3596
rect 260650 3584 260656 3596
rect 259512 3556 260656 3584
rect 259512 3544 259518 3556
rect 260650 3544 260656 3556
rect 260708 3544 260714 3596
rect 271230 3584 271236 3596
rect 267706 3556 271236 3584
rect 267706 3516 267734 3556
rect 271230 3544 271236 3556
rect 271288 3544 271294 3596
rect 244200 3488 267734 3516
rect 276014 3476 276020 3528
rect 276072 3516 276078 3528
rect 276842 3516 276848 3528
rect 276072 3488 276848 3516
rect 276072 3476 276078 3488
rect 276842 3476 276848 3488
rect 276900 3476 276906 3528
rect 307754 3476 307760 3528
rect 307812 3516 307818 3528
rect 309042 3516 309048 3528
rect 307812 3488 309048 3516
rect 307812 3476 307818 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 316126 3476 316132 3528
rect 316184 3516 316190 3528
rect 317322 3516 317328 3528
rect 316184 3488 317328 3516
rect 316184 3476 316190 3488
rect 317322 3476 317328 3488
rect 317380 3476 317386 3528
rect 324958 3476 324964 3528
rect 325016 3516 325022 3528
rect 325602 3516 325608 3528
rect 325016 3488 325608 3516
rect 325016 3476 325022 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 329190 3476 329196 3528
rect 329248 3516 329254 3528
rect 331214 3516 331220 3528
rect 329248 3488 331220 3516
rect 329248 3476 329254 3488
rect 331214 3476 331220 3488
rect 331272 3476 331278 3528
rect 332594 3476 332600 3528
rect 332652 3516 332658 3528
rect 333882 3516 333888 3528
rect 332652 3488 333888 3516
rect 332652 3476 332658 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 340874 3476 340880 3528
rect 340932 3516 340938 3528
rect 342162 3516 342168 3528
rect 340932 3488 342168 3516
rect 340932 3476 340938 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 350442 3476 350448 3528
rect 350500 3516 350506 3528
rect 360838 3516 360844 3528
rect 350500 3488 360844 3516
rect 350500 3476 350506 3488
rect 360838 3476 360844 3488
rect 360896 3476 360902 3528
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 202230 3448 202236 3460
rect 18288 3420 202236 3448
rect 18288 3408 18294 3420
rect 202230 3408 202236 3420
rect 202288 3408 202294 3460
rect 215938 3408 215944 3460
rect 215996 3448 216002 3460
rect 239306 3448 239312 3460
rect 215996 3420 239312 3448
rect 215996 3408 216002 3420
rect 239306 3408 239312 3420
rect 239364 3448 239370 3460
rect 286410 3448 286416 3460
rect 239364 3420 286416 3448
rect 239364 3408 239370 3420
rect 286410 3408 286416 3420
rect 286468 3408 286474 3460
rect 313826 3408 313832 3460
rect 313884 3448 313890 3460
rect 318886 3448 318892 3460
rect 313884 3420 318892 3448
rect 313884 3408 313890 3420
rect 318886 3408 318892 3420
rect 318944 3408 318950 3460
rect 342070 3408 342076 3460
rect 342128 3448 342134 3460
rect 500954 3448 500960 3460
rect 342128 3420 500960 3448
rect 342128 3408 342134 3420
rect 500954 3408 500960 3420
rect 501012 3408 501018 3460
rect 135254 3340 135260 3392
rect 135312 3380 135318 3392
rect 136450 3380 136456 3392
rect 135312 3352 136456 3380
rect 135312 3340 135318 3352
rect 136450 3340 136456 3352
rect 136508 3340 136514 3392
rect 267734 3340 267740 3392
rect 267792 3380 267798 3392
rect 274634 3380 274640 3392
rect 267792 3352 274640 3380
rect 267792 3340 267798 3352
rect 274634 3340 274640 3352
rect 274692 3340 274698 3392
rect 282178 3272 282184 3324
rect 282236 3312 282242 3324
rect 285398 3312 285404 3324
rect 282236 3284 285404 3312
rect 282236 3272 282242 3284
rect 285398 3272 285404 3284
rect 285456 3272 285462 3324
rect 235810 3000 235816 3052
rect 235868 3040 235874 3052
rect 238018 3040 238024 3052
rect 235868 3012 238024 3040
rect 235868 3000 235874 3012
rect 238018 3000 238024 3012
rect 238076 3000 238082 3052
rect 41322 2184 41328 2236
rect 41380 2224 41386 2236
rect 129366 2224 129372 2236
rect 41380 2196 129372 2224
rect 41380 2184 41386 2196
rect 129366 2184 129372 2196
rect 129424 2184 129430 2236
rect 111610 2116 111616 2168
rect 111668 2156 111674 2168
rect 294782 2156 294788 2168
rect 111668 2128 294788 2156
rect 111668 2116 111674 2128
rect 294782 2116 294788 2128
rect 294840 2116 294846 2168
rect 64322 2048 64328 2100
rect 64380 2088 64386 2100
rect 294690 2088 294696 2100
rect 64380 2060 294696 2088
rect 64380 2048 64386 2060
rect 294690 2048 294696 2060
rect 294748 2048 294754 2100
<< via1 >>
rect 201500 703332 201552 703384
rect 202788 703332 202840 703384
rect 77944 703264 77996 703316
rect 267648 703264 267700 703316
rect 95148 703196 95200 703248
rect 332508 703196 332560 703248
rect 109684 703128 109736 703180
rect 348792 703128 348844 703180
rect 111064 703060 111116 703112
rect 397460 703060 397512 703112
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 76564 702992 76616 703044
rect 364984 702992 365036 703044
rect 104808 702924 104860 702976
rect 413652 702924 413704 702976
rect 115848 702856 115900 702908
rect 462320 702856 462372 702908
rect 75184 702788 75236 702840
rect 429200 702788 429252 702840
rect 429844 702788 429896 702840
rect 117228 702720 117280 702772
rect 478512 702720 478564 702772
rect 113088 702652 113140 702704
rect 453948 702652 454000 702704
rect 492588 702652 492640 702704
rect 494796 702652 494848 702704
rect 79324 702584 79376 702636
rect 527180 702584 527232 702636
rect 108948 702516 109000 702568
rect 511908 702516 511960 702568
rect 550548 702516 550600 702568
rect 559656 702516 559708 702568
rect 68928 702448 68980 702500
rect 543464 702448 543516 702500
rect 364984 701700 365036 701752
rect 483664 701700 483716 701752
rect 71044 700340 71096 700392
rect 154120 700340 154172 700392
rect 162124 700340 162176 700392
rect 218980 700340 219032 700392
rect 62028 700272 62080 700324
rect 235172 700272 235224 700324
rect 238024 700272 238076 700324
rect 283840 700272 283892 700324
rect 450544 700272 450596 700324
rect 453948 700272 454000 700324
rect 492588 700272 492640 700324
rect 511908 700272 511960 700324
rect 550548 700272 550600 700324
rect 511264 699660 511316 699712
rect 511908 699660 511960 699712
rect 24308 698912 24360 698964
rect 106280 698912 106332 698964
rect 57888 697552 57940 697604
rect 170312 697552 170364 697604
rect 69020 696940 69072 696992
rect 580172 696940 580224 696992
rect 159364 683136 159416 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 15844 670692 15896 670744
rect 90364 670692 90416 670744
rect 580908 670692 580960 670744
rect 3516 656888 3568 656940
rect 11704 656888 11756 656940
rect 3516 632068 3568 632120
rect 58624 632068 58676 632120
rect 119344 630640 119396 630692
rect 580172 630640 580224 630692
rect 3516 618264 3568 618316
rect 93124 618264 93176 618316
rect 425704 616088 425756 616140
rect 580172 616088 580224 616140
rect 6920 598204 6972 598256
rect 46848 598204 46900 598256
rect 46848 597524 46900 597576
rect 85580 597524 85632 597576
rect 68836 596776 68888 596828
rect 238024 596776 238076 596828
rect 3424 595416 3476 595468
rect 42800 595416 42852 595468
rect 42800 594804 42852 594856
rect 44088 594804 44140 594856
rect 71872 594804 71924 594856
rect 3516 594056 3568 594108
rect 106464 594056 106516 594108
rect 68652 592628 68704 592680
rect 136640 592628 136692 592680
rect 82084 591268 82136 591320
rect 90364 591268 90416 591320
rect 40040 590656 40092 590708
rect 48228 590656 48280 590708
rect 74632 590656 74684 590708
rect 556804 590656 556856 590708
rect 579804 590656 579856 590708
rect 11704 588548 11756 588600
rect 87328 588548 87380 588600
rect 88340 588548 88392 588600
rect 117412 588548 117464 588600
rect 103520 586712 103572 586764
rect 104808 586712 104860 586764
rect 131304 586712 131356 586764
rect 85304 586644 85356 586696
rect 113272 586644 113324 586696
rect 49608 586576 49660 586628
rect 79324 586576 79376 586628
rect 91008 586576 91060 586628
rect 123024 586576 123076 586628
rect 52368 586508 52420 586560
rect 84292 586508 84344 586560
rect 94872 586508 94924 586560
rect 128452 586508 128504 586560
rect 112076 585760 112128 585812
rect 162124 585760 162176 585812
rect 93124 585352 93176 585404
rect 95884 585352 95936 585404
rect 115940 585352 115992 585404
rect 61936 585284 61988 585336
rect 80612 585284 80664 585336
rect 95148 585284 95200 585336
rect 120080 585284 120132 585336
rect 50712 585216 50764 585268
rect 76564 585216 76616 585268
rect 87328 585216 87380 585268
rect 87512 585216 87564 585268
rect 118792 585216 118844 585268
rect 49516 585148 49568 585200
rect 78036 585148 78088 585200
rect 97908 585148 97960 585200
rect 131120 585148 131172 585200
rect 88248 584196 88300 584248
rect 105636 584196 105688 584248
rect 98736 584128 98788 584180
rect 101404 584128 101456 584180
rect 39856 583992 39908 584044
rect 77852 584060 77904 584112
rect 79232 584060 79284 584112
rect 99288 584060 99340 584112
rect 129832 584060 129884 584112
rect 66168 583992 66220 584044
rect 70952 583992 71004 584044
rect 96528 583992 96580 584044
rect 110420 583992 110472 584044
rect 56508 583924 56560 583976
rect 70400 583924 70452 583976
rect 101312 583924 101364 583976
rect 116032 583924 116084 583976
rect 41236 583856 41288 583908
rect 73344 583856 73396 583908
rect 101864 583856 101916 583908
rect 113364 583856 113416 583908
rect 59176 583788 59228 583840
rect 96712 583788 96764 583840
rect 104440 583788 104492 583840
rect 125692 583788 125744 583840
rect 70308 583720 70360 583772
rect 83372 583720 83424 583772
rect 88984 583720 89036 583772
rect 102140 583720 102192 583772
rect 105268 583720 105320 583772
rect 114560 583720 114612 583772
rect 60004 582972 60056 583024
rect 71780 582972 71832 583024
rect 102140 582972 102192 583024
rect 121460 582972 121512 583024
rect 92848 582632 92900 582684
rect 109040 582632 109092 582684
rect 83280 582564 83332 582616
rect 110512 582564 110564 582616
rect 54484 582496 54536 582548
rect 76748 582496 76800 582548
rect 91560 582496 91612 582548
rect 120172 582496 120224 582548
rect 57796 582428 57848 582480
rect 84476 582428 84528 582480
rect 89628 582428 89680 582480
rect 122840 582428 122892 582480
rect 14464 582360 14516 582412
rect 107660 582360 107712 582412
rect 68468 581952 68520 582004
rect 71044 581952 71096 582004
rect 65524 581748 65576 581800
rect 75460 581748 75512 581800
rect 72240 581680 72292 581732
rect 53104 581204 53156 581256
rect 67640 581204 67692 581256
rect 50804 581136 50856 581188
rect 48044 581068 48096 581120
rect 78680 581680 78732 581732
rect 90272 581680 90324 581732
rect 35808 581000 35860 581052
rect 65524 581000 65576 581052
rect 100576 581680 100628 581732
rect 104992 581680 105044 581732
rect 108948 581680 109000 581732
rect 117320 581136 117372 581188
rect 108948 581068 109000 581120
rect 127072 581068 127124 581120
rect 122932 581000 122984 581052
rect 65524 579640 65576 579692
rect 68652 579640 68704 579692
rect 108212 579640 108264 579692
rect 111800 579640 111852 579692
rect 64604 578280 64656 578332
rect 67732 578280 67784 578332
rect 108856 578280 108908 578332
rect 133144 578280 133196 578332
rect 53656 578212 53708 578264
rect 67640 578212 67692 578264
rect 108948 578212 109000 578264
rect 135260 578212 135312 578264
rect 69112 576988 69164 577040
rect 69756 576988 69808 577040
rect 64512 576852 64564 576904
rect 67640 576852 67692 576904
rect 105636 576104 105688 576156
rect 118884 576104 118936 576156
rect 37188 575492 37240 575544
rect 67640 575492 67692 575544
rect 108948 575492 109000 575544
rect 122748 575492 122800 575544
rect 431224 575492 431276 575544
rect 61752 574132 61804 574184
rect 67732 574132 67784 574184
rect 56324 574064 56376 574116
rect 67640 574064 67692 574116
rect 108948 574064 109000 574116
rect 137284 574064 137336 574116
rect 122104 573996 122156 574048
rect 159364 573996 159416 574048
rect 108948 573316 109000 573368
rect 122104 573316 122156 573368
rect 108672 572976 108724 573028
rect 113180 572976 113232 573028
rect 34428 572772 34480 572824
rect 67640 572772 67692 572824
rect 105636 572772 105688 572824
rect 110604 572772 110656 572824
rect 108948 572704 109000 572756
rect 128636 572704 128688 572756
rect 66076 571548 66128 571600
rect 68284 571548 68336 571600
rect 108948 571344 109000 571396
rect 140780 571344 140832 571396
rect 66168 571276 66220 571328
rect 68284 571276 68336 571328
rect 63224 569916 63276 569968
rect 67640 569916 67692 569968
rect 108948 569916 109000 569968
rect 142160 569916 142212 569968
rect 107660 568624 107712 568676
rect 109776 568624 109828 568676
rect 66168 568556 66220 568608
rect 67640 568556 67692 568608
rect 108948 567536 109000 567588
rect 114744 567536 114796 567588
rect 64696 567264 64748 567316
rect 67640 567264 67692 567316
rect 63316 567196 63368 567248
rect 67732 567196 67784 567248
rect 108948 567196 109000 567248
rect 117964 567196 118016 567248
rect 108856 565904 108908 565956
rect 125784 565904 125836 565956
rect 3240 565836 3292 565888
rect 25504 565836 25556 565888
rect 63132 565836 63184 565888
rect 67640 565836 67692 565888
rect 108948 565836 109000 565888
rect 142252 565836 142304 565888
rect 431224 565088 431276 565140
rect 497464 565088 497516 565140
rect 504364 565088 504416 565140
rect 57704 564408 57756 564460
rect 67640 564408 67692 564460
rect 108856 564408 108908 564460
rect 133880 564408 133932 564460
rect 204904 564408 204956 564460
rect 108948 564340 109000 564392
rect 117228 564340 117280 564392
rect 124312 564340 124364 564392
rect 504364 563660 504416 563712
rect 580172 563660 580224 563712
rect 60464 563116 60516 563168
rect 67640 563116 67692 563168
rect 52276 563048 52328 563100
rect 67732 563048 67784 563100
rect 60740 562300 60792 562352
rect 62028 562300 62080 562352
rect 67640 562300 67692 562352
rect 61844 561688 61896 561740
rect 67640 561688 67692 561740
rect 108948 561688 109000 561740
rect 130016 561688 130068 561740
rect 52184 560940 52236 560992
rect 60740 560940 60792 560992
rect 106924 560940 106976 560992
rect 116124 560940 116176 560992
rect 59268 560328 59320 560380
rect 67732 560328 67784 560380
rect 107660 560328 107712 560380
rect 138112 560328 138164 560380
rect 50988 560260 51040 560312
rect 67640 560260 67692 560312
rect 108948 560260 109000 560312
rect 139492 560260 139544 560312
rect 136824 559512 136876 559564
rect 201500 559512 201552 559564
rect 108948 558968 109000 559020
rect 124220 558968 124272 559020
rect 42708 558900 42760 558952
rect 67640 558900 67692 558952
rect 108856 558900 108908 558952
rect 136824 558900 136876 558952
rect 37096 558152 37148 558204
rect 68836 558152 68888 558204
rect 108948 557744 109000 557796
rect 114652 557744 114704 557796
rect 30288 557540 30340 557592
rect 67640 557540 67692 557592
rect 48136 556248 48188 556300
rect 67640 556248 67692 556300
rect 43904 556180 43956 556232
rect 67732 556180 67784 556232
rect 108948 556180 109000 556232
rect 127624 556180 127676 556232
rect 108856 556112 108908 556164
rect 110604 556112 110656 556164
rect 110604 555432 110656 555484
rect 119436 555432 119488 555484
rect 57980 554820 58032 554872
rect 67640 554820 67692 554872
rect 35716 554752 35768 554804
rect 67732 554752 67784 554804
rect 3516 554684 3568 554736
rect 14464 554684 14516 554736
rect 141516 554004 141568 554056
rect 556804 554004 556856 554056
rect 65616 553392 65668 553444
rect 67640 553392 67692 553444
rect 108948 553392 109000 553444
rect 140964 553392 141016 553444
rect 141516 553392 141568 553444
rect 55036 552032 55088 552084
rect 67640 552032 67692 552084
rect 108948 552032 109000 552084
rect 138020 552032 138072 552084
rect 107660 550672 107712 550724
rect 110696 550672 110748 550724
rect 46756 550604 46808 550656
rect 67640 550604 67692 550656
rect 108948 550604 109000 550656
rect 125600 550604 125652 550656
rect 108856 549312 108908 549364
rect 135444 549312 135496 549364
rect 41144 549244 41196 549296
rect 67640 549244 67692 549296
rect 108948 549244 109000 549296
rect 139584 549244 139636 549296
rect 64788 547952 64840 548004
rect 67640 547952 67692 548004
rect 56416 547884 56468 547936
rect 67732 547884 67784 547936
rect 61660 546524 61712 546576
rect 67732 546524 67784 546576
rect 60556 546456 60608 546508
rect 67640 546456 67692 546508
rect 108948 546456 109000 546508
rect 132592 546456 132644 546508
rect 108948 545708 109000 545760
rect 112352 545708 112404 545760
rect 33048 545096 33100 545148
rect 68100 545096 68152 545148
rect 108948 545096 109000 545148
rect 134248 545096 134300 545148
rect 25504 544348 25556 544400
rect 68008 544348 68060 544400
rect 108948 544348 109000 544400
rect 115848 544348 115900 544400
rect 116216 544348 116268 544400
rect 108948 543736 109000 543788
rect 140872 543736 140924 543788
rect 63408 542444 63460 542496
rect 67640 542444 67692 542496
rect 45468 542376 45520 542428
rect 68008 542376 68060 542428
rect 107844 542376 107896 542428
rect 134156 542376 134208 542428
rect 61936 541628 61988 541680
rect 69664 541628 69716 541680
rect 60648 540948 60700 541000
rect 67640 540948 67692 541000
rect 108304 540744 108356 540796
rect 109684 540744 109736 540796
rect 62028 539588 62080 539640
rect 67640 539588 67692 539640
rect 106832 539588 106884 539640
rect 142436 539588 142488 539640
rect 3424 539520 3476 539572
rect 98368 539520 98420 539572
rect 425060 539520 425112 539572
rect 425704 539520 425756 539572
rect 58624 539452 58676 539504
rect 99012 539452 99064 539504
rect 70308 539044 70360 539096
rect 71964 539044 72016 539096
rect 95148 538976 95200 539028
rect 109132 538976 109184 539028
rect 99288 538908 99340 538960
rect 121552 538908 121604 538960
rect 99012 538840 99064 538892
rect 129924 538840 129976 538892
rect 41328 538228 41380 538280
rect 60004 538228 60056 538280
rect 109684 538228 109736 538280
rect 123484 538228 123536 538280
rect 425060 538228 425112 538280
rect 73896 538160 73948 538212
rect 80336 538160 80388 538212
rect 111064 538160 111116 538212
rect 204904 538160 204956 538212
rect 580172 538160 580224 538212
rect 100944 538092 100996 538144
rect 119344 538092 119396 538144
rect 53748 537684 53800 537736
rect 82912 537684 82964 537736
rect 97080 537684 97132 537736
rect 102140 537684 102192 537736
rect 102232 537684 102284 537736
rect 110604 537684 110656 537736
rect 46664 537616 46716 537668
rect 79692 537616 79744 537668
rect 84108 537616 84160 537668
rect 89996 537616 90048 537668
rect 102876 537616 102928 537668
rect 128544 537616 128596 537668
rect 53196 537548 53248 537600
rect 86132 537548 86184 537600
rect 95792 537548 95844 537600
rect 121644 537548 121696 537600
rect 15844 537480 15896 537532
rect 57520 537480 57572 537532
rect 91284 537480 91336 537532
rect 100300 537480 100352 537532
rect 132684 537480 132736 537532
rect 83464 536800 83516 536852
rect 85488 536800 85540 536852
rect 94504 536800 94556 536852
rect 117412 536732 117464 536784
rect 101956 536664 102008 536716
rect 105544 536664 105596 536716
rect 38476 536052 38528 536104
rect 71320 536052 71372 536104
rect 117412 535440 117464 535492
rect 118700 535440 118752 535492
rect 57796 534964 57848 535016
rect 75184 534964 75236 535016
rect 52000 534896 52052 534948
rect 78404 534896 78456 534948
rect 50896 534828 50948 534880
rect 83556 534828 83608 534880
rect 45284 534760 45336 534812
rect 77760 534760 77812 534812
rect 91008 534760 91060 534812
rect 115940 534760 115992 534812
rect 39948 534692 40000 534744
rect 73252 534692 73304 534744
rect 93860 534692 93912 534744
rect 128360 534692 128412 534744
rect 420920 534692 420972 534744
rect 429200 534692 429252 534744
rect 52368 533332 52420 533384
rect 69296 533332 69348 533384
rect 69756 533332 69808 533384
rect 72424 533264 72476 533316
rect 52092 532176 52144 532228
rect 72608 532176 72660 532228
rect 55128 532108 55180 532160
rect 76472 532108 76524 532160
rect 45376 532040 45428 532092
rect 75092 532040 75144 532092
rect 84844 532040 84896 532092
rect 111984 532040 112036 532092
rect 39672 531972 39724 532024
rect 71872 531972 71924 532024
rect 93768 531972 93820 532024
rect 123024 531972 123076 532024
rect 41052 529252 41104 529304
rect 70400 529252 70452 529304
rect 42524 529184 42576 529236
rect 77116 529184 77168 529236
rect 110696 529184 110748 529236
rect 116676 529184 116728 529236
rect 3148 528504 3200 528556
rect 110696 528572 110748 528624
rect 69204 525716 69256 525768
rect 579804 525716 579856 525768
rect 2780 514768 2832 514820
rect 4804 514768 4856 514820
rect 431224 510620 431276 510672
rect 580172 510620 580224 510672
rect 87420 499468 87472 499520
rect 114836 499536 114888 499588
rect 131212 499536 131264 499588
rect 89352 498856 89404 498908
rect 113548 498856 113600 498908
rect 69664 498788 69716 498840
rect 74540 498788 74592 498840
rect 80612 498788 80664 498840
rect 88064 498788 88116 498840
rect 128452 498788 128504 498840
rect 4804 498108 4856 498160
rect 59176 498108 59228 498160
rect 59176 497632 59228 497684
rect 91100 497632 91152 497684
rect 93216 497632 93268 497684
rect 117504 497632 117556 497684
rect 85580 497564 85632 497616
rect 120172 497564 120224 497616
rect 126980 497564 127032 497616
rect 84108 497496 84160 497548
rect 120264 497496 120316 497548
rect 83280 497428 83332 497480
rect 122932 497428 122984 497480
rect 131396 497428 131448 497480
rect 53656 496748 53708 496800
rect 58072 496748 58124 496800
rect 430580 496748 430632 496800
rect 53656 496272 53708 496324
rect 83464 496272 83516 496324
rect 81532 496204 81584 496256
rect 116124 496204 116176 496256
rect 430580 496204 430632 496256
rect 431224 496204 431276 496256
rect 79692 496136 79744 496188
rect 113272 496136 113324 496188
rect 116584 496136 116636 496188
rect 49424 496068 49476 496120
rect 80980 496068 81032 496120
rect 95056 496068 95108 496120
rect 131120 496068 131172 496120
rect 141056 496068 141108 496120
rect 78404 495456 78456 495508
rect 112076 495456 112128 495508
rect 116124 495456 116176 495508
rect 121552 495456 121604 495508
rect 3424 495388 3476 495440
rect 83280 495388 83332 495440
rect 75184 494980 75236 495032
rect 78404 494980 78456 495032
rect 94964 494980 95016 495032
rect 111892 494980 111944 495032
rect 114836 494980 114888 495032
rect 98644 494912 98696 494964
rect 120356 494912 120408 494964
rect 94872 494844 94924 494896
rect 116032 494844 116084 494896
rect 132500 494844 132552 494896
rect 80980 494776 81032 494828
rect 118792 494776 118844 494828
rect 125876 494776 125928 494828
rect 82912 494708 82964 494760
rect 122840 494708 122892 494760
rect 130108 494708 130160 494760
rect 92480 494028 92532 494080
rect 93768 494028 93820 494080
rect 110696 494028 110748 494080
rect 91928 493824 91980 493876
rect 95056 493824 95108 493876
rect 95792 493484 95844 493536
rect 90272 493416 90324 493468
rect 110420 493416 110472 493468
rect 113364 493416 113416 493468
rect 127164 493416 127216 493468
rect 54116 493348 54168 493400
rect 54944 493348 54996 493400
rect 74816 493348 74868 493400
rect 88708 493348 88760 493400
rect 120080 493348 120132 493400
rect 122840 493348 122892 493400
rect 43996 493280 44048 493332
rect 49516 493280 49568 493332
rect 71688 493280 71740 493332
rect 93216 493280 93268 493332
rect 129832 493280 129884 493332
rect 139400 493280 139452 493332
rect 75828 493008 75880 493060
rect 81532 493008 81584 493060
rect 81624 492804 81676 492856
rect 96528 492804 96580 492856
rect 46572 492736 46624 492788
rect 53840 492736 53892 492788
rect 57888 492736 57940 492788
rect 90272 492736 90324 492788
rect 39856 492668 39908 492720
rect 70952 492668 71004 492720
rect 77760 492668 77812 492720
rect 120080 492668 120132 492720
rect 72424 492600 72476 492652
rect 84844 492600 84896 492652
rect 92480 492600 92532 492652
rect 97724 492600 97776 492652
rect 99288 492600 99340 492652
rect 53840 492124 53892 492176
rect 54484 492124 54536 492176
rect 70400 492124 70452 492176
rect 50712 492056 50764 492108
rect 70032 492056 70084 492108
rect 86132 492056 86184 492108
rect 87144 492056 87196 492108
rect 89904 492056 89956 492108
rect 92020 492056 92072 492108
rect 102416 492056 102468 492108
rect 114468 492056 114520 492108
rect 125692 492056 125744 492108
rect 39764 491988 39816 492040
rect 48044 491988 48096 492040
rect 72240 491988 72292 492040
rect 76472 491988 76524 492040
rect 110512 491988 110564 492040
rect 123024 491988 123076 492040
rect 56140 491920 56192 491972
rect 90640 491920 90692 491972
rect 97080 491920 97132 491972
rect 131304 491920 131356 491972
rect 143540 491920 143592 491972
rect 89996 491784 90048 491836
rect 91008 491784 91060 491836
rect 92572 491648 92624 491700
rect 94964 491648 95016 491700
rect 95148 491648 95200 491700
rect 96344 491648 96396 491700
rect 91008 491512 91060 491564
rect 99932 491512 99984 491564
rect 71780 491444 71832 491496
rect 76748 491444 76800 491496
rect 86776 491444 86828 491496
rect 96436 491444 96488 491496
rect 99012 491444 99064 491496
rect 110420 491444 110472 491496
rect 54852 491376 54904 491428
rect 65616 491376 65668 491428
rect 65984 491376 66036 491428
rect 98368 491376 98420 491428
rect 113456 491376 113508 491428
rect 114468 491376 114520 491428
rect 80060 491308 80112 491360
rect 93860 491308 93912 491360
rect 99288 491308 99340 491360
rect 99656 491308 99708 491360
rect 114560 491308 114612 491360
rect 46848 491240 46900 491292
rect 48964 491240 49016 491292
rect 96528 491240 96580 491292
rect 115112 491240 115164 491292
rect 118884 491240 118936 491292
rect 110420 491172 110472 491224
rect 111708 491172 111760 491224
rect 127072 491172 127124 491224
rect 89904 490696 89956 490748
rect 99380 490696 99432 490748
rect 58992 490628 59044 490680
rect 79048 490628 79100 490680
rect 96252 490628 96304 490680
rect 113364 490628 113416 490680
rect 42616 490560 42668 490612
rect 49608 490560 49660 490612
rect 73252 490560 73304 490612
rect 86868 490560 86920 490612
rect 109132 490560 109184 490612
rect 104900 489880 104952 489932
rect 35808 489812 35860 489864
rect 67640 489812 67692 489864
rect 91560 489812 91612 489864
rect 102048 489812 102100 489864
rect 109040 489812 109092 489864
rect 109316 489812 109368 489864
rect 118792 489812 118844 489864
rect 121460 489812 121512 489864
rect 103428 489132 103480 489184
rect 117412 489132 117464 489184
rect 121460 489132 121512 489184
rect 579620 489132 579672 489184
rect 34336 488520 34388 488572
rect 35808 488520 35860 488572
rect 103428 488452 103480 488504
rect 111800 488452 111852 488504
rect 109040 488384 109092 488436
rect 110328 488384 110380 488436
rect 117320 488384 117372 488436
rect 111800 487840 111852 487892
rect 128452 487840 128504 487892
rect 48228 487772 48280 487824
rect 57796 487772 57848 487824
rect 103428 487772 103480 487824
rect 133144 487772 133196 487824
rect 136732 487772 136784 487824
rect 114560 487500 114612 487552
rect 118792 487500 118844 487552
rect 57612 487160 57664 487212
rect 57796 487160 57848 487212
rect 67640 487160 67692 487212
rect 103428 487092 103480 487144
rect 135260 487092 135312 487144
rect 136548 487092 136600 487144
rect 136548 486480 136600 486532
rect 150532 486480 150584 486532
rect 41236 486412 41288 486464
rect 67640 486412 67692 486464
rect 103428 486412 103480 486464
rect 106188 486412 106240 486464
rect 135352 486412 135404 486464
rect 50804 485732 50856 485784
rect 65616 485800 65668 485852
rect 67640 485800 67692 485852
rect 102140 485052 102192 485104
rect 111800 485052 111852 485104
rect 112628 485052 112680 485104
rect 67272 484576 67324 484628
rect 68652 484576 68704 484628
rect 44088 484304 44140 484356
rect 47584 484440 47636 484492
rect 67640 484440 67692 484492
rect 99656 484372 99708 484424
rect 112536 484372 112588 484424
rect 112628 484372 112680 484424
rect 121460 484372 121512 484424
rect 56232 484304 56284 484356
rect 56508 484304 56560 484356
rect 99932 484304 99984 484356
rect 103520 484304 103572 484356
rect 56232 483624 56284 483676
rect 67640 483624 67692 483676
rect 102140 483624 102192 483676
rect 122932 483624 122984 483676
rect 37004 483012 37056 483064
rect 137284 483012 137336 483064
rect 147956 483012 148008 483064
rect 53104 482944 53156 482996
rect 67640 482944 67692 482996
rect 102140 482944 102192 482996
rect 48044 481652 48096 481704
rect 65524 481652 65576 481704
rect 65984 481652 66036 481704
rect 102140 481652 102192 481704
rect 117044 481652 117096 481704
rect 64604 481584 64656 481636
rect 68008 481584 68060 481636
rect 102324 481584 102376 481636
rect 128636 481584 128688 481636
rect 65984 481516 66036 481568
rect 67640 481516 67692 481568
rect 102140 480904 102192 480956
rect 113180 480904 113232 480956
rect 128636 480904 128688 480956
rect 146300 480904 146352 480956
rect 59176 480156 59228 480208
rect 67640 480156 67692 480208
rect 102140 480156 102192 480208
rect 140780 480156 140832 480208
rect 102140 479680 102192 479732
rect 104992 479680 105044 479732
rect 106188 479680 106240 479732
rect 112536 479476 112588 479528
rect 117320 479476 117372 479528
rect 140780 479476 140832 479528
rect 145012 479476 145064 479528
rect 109776 478864 109828 478916
rect 136640 478864 136692 478916
rect 63040 477572 63092 477624
rect 63224 477572 63276 477624
rect 102140 477504 102192 477556
rect 115848 477504 115900 477556
rect 61752 477436 61804 477488
rect 63224 477436 63276 477488
rect 67732 477436 67784 477488
rect 102324 477436 102376 477488
rect 114744 477436 114796 477488
rect 116032 477436 116084 477488
rect 102140 477368 102192 477420
rect 109776 477368 109828 477420
rect 106188 476756 106240 476808
rect 151820 476756 151872 476808
rect 35808 476076 35860 476128
rect 67640 476076 67692 476128
rect 117964 476076 118016 476128
rect 120172 476076 120224 476128
rect 102416 476008 102468 476060
rect 103428 476008 103480 476060
rect 142160 476008 142212 476060
rect 102324 475940 102376 475992
rect 125784 475940 125836 475992
rect 131764 475940 131816 475992
rect 102140 475872 102192 475924
rect 117964 475872 118016 475924
rect 55956 475328 56008 475380
rect 56324 475328 56376 475380
rect 67640 475328 67692 475380
rect 105636 474852 105688 474904
rect 107936 474852 107988 474904
rect 3424 474716 3476 474768
rect 25504 474716 25556 474768
rect 34428 474648 34480 474700
rect 64236 474648 64288 474700
rect 67640 474716 67692 474768
rect 102140 474648 102192 474700
rect 142252 474648 142304 474700
rect 150624 474648 150676 474700
rect 66076 473288 66128 473340
rect 67640 473288 67692 473340
rect 102324 473288 102376 473340
rect 106372 473288 106424 473340
rect 107568 473288 107620 473340
rect 99564 472744 99616 472796
rect 110604 472744 110656 472796
rect 107568 472676 107620 472728
rect 118884 472676 118936 472728
rect 48228 472608 48280 472660
rect 66076 472608 66128 472660
rect 102140 472608 102192 472660
rect 133880 472608 133932 472660
rect 102140 471928 102192 471980
rect 124312 471928 124364 471980
rect 129740 471928 129792 471980
rect 64972 471588 65024 471640
rect 67640 471588 67692 471640
rect 118884 471316 118936 471368
rect 146392 471316 146444 471368
rect 50804 471248 50856 471300
rect 63040 471248 63092 471300
rect 67640 471248 67692 471300
rect 102876 471248 102928 471300
rect 139492 471248 139544 471300
rect 59084 470568 59136 470620
rect 64972 470568 65024 470620
rect 102324 470568 102376 470620
rect 107568 470568 107620 470620
rect 112628 470568 112680 470620
rect 139492 470568 139544 470620
rect 142344 470568 142396 470620
rect 146392 470568 146444 470620
rect 579896 470568 579948 470620
rect 102140 470500 102192 470552
rect 130016 470500 130068 470552
rect 130016 469888 130068 469940
rect 152004 469888 152056 469940
rect 103612 469820 103664 469872
rect 138112 469820 138164 469872
rect 142252 469820 142304 469872
rect 64512 469480 64564 469532
rect 66168 469480 66220 469532
rect 67732 469480 67784 469532
rect 43812 469208 43864 469260
rect 66076 469208 66128 469260
rect 67640 469208 67692 469260
rect 64696 469072 64748 469124
rect 66076 469072 66128 469124
rect 66076 468188 66128 468240
rect 67640 468188 67692 468240
rect 60372 467848 60424 467900
rect 63316 467848 63368 467900
rect 67732 467848 67784 467900
rect 61752 466760 61804 466812
rect 63132 466760 63184 466812
rect 67640 466760 67692 466812
rect 102140 466488 102192 466540
rect 115204 466488 115256 466540
rect 115848 466488 115900 466540
rect 103152 466420 103204 466472
rect 102140 466352 102192 466404
rect 119988 466352 120040 466404
rect 136824 466352 136876 466404
rect 115848 466284 115900 466336
rect 124220 466284 124272 466336
rect 114652 466216 114704 466268
rect 121736 466216 121788 466268
rect 102140 465672 102192 465724
rect 103336 465672 103388 465724
rect 107752 465672 107804 465724
rect 57704 464992 57756 465044
rect 65524 465060 65576 465112
rect 67732 465060 67784 465112
rect 127624 465060 127676 465112
rect 138112 465060 138164 465112
rect 102140 464992 102192 465044
rect 101404 464924 101456 464976
rect 102232 464924 102284 464976
rect 108488 464380 108540 464432
rect 111984 464380 112036 464432
rect 427820 464312 427872 464364
rect 497464 464312 497516 464364
rect 102140 464108 102192 464160
rect 105636 464108 105688 464160
rect 60464 463768 60516 463820
rect 64144 463768 64196 463820
rect 67640 463768 67692 463820
rect 52276 463632 52328 463684
rect 53104 463632 53156 463684
rect 67824 463700 67876 463752
rect 60464 463632 60516 463684
rect 61844 463632 61896 463684
rect 67732 463632 67784 463684
rect 102140 463632 102192 463684
rect 119436 463632 119488 463684
rect 124220 463700 124272 463752
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 52276 462272 52328 462324
rect 53196 462272 53248 462324
rect 59176 462272 59228 462324
rect 67640 462340 67692 462392
rect 107568 462340 107620 462392
rect 140964 462340 141016 462392
rect 102232 462272 102284 462324
rect 124404 462272 124456 462324
rect 125968 462272 126020 462324
rect 59268 462204 59320 462256
rect 63224 462204 63276 462256
rect 102140 462204 102192 462256
rect 107568 462204 107620 462256
rect 52184 461592 52236 461644
rect 59176 461592 59228 461644
rect 63224 460912 63276 460964
rect 67640 460912 67692 460964
rect 102140 460844 102192 460896
rect 107016 460912 107068 460964
rect 147864 460912 147916 460964
rect 50988 460232 51040 460284
rect 67640 460232 67692 460284
rect 42708 460164 42760 460216
rect 67732 460164 67784 460216
rect 50712 459552 50764 459604
rect 50988 459552 51040 459604
rect 102232 459552 102284 459604
rect 107476 459552 107528 459604
rect 116676 459552 116728 459604
rect 133972 459552 134024 459604
rect 138020 459484 138072 459536
rect 102140 459416 102192 459468
rect 116676 459416 116728 459468
rect 35164 458872 35216 458924
rect 42708 458872 42760 458924
rect 37096 458804 37148 458856
rect 67456 458804 67508 458856
rect 67640 458804 67692 458856
rect 107568 458804 107620 458856
rect 135444 458804 135496 458856
rect 30288 458124 30340 458176
rect 33784 458260 33836 458312
rect 67640 458260 67692 458312
rect 135444 458192 135496 458244
rect 139492 458192 139544 458244
rect 43720 458124 43772 458176
rect 48136 458124 48188 458176
rect 67732 458124 67784 458176
rect 103244 458124 103296 458176
rect 125600 458124 125652 458176
rect 102140 458056 102192 458108
rect 107568 458056 107620 458108
rect 43904 457444 43956 457496
rect 44088 457444 44140 457496
rect 67640 457444 67692 457496
rect 431960 457444 432012 457496
rect 579620 457444 579672 457496
rect 106188 456764 106240 456816
rect 151912 456764 151964 456816
rect 42432 456696 42484 456748
rect 44088 456696 44140 456748
rect 102140 456696 102192 456748
rect 139584 456696 139636 456748
rect 140320 456696 140372 456748
rect 102232 456628 102284 456680
rect 105544 456628 105596 456680
rect 106188 456628 106240 456680
rect 35716 456016 35768 456068
rect 67640 456016 67692 456068
rect 140320 456016 140372 456068
rect 149152 456016 149204 456068
rect 105544 455948 105596 456000
rect 109132 455948 109184 456000
rect 56508 455812 56560 455864
rect 57980 455812 58032 455864
rect 35716 455336 35768 455388
rect 36636 455336 36688 455388
rect 57980 455336 58032 455388
rect 67640 455336 67692 455388
rect 102140 455336 102192 455388
rect 132592 455404 132644 455456
rect 107660 455336 107712 455388
rect 108304 455336 108356 455388
rect 102140 454792 102192 454844
rect 107660 454792 107712 454844
rect 100668 454724 100720 454776
rect 113180 454724 113232 454776
rect 106188 454656 106240 454708
rect 134248 454656 134300 454708
rect 143724 454656 143776 454708
rect 46848 453976 46900 454028
rect 54852 453976 54904 454028
rect 67640 453976 67692 454028
rect 54484 453296 54536 453348
rect 55036 453296 55088 453348
rect 67640 453296 67692 453348
rect 102876 453296 102928 453348
rect 125600 453296 125652 453348
rect 102140 453228 102192 453280
rect 106188 453228 106240 453280
rect 102140 452548 102192 452600
rect 116216 452548 116268 452600
rect 124864 452548 124916 452600
rect 103612 451868 103664 451920
rect 134156 451868 134208 451920
rect 147772 451868 147824 451920
rect 103704 451664 103756 451716
rect 107844 451664 107896 451716
rect 69204 451256 69256 451308
rect 46756 451188 46808 451240
rect 62764 451188 62816 451240
rect 41144 449828 41196 449880
rect 61384 449896 61436 449948
rect 67640 449896 67692 449948
rect 106924 449896 106976 449948
rect 140780 449896 140832 449948
rect 102140 449828 102192 449880
rect 56416 449148 56468 449200
rect 67640 449148 67692 449200
rect 106188 449148 106240 449200
rect 142436 449148 142488 449200
rect 143816 449148 143868 449200
rect 3148 448536 3200 448588
rect 50344 448536 50396 448588
rect 55864 448536 55916 448588
rect 56416 448536 56468 448588
rect 102232 448468 102284 448520
rect 107476 448468 107528 448520
rect 102140 448400 102192 448452
rect 106188 448400 106240 448452
rect 107476 448060 107528 448112
rect 113456 448060 113508 448112
rect 61660 447176 61712 447228
rect 66260 447176 66312 447228
rect 67640 447176 67692 447228
rect 64788 447108 64840 447160
rect 66168 447108 66220 447160
rect 67732 447108 67784 447160
rect 33048 446360 33100 446412
rect 67640 446360 67692 446412
rect 104164 445816 104216 445868
rect 108396 445816 108448 445868
rect 60556 445748 60608 445800
rect 64604 445748 64656 445800
rect 67732 445748 67784 445800
rect 101956 445748 102008 445800
rect 138204 445748 138256 445800
rect 103152 445068 103204 445120
rect 104164 445068 104216 445120
rect 102600 445000 102652 445052
rect 128544 445000 128596 445052
rect 142160 445000 142212 445052
rect 99472 444388 99524 444440
rect 100760 444388 100812 444440
rect 45468 443640 45520 443692
rect 67640 443640 67692 443692
rect 61936 442892 61988 442944
rect 63408 442892 63460 442944
rect 67640 442892 67692 442944
rect 38568 442212 38620 442264
rect 67640 442212 67692 442264
rect 102692 441668 102744 441720
rect 112536 441668 112588 441720
rect 103152 441600 103204 441652
rect 132868 441600 132920 441652
rect 60648 441532 60700 441584
rect 67640 441532 67692 441584
rect 62028 440988 62080 441040
rect 67640 440988 67692 441040
rect 52092 440920 52144 440972
rect 45284 440852 45336 440904
rect 112076 440920 112128 440972
rect 72148 440648 72200 440700
rect 72332 440648 72384 440700
rect 92388 440648 92440 440700
rect 94136 440648 94188 440700
rect 117504 440852 117556 440904
rect 103152 440308 103204 440360
rect 127072 440308 127124 440360
rect 132684 440308 132736 440360
rect 102140 440240 102192 440292
rect 133880 440240 133932 440292
rect 67272 439560 67324 439612
rect 75184 439560 75236 439612
rect 89812 439560 89864 439612
rect 113548 439560 113600 439612
rect 53656 439492 53708 439544
rect 83464 439492 83516 439544
rect 85764 439492 85816 439544
rect 96528 439492 96580 439544
rect 120264 439492 120316 439544
rect 56140 439016 56192 439068
rect 59268 439016 59320 439068
rect 90916 439016 90968 439068
rect 88708 438948 88760 439000
rect 123484 438948 123536 439000
rect 123760 438948 123812 439000
rect 25504 438880 25556 438932
rect 96436 438880 96488 438932
rect 4804 438812 4856 438864
rect 50896 438812 50948 438864
rect 89996 438812 90048 438864
rect 95884 438812 95936 438864
rect 96528 438812 96580 438864
rect 99656 438812 99708 438864
rect 122932 438880 122984 438932
rect 129924 438880 129976 438932
rect 46664 438744 46716 438796
rect 78772 438744 78824 438796
rect 96436 438744 96488 438796
rect 121644 438744 121696 438796
rect 52184 438676 52236 438728
rect 53748 438676 53800 438728
rect 82912 438676 82964 438728
rect 99012 438676 99064 438728
rect 120356 438676 120408 438728
rect 120908 438676 120960 438728
rect 87604 438608 87656 438660
rect 105544 438608 105596 438660
rect 97080 438540 97132 438592
rect 113364 438540 113416 438592
rect 114468 438540 114520 438592
rect 50344 438472 50396 438524
rect 99472 438472 99524 438524
rect 53104 438268 53156 438320
rect 73896 438268 73948 438320
rect 88064 438268 88116 438320
rect 88984 438268 89036 438320
rect 121644 438268 121696 438320
rect 125784 438268 125836 438320
rect 44272 438200 44324 438252
rect 71320 438200 71372 438252
rect 50896 438132 50948 438184
rect 52092 438132 52144 438184
rect 83556 438200 83608 438252
rect 92572 438200 92624 438252
rect 97908 438200 97960 438252
rect 101404 438200 101456 438252
rect 120908 438200 120960 438252
rect 129924 438200 129976 438252
rect 75460 438132 75512 438184
rect 82268 438132 82320 438184
rect 84844 438132 84896 438184
rect 97724 438132 97776 438184
rect 114468 438132 114520 438184
rect 135260 438132 135312 438184
rect 78772 437860 78824 437912
rect 79692 437860 79744 437912
rect 81624 437452 81676 437504
rect 82820 437452 82872 437504
rect 38476 437384 38528 437436
rect 44272 437384 44324 437436
rect 44824 437384 44876 437436
rect 52276 437384 52328 437436
rect 86224 437384 86276 437436
rect 86776 437384 86828 437436
rect 94504 437384 94556 437436
rect 128360 437384 128412 437436
rect 49424 437316 49476 437368
rect 81624 437316 81676 437368
rect 95148 437316 95200 437368
rect 118700 437316 118752 437368
rect 39672 437248 39724 437300
rect 71964 437248 72016 437300
rect 72148 437248 72200 437300
rect 77300 437248 77352 437300
rect 77760 437248 77812 437300
rect 41328 437180 41380 437232
rect 53104 437180 53156 437232
rect 58992 437180 59044 437232
rect 78864 437180 78916 437232
rect 79048 437180 79100 437232
rect 65616 436704 65668 436756
rect 76564 436704 76616 436756
rect 97724 436704 97776 436756
rect 107384 436704 107436 436756
rect 108488 436704 108540 436756
rect 57520 436024 57572 436076
rect 91744 436024 91796 436076
rect 45376 435956 45428 436008
rect 74632 435956 74684 436008
rect 75828 435956 75880 436008
rect 42524 435412 42576 435464
rect 44088 435412 44140 435464
rect 77116 435412 77168 435464
rect 40684 435344 40736 435396
rect 73252 435344 73304 435396
rect 39948 434664 40000 434716
rect 40684 434664 40736 434716
rect 52000 434664 52052 434716
rect 69020 434664 69072 434716
rect 78588 434664 78640 434716
rect 82912 434664 82964 434716
rect 38476 433236 38528 433288
rect 41052 433236 41104 433288
rect 70676 433236 70728 433288
rect 55128 433168 55180 433220
rect 76472 433168 76524 433220
rect 82912 431876 82964 431928
rect 579804 431876 579856 431928
rect 101496 431808 101548 431860
rect 140872 431808 140924 431860
rect 140872 431196 140924 431248
rect 150716 431196 150768 431248
rect 3424 429836 3476 429888
rect 101496 429836 101548 429888
rect 69204 428408 69256 428460
rect 579620 428408 579672 428460
rect 3516 422288 3568 422340
rect 118792 422220 118844 422272
rect 118792 420928 118844 420980
rect 119344 420928 119396 420980
rect 525064 418752 525116 418804
rect 579620 418752 579672 418804
rect 579988 418752 580040 418804
rect 87696 404336 87748 404388
rect 579620 404336 579672 404388
rect 104256 403656 104308 403708
rect 128636 403656 128688 403708
rect 96620 403588 96672 403640
rect 127256 403588 127308 403640
rect 61844 402976 61896 403028
rect 289084 402976 289136 403028
rect 93768 402228 93820 402280
rect 130016 402228 130068 402280
rect 70400 401616 70452 401668
rect 71044 401616 71096 401668
rect 358820 401616 358872 401668
rect 104164 401004 104216 401056
rect 132776 401004 132828 401056
rect 86224 400936 86276 400988
rect 123116 400936 123168 400988
rect 93676 400868 93728 400920
rect 131304 400868 131356 400920
rect 50804 400120 50856 400172
rect 69112 400188 69164 400240
rect 357440 400188 357492 400240
rect 107568 399508 107620 399560
rect 117504 399508 117556 399560
rect 91744 399440 91796 399492
rect 124312 399440 124364 399492
rect 94136 398896 94188 398948
rect 115112 398896 115164 398948
rect 50988 398828 51040 398880
rect 107016 398828 107068 398880
rect 114836 398828 114888 398880
rect 160744 398828 160796 398880
rect 108396 398216 108448 398268
rect 136824 398216 136876 398268
rect 56232 398148 56284 398200
rect 71044 398148 71096 398200
rect 108304 398148 108356 398200
rect 140872 398148 140924 398200
rect 3148 398080 3200 398132
rect 116032 398080 116084 398132
rect 98644 397536 98696 397588
rect 188344 397536 188396 397588
rect 67364 397468 67416 397520
rect 202144 397468 202196 397520
rect 95884 396856 95936 396908
rect 120724 396856 120776 396908
rect 69664 396788 69716 396840
rect 94504 396788 94556 396840
rect 101128 396788 101180 396840
rect 131212 396788 131264 396840
rect 46756 396720 46808 396772
rect 77300 396720 77352 396772
rect 95148 396720 95200 396772
rect 125692 396720 125744 396772
rect 178684 396720 178736 396772
rect 72424 396040 72476 396092
rect 146944 396040 146996 396092
rect 116584 395972 116636 396024
rect 120264 395972 120316 396024
rect 46572 395360 46624 395412
rect 81808 395360 81860 395412
rect 110604 395360 110656 395412
rect 127164 395360 127216 395412
rect 42616 395292 42668 395344
rect 84844 395292 84896 395344
rect 88340 395292 88392 395344
rect 123024 395292 123076 395344
rect 170404 395292 170456 395344
rect 39580 394816 39632 394868
rect 110604 394816 110656 394868
rect 81808 394748 81860 394800
rect 154580 394748 154632 394800
rect 84844 394680 84896 394732
rect 85120 394680 85172 394732
rect 195244 394680 195296 394732
rect 77852 394136 77904 394188
rect 87696 394136 87748 394188
rect 105636 394136 105688 394188
rect 117596 394136 117648 394188
rect 57704 394068 57756 394120
rect 83464 394068 83516 394120
rect 103336 394068 103388 394120
rect 116124 394068 116176 394120
rect 47952 394000 48004 394052
rect 78772 394000 78824 394052
rect 99288 394000 99340 394052
rect 135444 394000 135496 394052
rect 39856 393932 39908 393984
rect 83004 393932 83056 393984
rect 98552 393932 98604 393984
rect 126980 393932 127032 393984
rect 196624 393932 196676 393984
rect 83004 393388 83056 393440
rect 150440 393388 150492 393440
rect 53656 393252 53708 393304
rect 147680 393320 147732 393372
rect 60648 392640 60700 392692
rect 89812 392640 89864 392692
rect 97448 392640 97500 392692
rect 131396 392640 131448 392692
rect 139584 392640 139636 392692
rect 43996 392572 44048 392624
rect 82912 392572 82964 392624
rect 88248 392572 88300 392624
rect 121552 392572 121604 392624
rect 186964 392572 187016 392624
rect 91560 392096 91612 392148
rect 92388 392096 92440 392148
rect 121552 392096 121604 392148
rect 82912 392028 82964 392080
rect 83648 392028 83700 392080
rect 138020 392028 138072 392080
rect 51724 391960 51776 392012
rect 121644 391892 121696 391944
rect 109408 391620 109460 391672
rect 110696 391620 110748 391672
rect 39764 391280 39816 391332
rect 52460 391280 52512 391332
rect 57612 391280 57664 391332
rect 78220 391280 78272 391332
rect 112536 391280 112588 391332
rect 131212 391280 131264 391332
rect 47584 391212 47636 391264
rect 75552 391212 75604 391264
rect 110696 391212 110748 391264
rect 228364 391212 228416 391264
rect 52460 390736 52512 390788
rect 53196 390736 53248 390788
rect 84476 390736 84528 390788
rect 111708 390736 111760 390788
rect 114928 390736 114980 390788
rect 34336 390668 34388 390720
rect 36544 390668 36596 390720
rect 80060 390668 80112 390720
rect 94044 390668 94096 390720
rect 123484 390668 123536 390720
rect 125876 390668 125928 390720
rect 78220 390600 78272 390652
rect 126980 390600 127032 390652
rect 75552 390532 75604 390584
rect 137284 390532 137336 390584
rect 107476 390464 107528 390516
rect 114284 390464 114336 390516
rect 103244 389852 103296 389904
rect 115296 389852 115348 389904
rect 130384 389852 130436 389904
rect 139400 389852 139452 389904
rect 49516 389784 49568 389836
rect 82820 389784 82872 389836
rect 96528 389784 96580 389836
rect 130108 389784 130160 389836
rect 142436 389784 142488 389836
rect 57796 389308 57848 389360
rect 104532 389308 104584 389360
rect 114284 389308 114336 389360
rect 118792 389308 118844 389360
rect 119344 389308 119396 389360
rect 128544 389308 128596 389360
rect 57244 389240 57296 389292
rect 57612 389240 57664 389292
rect 79324 389240 79376 389292
rect 101036 389240 101088 389292
rect 102048 389240 102100 389292
rect 128360 389240 128412 389292
rect 102600 389172 102652 389224
rect 136916 389172 136968 389224
rect 198096 389172 198148 389224
rect 37096 389104 37148 389156
rect 71044 389104 71096 389156
rect 74816 389104 74868 389156
rect 115756 389104 115808 389156
rect 119344 389104 119396 389156
rect 72424 389036 72476 389088
rect 98460 388628 98512 388680
rect 109408 388628 109460 388680
rect 97908 388560 97960 388612
rect 111800 388560 111852 388612
rect 91008 388492 91060 388544
rect 120080 388492 120132 388544
rect 122012 388492 122064 388544
rect 4804 388424 4856 388476
rect 37096 388424 37148 388476
rect 41144 388424 41196 388476
rect 48044 388424 48096 388476
rect 71780 388424 71832 388476
rect 86408 388424 86460 388476
rect 98644 388424 98696 388476
rect 106924 388424 106976 388476
rect 141056 388424 141108 388476
rect 204904 388424 204956 388476
rect 74908 388084 74960 388136
rect 184204 388084 184256 388136
rect 112168 388016 112220 388068
rect 112444 388016 112496 388068
rect 119344 388016 119396 388068
rect 58532 387948 58584 388000
rect 87052 387948 87104 388000
rect 48964 387880 49016 387932
rect 52368 387880 52420 387932
rect 92940 387880 92992 387932
rect 109592 387880 109644 387932
rect 110328 387880 110380 387932
rect 200764 387880 200816 387932
rect 54944 387812 54996 387864
rect 55128 387812 55180 387864
rect 69756 387812 69808 387864
rect 92848 387812 92900 387864
rect 108948 387812 109000 387864
rect 115848 387812 115900 387864
rect 120264 387744 120316 387796
rect 56416 387200 56468 387252
rect 71964 387200 72016 387252
rect 70124 387132 70176 387184
rect 87604 387132 87656 387184
rect 107384 387132 107436 387184
rect 124404 387132 124456 387184
rect 48044 387064 48096 387116
rect 74632 387064 74684 387116
rect 88984 387064 89036 387116
rect 118700 387064 118752 387116
rect 50896 386520 50948 386572
rect 80612 386520 80664 386572
rect 103888 386520 103940 386572
rect 122104 386520 122156 386572
rect 39764 386452 39816 386504
rect 103796 386452 103848 386504
rect 103980 386452 104032 386504
rect 110328 386452 110380 386504
rect 132500 386452 132552 386504
rect 74816 386384 74868 386436
rect 286324 386384 286376 386436
rect 104900 386316 104952 386368
rect 105912 386316 105964 386368
rect 41236 385772 41288 385824
rect 50804 385772 50856 385824
rect 46664 385704 46716 385756
rect 78864 385704 78916 385756
rect 112720 385704 112772 385756
rect 117412 385704 117464 385756
rect 43996 385636 44048 385688
rect 100668 385636 100720 385688
rect 120264 385636 120316 385688
rect 50804 385024 50856 385076
rect 77484 385296 77536 385348
rect 90272 385296 90324 385348
rect 100024 385296 100076 385348
rect 106280 385296 106332 385348
rect 120080 385160 120132 385212
rect 287704 385092 287756 385144
rect 308404 385024 308456 385076
rect 115940 384956 115992 385008
rect 128452 384956 128504 385008
rect 63132 383732 63184 383784
rect 65892 383732 65944 383784
rect 34428 383664 34480 383716
rect 68744 383664 68796 383716
rect 118516 383664 118568 383716
rect 360844 383664 360896 383716
rect 118608 383596 118660 383648
rect 136732 383596 136784 383648
rect 136732 382916 136784 382968
rect 145104 382916 145156 382968
rect 41328 382236 41380 382288
rect 67640 382236 67692 382288
rect 118608 381488 118660 381540
rect 135352 381488 135404 381540
rect 49608 380808 49660 380860
rect 67640 380808 67692 380860
rect 118608 380808 118660 380860
rect 121460 380808 121512 380860
rect 122196 380808 122248 380860
rect 48136 380264 48188 380316
rect 49608 380264 49660 380316
rect 118332 380128 118384 380180
rect 295984 380128 296036 380180
rect 64236 379516 64288 379568
rect 65984 379516 66036 379568
rect 67640 379516 67692 379568
rect 118608 378836 118660 378888
rect 122840 378836 122892 378888
rect 123024 378836 123076 378888
rect 119344 378768 119396 378820
rect 276664 378768 276716 378820
rect 519544 378768 519596 378820
rect 579620 378768 579672 378820
rect 118608 378156 118660 378208
rect 122196 378156 122248 378208
rect 147956 378088 148008 378140
rect 48228 377408 48280 377460
rect 67640 377408 67692 377460
rect 147956 377408 148008 377460
rect 441620 377408 441672 377460
rect 118424 376728 118476 376780
rect 143632 376728 143684 376780
rect 118608 376660 118660 376712
rect 146300 376660 146352 376712
rect 149060 376660 149112 376712
rect 117780 376252 117832 376304
rect 120264 376252 120316 376304
rect 42616 375368 42668 375420
rect 48228 375368 48280 375420
rect 43812 375300 43864 375352
rect 69112 375300 69164 375352
rect 118608 375300 118660 375352
rect 145012 375300 145064 375352
rect 146208 375300 146260 375352
rect 64512 374620 64564 374672
rect 64788 374620 64840 374672
rect 67640 374620 67692 374672
rect 60372 373940 60424 373992
rect 65892 373940 65944 373992
rect 118608 373940 118660 373992
rect 151820 373940 151872 373992
rect 3240 372512 3292 372564
rect 51724 372512 51776 372564
rect 61844 372512 61896 372564
rect 67640 372512 67692 372564
rect 66076 371900 66128 371952
rect 67732 371900 67784 371952
rect 60556 371832 60608 371884
rect 69664 371832 69716 371884
rect 117872 370472 117924 370524
rect 136732 370472 136784 370524
rect 65524 370132 65576 370184
rect 68376 370132 68428 370184
rect 116032 369860 116084 369912
rect 116216 369860 116268 369912
rect 118056 369860 118108 369912
rect 151820 369860 151872 369912
rect 53656 369792 53708 369844
rect 67640 369792 67692 369844
rect 117320 369112 117372 369164
rect 120172 369112 120224 369164
rect 131120 369112 131172 369164
rect 117412 368568 117464 368620
rect 117688 368568 117740 368620
rect 131396 368500 131448 368552
rect 131764 368500 131816 368552
rect 146300 368500 146352 368552
rect 117412 368432 117464 368484
rect 150624 368432 150676 368484
rect 151176 368432 151228 368484
rect 117320 368364 117372 368416
rect 131396 368364 131448 368416
rect 60372 367752 60424 367804
rect 69756 367752 69808 367804
rect 151176 367684 151228 367736
rect 152096 367684 152148 367736
rect 60464 367004 60516 367056
rect 68008 367004 68060 367056
rect 117320 367004 117372 367056
rect 134064 367004 134116 367056
rect 136640 367004 136692 367056
rect 59176 366324 59228 366376
rect 67640 366324 67692 366376
rect 136732 366324 136784 366376
rect 579620 366324 579672 366376
rect 63224 365644 63276 365696
rect 64696 365644 64748 365696
rect 119068 365644 119120 365696
rect 129740 365644 129792 365696
rect 34336 365576 34388 365628
rect 35164 365576 35216 365628
rect 119896 365032 119948 365084
rect 146392 365032 146444 365084
rect 122104 364964 122156 365016
rect 305644 364964 305696 365016
rect 117320 364828 117372 364880
rect 119896 364828 119948 364880
rect 64696 364352 64748 364404
rect 67640 364352 67692 364404
rect 50712 364284 50764 364336
rect 67732 364284 67784 364336
rect 34336 363604 34388 363656
rect 67640 363604 67692 363656
rect 117688 363604 117740 363656
rect 307024 363604 307076 363656
rect 48228 362992 48280 363044
rect 50712 362992 50764 363044
rect 42432 362924 42484 362976
rect 59084 362924 59136 362976
rect 117320 362856 117372 362908
rect 152004 362856 152056 362908
rect 153108 362856 153160 362908
rect 35716 362176 35768 362228
rect 42432 362176 42484 362228
rect 117320 362176 117372 362228
rect 121368 362176 121420 362228
rect 142344 362176 142396 362228
rect 153108 362176 153160 362228
rect 191104 362176 191156 362228
rect 59084 361496 59136 361548
rect 67640 361496 67692 361548
rect 141792 361496 141844 361548
rect 142252 361496 142304 361548
rect 118884 360272 118936 360324
rect 119988 360272 120040 360324
rect 134064 360272 134116 360324
rect 117320 360204 117372 360256
rect 141424 360204 141476 360256
rect 141792 360204 141844 360256
rect 43720 359456 43772 359508
rect 59084 359456 59136 359508
rect 59084 358776 59136 358828
rect 67640 358776 67692 358828
rect 117872 358776 117924 358828
rect 206284 358776 206336 358828
rect 36636 358028 36688 358080
rect 53840 358028 53892 358080
rect 56508 358028 56560 358080
rect 67640 358028 67692 358080
rect 118608 358028 118660 358080
rect 121644 358028 121696 358080
rect 143540 358028 143592 358080
rect 3148 357416 3200 357468
rect 43444 357416 43496 357468
rect 53840 357416 53892 357468
rect 54944 357416 54996 357468
rect 67732 357416 67784 357468
rect 131396 356668 131448 356720
rect 138112 356668 138164 356720
rect 118608 356124 118660 356176
rect 131396 356124 131448 356176
rect 131764 356124 131816 356176
rect 52276 356056 52328 356108
rect 60004 356056 60056 356108
rect 54484 355988 54536 356040
rect 118148 356056 118200 356108
rect 308496 356056 308548 356108
rect 46848 355920 46900 355972
rect 60004 355920 60056 355972
rect 67640 355988 67692 356040
rect 67732 355920 67784 355972
rect 118608 355308 118660 355360
rect 280804 355308 280856 355360
rect 118516 354628 118568 354680
rect 140964 354628 141016 354680
rect 118608 354016 118660 354068
rect 124220 354016 124272 354068
rect 119344 353948 119396 354000
rect 580356 353948 580408 354000
rect 62764 353268 62816 353320
rect 67364 353268 67416 353320
rect 67640 353268 67692 353320
rect 124220 353268 124272 353320
rect 125600 353268 125652 353320
rect 140964 353268 141016 353320
rect 142252 353268 142304 353320
rect 61384 352588 61436 352640
rect 67640 352588 67692 352640
rect 42800 352520 42852 352572
rect 43904 352520 43956 352572
rect 68928 352520 68980 352572
rect 118608 352520 118660 352572
rect 124220 352520 124272 352572
rect 125968 352520 126020 352572
rect 504364 352520 504416 352572
rect 579620 352520 579672 352572
rect 7564 351908 7616 351960
rect 42800 351908 42852 351960
rect 61384 351908 61436 351960
rect 61844 351908 61896 351960
rect 118056 351840 118108 351892
rect 147864 351840 147916 351892
rect 118608 351228 118660 351280
rect 158720 351228 158772 351280
rect 63316 351160 63368 351212
rect 67916 351160 67968 351212
rect 147864 351160 147916 351212
rect 213184 351160 213236 351212
rect 46848 350548 46900 350600
rect 55864 350480 55916 350532
rect 67640 350480 67692 350532
rect 118608 349800 118660 349852
rect 133972 349800 134024 349852
rect 66168 349732 66220 349784
rect 68376 349732 68428 349784
rect 63316 349120 63368 349172
rect 66260 349120 66312 349172
rect 67640 349052 67692 349104
rect 118608 349052 118660 349104
rect 139492 349052 139544 349104
rect 139768 349052 139820 349104
rect 139768 348372 139820 348424
rect 180064 348372 180116 348424
rect 57888 347760 57940 347812
rect 117872 347760 117924 347812
rect 297364 347760 297416 347812
rect 67732 347692 67784 347744
rect 117412 347692 117464 347744
rect 149152 347692 149204 347744
rect 149704 347692 149756 347744
rect 149704 347080 149756 347132
rect 215944 347080 215996 347132
rect 64604 347012 64656 347064
rect 67640 347012 67692 347064
rect 158720 347012 158772 347064
rect 347044 347012 347096 347064
rect 43444 346332 43496 346384
rect 68192 346332 68244 346384
rect 118608 346332 118660 346384
rect 132592 346332 132644 346384
rect 133788 346332 133840 346384
rect 2780 346264 2832 346316
rect 4804 346264 4856 346316
rect 118516 345652 118568 345704
rect 122104 345652 122156 345704
rect 151912 345720 151964 345772
rect 133788 345652 133840 345704
rect 209044 345652 209096 345704
rect 53656 345040 53708 345092
rect 68652 345040 68704 345092
rect 118608 344972 118660 345024
rect 140872 344972 140924 345024
rect 45468 344292 45520 344344
rect 49424 344292 49476 344344
rect 140872 344292 140924 344344
rect 305736 344292 305788 344344
rect 49424 343612 49476 343664
rect 67640 343612 67692 343664
rect 117780 343544 117832 343596
rect 143724 343544 143776 343596
rect 144828 343544 144880 343596
rect 118608 342864 118660 342916
rect 126152 342864 126204 342916
rect 144828 342864 144880 342916
rect 278044 342864 278096 342916
rect 126152 342320 126204 342372
rect 128452 342320 128504 342372
rect 61936 342252 61988 342304
rect 67272 342252 67324 342304
rect 67640 342252 67692 342304
rect 118608 342184 118660 342236
rect 124864 342184 124916 342236
rect 140872 342252 140924 342304
rect 115756 341572 115808 341624
rect 128636 341572 128688 341624
rect 38568 341504 38620 341556
rect 68652 341504 68704 341556
rect 124864 341504 124916 341556
rect 133972 341504 134024 341556
rect 485044 341504 485096 341556
rect 117504 340212 117556 340264
rect 150716 340212 150768 340264
rect 62028 340144 62080 340196
rect 67916 340144 67968 340196
rect 118424 340144 118476 340196
rect 147772 340144 147824 340196
rect 377404 340144 377456 340196
rect 70400 339940 70452 339992
rect 71044 339940 71096 339992
rect 56416 339532 56468 339584
rect 73252 339532 73304 339584
rect 107936 339532 107988 339584
rect 131212 339532 131264 339584
rect 47952 339464 48004 339516
rect 81624 339464 81676 339516
rect 113272 339464 113324 339516
rect 113824 339464 113876 339516
rect 143816 339464 143868 339516
rect 52092 339396 52144 339448
rect 86224 339396 86276 339448
rect 107384 339396 107436 339448
rect 107568 339396 107620 339448
rect 132868 339396 132920 339448
rect 40684 339328 40736 339380
rect 73896 339328 73948 339380
rect 53748 339260 53800 339312
rect 86776 339260 86828 339312
rect 60372 339192 60424 339244
rect 89996 339192 90048 339244
rect 90364 339192 90416 339244
rect 113088 338920 113140 338972
rect 118792 338920 118844 338972
rect 70308 338852 70360 338904
rect 98644 338852 98696 338904
rect 112444 338852 112496 338904
rect 122196 338852 122248 338904
rect 70492 338784 70544 338836
rect 309784 338784 309836 338836
rect 97908 338716 97960 338768
rect 124404 338716 124456 338768
rect 506480 338716 506532 338768
rect 580264 338716 580316 338768
rect 38476 338036 38528 338088
rect 70676 338104 70728 338156
rect 70032 338036 70084 338088
rect 71780 338036 71832 338088
rect 87420 338036 87472 338088
rect 96712 338036 96764 338088
rect 97908 338036 97960 338088
rect 102140 338036 102192 338088
rect 109960 338036 110012 338088
rect 112536 338036 112588 338088
rect 138112 338036 138164 338088
rect 48044 337968 48096 338020
rect 76472 337968 76524 338020
rect 86776 337968 86828 338020
rect 87604 337968 87656 338020
rect 115112 337968 115164 338020
rect 140780 337968 140832 338020
rect 44824 337900 44876 337952
rect 71320 337900 71372 337952
rect 100300 337900 100352 337952
rect 125784 337900 125836 337952
rect 126888 337900 126940 337952
rect 53104 337832 53156 337884
rect 74540 337832 74592 337884
rect 75184 337832 75236 337884
rect 95792 337832 95844 337884
rect 120172 337832 120224 337884
rect 76564 337696 76616 337748
rect 78404 337696 78456 337748
rect 91284 337696 91336 337748
rect 93676 337696 93728 337748
rect 73252 337560 73304 337612
rect 91008 337560 91060 337612
rect 70676 337492 70728 337544
rect 93308 337492 93360 337544
rect 126888 337492 126940 337544
rect 140780 337492 140832 337544
rect 58992 337424 59044 337476
rect 84200 337424 84252 337476
rect 99656 337424 99708 337476
rect 102048 337424 102100 337476
rect 125692 337424 125744 337476
rect 138112 337424 138164 337476
rect 177304 337424 177356 337476
rect 81624 337356 81676 337408
rect 211804 337356 211856 337408
rect 97080 337016 97132 337068
rect 100024 337016 100076 337068
rect 71320 336880 71372 336932
rect 76656 336880 76708 336932
rect 120172 336744 120224 336796
rect 320824 336744 320876 336796
rect 49516 336676 49568 336728
rect 52184 336608 52236 336660
rect 53748 336608 53800 336660
rect 39672 336540 39724 336592
rect 46756 336472 46808 336524
rect 79140 336608 79192 336660
rect 79324 336676 79376 336728
rect 79692 336676 79744 336728
rect 106096 336676 106148 336728
rect 127072 336676 127124 336728
rect 83464 336608 83516 336660
rect 104164 336608 104216 336660
rect 104808 336608 104860 336660
rect 122932 336608 122984 336660
rect 71964 336540 72016 336592
rect 57704 336472 57756 336524
rect 88984 336472 89036 336524
rect 56324 336404 56376 336456
rect 79324 336404 79376 336456
rect 53748 335996 53800 336048
rect 84844 335996 84896 336048
rect 60556 335248 60608 335300
rect 98368 335248 98420 335300
rect 103520 335248 103572 335300
rect 129924 335248 129976 335300
rect 42708 335180 42760 335232
rect 75828 335180 75880 335232
rect 93676 335180 93728 335232
rect 118700 335180 118752 335232
rect 44088 335112 44140 335164
rect 76564 335112 76616 335164
rect 59268 334704 59320 334756
rect 62028 334704 62080 334756
rect 94504 334704 94556 334756
rect 59176 334636 59228 334688
rect 134616 334636 134668 334688
rect 71780 334568 71832 334620
rect 291844 334568 291896 334620
rect 75276 334092 75328 334144
rect 75828 334092 75880 334144
rect 56416 333956 56468 334008
rect 60556 333956 60608 334008
rect 129740 333956 129792 334008
rect 129924 333956 129976 334008
rect 46664 333888 46716 333940
rect 80704 333888 80756 333940
rect 95056 333888 95108 333940
rect 124312 333888 124364 333940
rect 60648 333820 60700 333872
rect 92572 333820 92624 333872
rect 61844 333276 61896 333328
rect 162124 333276 162176 333328
rect 71964 333208 72016 333260
rect 309140 333208 309192 333260
rect 92572 332596 92624 332648
rect 93124 332596 93176 332648
rect 113916 332528 113968 332580
rect 144920 332528 144972 332580
rect 146208 332528 146260 332580
rect 113180 332052 113232 332104
rect 113916 332052 113968 332104
rect 55036 331984 55088 332036
rect 82268 331984 82320 332036
rect 95148 331984 95200 332036
rect 113272 331984 113324 332036
rect 76472 331916 76524 331968
rect 116584 331916 116636 331968
rect 54944 331848 54996 331900
rect 117964 331848 118016 331900
rect 146208 331848 146260 331900
rect 499580 331848 499632 331900
rect 67364 330488 67416 330540
rect 77300 330488 77352 330540
rect 120172 329808 120224 329860
rect 120724 329808 120776 329860
rect 125784 329808 125836 329860
rect 100944 329740 100996 329792
rect 135260 329740 135312 329792
rect 136548 329740 136600 329792
rect 93216 329672 93268 329724
rect 120172 329672 120224 329724
rect 93768 329060 93820 329112
rect 115112 329060 115164 329112
rect 136548 329060 136600 329112
rect 282184 329060 282236 329112
rect 89352 328380 89404 328432
rect 123116 328380 123168 328432
rect 124128 328380 124180 328432
rect 97724 328312 97776 328364
rect 130016 328312 130068 328364
rect 130384 328312 130436 328364
rect 124128 327768 124180 327820
rect 242164 327768 242216 327820
rect 130384 327700 130436 327752
rect 284944 327700 284996 327752
rect 110604 327020 110656 327072
rect 136824 327020 136876 327072
rect 137100 327020 137152 327072
rect 65984 326340 66036 326392
rect 115296 326340 115348 326392
rect 72424 325660 72476 325712
rect 108304 325660 108356 325712
rect 111248 325592 111300 325644
rect 132684 325592 132736 325644
rect 133788 325592 133840 325644
rect 106188 325048 106240 325100
rect 115940 325048 115992 325100
rect 80704 324980 80756 325032
rect 198004 324980 198056 325032
rect 48044 324912 48096 324964
rect 107660 324912 107712 324964
rect 133788 324912 133840 324964
rect 340144 324912 340196 324964
rect 14464 324300 14516 324352
rect 48044 324300 48096 324352
rect 67456 323688 67508 323740
rect 121460 323688 121512 323740
rect 93308 323620 93360 323672
rect 265624 323620 265676 323672
rect 76656 323552 76708 323604
rect 345664 323552 345716 323604
rect 86224 322260 86276 322312
rect 147772 322260 147824 322312
rect 88984 322192 89036 322244
rect 217324 322192 217376 322244
rect 105452 321512 105504 321564
rect 133880 321512 133932 321564
rect 135168 321512 135220 321564
rect 67272 320900 67324 320952
rect 207664 320900 207716 320952
rect 65984 320832 66036 320884
rect 112444 320832 112496 320884
rect 135168 320832 135220 320884
rect 349804 320832 349856 320884
rect 100024 320084 100076 320136
rect 131304 320084 131356 320136
rect 131672 320084 131724 320136
rect 75184 319472 75236 319524
rect 115388 319472 115440 319524
rect 69204 319404 69256 319456
rect 121644 319404 121696 319456
rect 106096 318112 106148 318164
rect 113824 318112 113876 318164
rect 83464 318044 83516 318096
rect 351920 318044 351972 318096
rect 60004 316752 60056 316804
rect 128636 316752 128688 316804
rect 84292 316684 84344 316736
rect 113916 316684 113968 316736
rect 115204 316684 115256 316736
rect 204996 316684 205048 316736
rect 91928 315936 91980 315988
rect 124404 315936 124456 315988
rect 73160 315256 73212 315308
rect 116032 315256 116084 315308
rect 69112 313896 69164 313948
rect 282276 313896 282328 313948
rect 69020 313284 69072 313336
rect 122564 313284 122616 313336
rect 395344 313284 395396 313336
rect 102232 313216 102284 313268
rect 127256 313216 127308 313268
rect 71136 312536 71188 312588
rect 129832 312536 129884 312588
rect 410524 312536 410576 312588
rect 81440 311856 81492 311908
rect 356060 311856 356112 311908
rect 102876 311788 102928 311840
rect 135444 311788 135496 311840
rect 136548 311788 136600 311840
rect 117964 311720 118016 311772
rect 125508 311720 125560 311772
rect 79324 311312 79376 311364
rect 120172 311312 120224 311364
rect 91100 311244 91152 311296
rect 121552 311244 121604 311296
rect 159364 311244 159416 311296
rect 70308 311176 70360 311228
rect 104164 311176 104216 311228
rect 136548 311176 136600 311228
rect 273904 311176 273956 311228
rect 114468 311108 114520 311160
rect 141424 311108 141476 311160
rect 464344 311108 464396 311160
rect 539508 311108 539560 311160
rect 580172 311108 580224 311160
rect 124312 310496 124364 310548
rect 125508 310496 125560 310548
rect 538220 310496 538272 310548
rect 539508 310496 539560 310548
rect 3424 310428 3476 310480
rect 48136 310428 48188 310480
rect 80060 309884 80112 309936
rect 91100 309884 91152 309936
rect 107660 309884 107712 309936
rect 134524 309884 134576 309936
rect 135168 309884 135220 309936
rect 76564 309816 76616 309868
rect 192484 309816 192536 309868
rect 48136 309748 48188 309800
rect 116676 309748 116728 309800
rect 135168 309748 135220 309800
rect 521660 309748 521712 309800
rect 75184 309204 75236 309256
rect 228456 309204 228508 309256
rect 89720 309136 89772 309188
rect 304264 309136 304316 309188
rect 108304 309068 108356 309120
rect 142160 309068 142212 309120
rect 143448 309068 143500 309120
rect 75920 308456 75972 308508
rect 216036 308456 216088 308508
rect 84384 308388 84436 308440
rect 114468 308388 114520 308440
rect 143448 308388 143500 308440
rect 475384 308388 475436 308440
rect 102048 307776 102100 307828
rect 103704 307776 103756 307828
rect 467104 307776 467156 307828
rect 93676 307028 93728 307080
rect 279424 307028 279476 307080
rect 86960 306484 87012 306536
rect 213276 306484 213328 306536
rect 85580 306416 85632 306468
rect 240784 306416 240836 306468
rect 106280 306348 106332 306400
rect 118884 306348 118936 306400
rect 514760 306348 514812 306400
rect 3424 306212 3476 306264
rect 7564 306212 7616 306264
rect 59084 305736 59136 305788
rect 123668 305736 123720 305788
rect 90364 305668 90416 305720
rect 275284 305668 275336 305720
rect 93124 305600 93176 305652
rect 294604 305600 294656 305652
rect 81900 305056 81952 305108
rect 221464 305056 221516 305108
rect 49424 304920 49476 304972
rect 77392 304920 77444 304972
rect 367744 304988 367796 305040
rect 107568 304308 107620 304360
rect 127624 304308 127676 304360
rect 60648 304240 60700 304292
rect 124864 304240 124916 304292
rect 146944 303900 146996 303952
rect 196716 303900 196768 303952
rect 233884 303832 233936 303884
rect 94504 303764 94556 303816
rect 95056 303764 95108 303816
rect 96620 303764 96672 303816
rect 315304 303764 315356 303816
rect 86316 303696 86368 303748
rect 318064 303696 318116 303748
rect 56508 303560 56560 303612
rect 66904 303560 66956 303612
rect 482284 303628 482336 303680
rect 93952 302880 94004 302932
rect 122840 302880 122892 302932
rect 90272 302472 90324 302524
rect 135904 302472 135956 302524
rect 66168 302404 66220 302456
rect 169024 302404 169076 302456
rect 115940 302336 115992 302388
rect 116676 302336 116728 302388
rect 232596 302336 232648 302388
rect 75920 302268 75972 302320
rect 193864 302268 193916 302320
rect 71780 302200 71832 302252
rect 325700 302200 325752 302252
rect 105636 301520 105688 301572
rect 43904 301452 43956 301504
rect 124404 301452 124456 301504
rect 145104 301452 145156 301504
rect 238024 301452 238076 301504
rect 104900 301384 104952 301436
rect 106188 301384 106240 301436
rect 106188 301044 106240 301096
rect 187056 301044 187108 301096
rect 79324 300976 79376 301028
rect 214656 300976 214708 301028
rect 88340 300908 88392 300960
rect 347780 300908 347832 300960
rect 88432 300840 88484 300892
rect 350540 300840 350592 300892
rect 59268 300092 59320 300144
rect 70308 300092 70360 300144
rect 226984 300160 227036 300212
rect 87604 300092 87656 300144
rect 344284 300092 344336 300144
rect 94044 300024 94096 300076
rect 95148 300024 95200 300076
rect 113916 299684 113968 299736
rect 130384 299684 130436 299736
rect 95148 299616 95200 299668
rect 166264 299616 166316 299668
rect 110420 299548 110472 299600
rect 266360 299548 266412 299600
rect 109040 299480 109092 299532
rect 331864 299480 331916 299532
rect 74448 298732 74500 298784
rect 128544 298732 128596 298784
rect 195336 298732 195388 298784
rect 419540 298732 419592 298784
rect 580264 298732 580316 298784
rect 83556 298392 83608 298444
rect 147036 298392 147088 298444
rect 117688 298324 117740 298376
rect 191196 298324 191248 298376
rect 67548 298256 67600 298308
rect 220084 298256 220136 298308
rect 93216 298188 93268 298240
rect 246304 298188 246356 298240
rect 102876 298120 102928 298172
rect 276020 298120 276072 298172
rect 91928 297032 91980 297084
rect 133144 297032 133196 297084
rect 98644 296964 98696 297016
rect 160836 296964 160888 297016
rect 67640 296896 67692 296948
rect 224316 296896 224368 296948
rect 82912 296828 82964 296880
rect 249800 296828 249852 296880
rect 75184 296760 75236 296812
rect 251824 296760 251876 296812
rect 113456 296692 113508 296744
rect 113824 296692 113876 296744
rect 378784 296692 378836 296744
rect 69112 295944 69164 295996
rect 94504 295944 94556 295996
rect 92572 295672 92624 295724
rect 93768 295672 93820 295724
rect 125692 295672 125744 295724
rect 99656 295604 99708 295656
rect 144184 295604 144236 295656
rect 88064 295536 88116 295588
rect 155224 295536 155276 295588
rect 74540 295468 74592 295520
rect 225604 295468 225656 295520
rect 69848 295400 69900 295452
rect 244924 295400 244976 295452
rect 106740 295332 106792 295384
rect 333980 295332 334032 295384
rect 70032 295196 70084 295248
rect 75092 295196 75144 295248
rect 99012 294720 99064 294772
rect 113180 294720 113232 294772
rect 84200 294652 84252 294704
rect 113916 294652 113968 294704
rect 119620 294652 119672 294704
rect 146944 294652 146996 294704
rect 512000 294652 512052 294704
rect 580908 294652 580960 294704
rect 109960 294584 110012 294636
rect 152096 294584 152148 294636
rect 525800 294584 525852 294636
rect 71320 294380 71372 294432
rect 72424 294380 72476 294432
rect 73160 294312 73212 294364
rect 73620 294312 73672 294364
rect 77300 294312 77352 294364
rect 78036 294312 78088 294364
rect 84292 294312 84344 294364
rect 85212 294312 85264 294364
rect 88340 294312 88392 294364
rect 89076 294312 89128 294364
rect 93952 294312 94004 294364
rect 94780 294312 94832 294364
rect 72608 294244 72660 294296
rect 74448 294244 74500 294296
rect 115112 294244 115164 294296
rect 115388 294244 115440 294296
rect 123576 294244 123628 294296
rect 103520 294176 103572 294228
rect 117228 294176 117280 294228
rect 115296 294108 115348 294160
rect 123760 294108 123812 294160
rect 57796 294040 57848 294092
rect 79048 294040 79100 294092
rect 80980 294040 81032 294092
rect 117136 294040 117188 294092
rect 44088 293972 44140 294024
rect 96436 293972 96488 294024
rect 113824 293972 113876 294024
rect 357532 293972 357584 294024
rect 3056 293904 3108 293956
rect 14464 293904 14516 293956
rect 113088 293360 113140 293412
rect 126244 293360 126296 293412
rect 77116 293292 77168 293344
rect 116584 293292 116636 293344
rect 131120 293292 131172 293344
rect 21364 293224 21416 293276
rect 53196 293224 53248 293276
rect 97080 293224 97132 293276
rect 117228 293224 117280 293276
rect 311164 293224 311216 293276
rect 93860 292680 93912 292732
rect 142804 292680 142856 292732
rect 112536 292612 112588 292664
rect 220176 292612 220228 292664
rect 102232 292544 102284 292596
rect 229744 292544 229796 292596
rect 118332 292476 118384 292528
rect 119804 292476 119856 292528
rect 135352 292476 135404 292528
rect 117136 291932 117188 291984
rect 103980 291864 104032 291916
rect 4068 291796 4120 291848
rect 57796 291796 57848 291848
rect 117228 291864 117280 291916
rect 119344 291864 119396 291916
rect 119988 291864 120040 291916
rect 119896 291796 119948 291848
rect 224224 291796 224276 291848
rect 121552 291728 121604 291780
rect 123484 291728 123536 291780
rect 124864 291728 124916 291780
rect 231216 291320 231268 291372
rect 119988 291252 120040 291304
rect 345112 291252 345164 291304
rect 119896 291184 119948 291236
rect 353392 291184 353444 291236
rect 22744 290436 22796 290488
rect 65984 290436 66036 290488
rect 67732 290436 67784 290488
rect 121552 289824 121604 289876
rect 214564 289824 214616 289876
rect 123484 289756 123536 289808
rect 123668 289756 123720 289808
rect 123484 289076 123536 289128
rect 512000 289076 512052 289128
rect 122380 288464 122432 288516
rect 222844 288464 222896 288516
rect 39948 288396 40000 288448
rect 67640 288396 67692 288448
rect 121736 288396 121788 288448
rect 328460 288396 328512 288448
rect 65616 288328 65668 288380
rect 67824 288328 67876 288380
rect 121552 288328 121604 288380
rect 142436 288328 142488 288380
rect 143448 288328 143500 288380
rect 143448 287648 143500 287700
rect 507860 287648 507912 287700
rect 65524 287376 65576 287428
rect 67824 287376 67876 287428
rect 121828 287036 121880 287088
rect 325792 287036 325844 287088
rect 121552 286968 121604 287020
rect 134064 286968 134116 287020
rect 124404 286764 124456 286816
rect 128544 286764 128596 286816
rect 122748 286356 122800 286408
rect 125784 286356 125836 286408
rect 121552 286288 121604 286340
rect 124404 286288 124456 286340
rect 134064 286288 134116 286340
rect 382924 286288 382976 286340
rect 121552 284384 121604 284436
rect 322940 284384 322992 284436
rect 121644 284316 121696 284368
rect 495440 284316 495492 284368
rect 50804 284248 50856 284300
rect 67640 284248 67692 284300
rect 121552 283568 121604 283620
rect 124956 283568 125008 283620
rect 121552 282888 121604 282940
rect 342352 282888 342404 282940
rect 128544 282140 128596 282192
rect 448520 282140 448572 282192
rect 121644 281596 121696 281648
rect 246396 281596 246448 281648
rect 121552 281528 121604 281580
rect 249064 281528 249116 281580
rect 122748 280780 122800 280832
rect 407764 280780 407816 280832
rect 56508 280236 56560 280288
rect 67732 280236 67784 280288
rect 121552 280236 121604 280288
rect 240876 280236 240928 280288
rect 45468 280168 45520 280220
rect 67640 280168 67692 280220
rect 121644 280168 121696 280220
rect 353300 280168 353352 280220
rect 44180 280100 44232 280152
rect 45376 280100 45428 280152
rect 68008 280100 68060 280152
rect 55128 280032 55180 280084
rect 67640 280032 67692 280084
rect 35164 279420 35216 279472
rect 44180 279420 44232 279472
rect 121552 278808 121604 278860
rect 236644 278808 236696 278860
rect 121644 278740 121696 278792
rect 319444 278740 319496 278792
rect 123760 277992 123812 278044
rect 496820 277992 496872 278044
rect 47952 277448 48004 277500
rect 67640 277448 67692 277500
rect 42708 277380 42760 277432
rect 67732 277380 67784 277432
rect 121552 277380 121604 277432
rect 316684 277380 316736 277432
rect 63316 276088 63368 276140
rect 67640 276088 67692 276140
rect 52184 276020 52236 276072
rect 67732 276020 67784 276072
rect 121552 276020 121604 276072
rect 335360 276020 335412 276072
rect 121644 275952 121696 276004
rect 131120 275952 131172 276004
rect 121736 275340 121788 275392
rect 406384 275340 406436 275392
rect 131120 275272 131172 275324
rect 493324 275272 493376 275324
rect 55128 274728 55180 274780
rect 67732 274728 67784 274780
rect 50804 274660 50856 274712
rect 67640 274660 67692 274712
rect 121552 274660 121604 274712
rect 222936 274660 222988 274712
rect 39764 274592 39816 274644
rect 68008 274592 68060 274644
rect 121552 274524 121604 274576
rect 124312 274524 124364 274576
rect 48136 273232 48188 273284
rect 67640 273232 67692 273284
rect 121552 273232 121604 273284
rect 267740 273232 267792 273284
rect 124956 273164 125008 273216
rect 150440 273164 150492 273216
rect 121552 273096 121604 273148
rect 129832 273096 129884 273148
rect 129832 272552 129884 272604
rect 251916 272552 251968 272604
rect 150440 272484 150492 272536
rect 417424 272484 417476 272536
rect 66076 271940 66128 271992
rect 68192 271940 68244 271992
rect 64512 271872 64564 271924
rect 67640 271872 67692 271924
rect 121552 271872 121604 271924
rect 164884 271872 164936 271924
rect 419448 271872 419500 271924
rect 579804 271872 579856 271924
rect 160836 271124 160888 271176
rect 447784 271124 447836 271176
rect 43904 270512 43956 270564
rect 67640 270512 67692 270564
rect 121552 270512 121604 270564
rect 233976 270512 234028 270564
rect 46756 269764 46808 269816
rect 68284 269764 68336 269816
rect 49516 269152 49568 269204
rect 67732 269152 67784 269204
rect 121552 269152 121604 269204
rect 231124 269152 231176 269204
rect 45376 269084 45428 269136
rect 67640 269084 67692 269136
rect 121644 269084 121696 269136
rect 252560 269084 252612 269136
rect 53656 269016 53708 269068
rect 54944 269016 54996 269068
rect 129648 268404 129700 268456
rect 139584 268404 139636 268456
rect 119988 268336 120040 268388
rect 434720 268336 434772 268388
rect 61936 267792 61988 267844
rect 67732 267792 67784 267844
rect 121644 267792 121696 267844
rect 129648 267792 129700 267844
rect 39580 267656 39632 267708
rect 51724 267656 51776 267708
rect 67640 267724 67692 267776
rect 121552 267724 121604 267776
rect 338120 267724 338172 267776
rect 52368 267044 52420 267096
rect 59176 267044 59228 267096
rect 54944 266976 54996 267028
rect 67640 266976 67692 267028
rect 320824 266976 320876 267028
rect 351184 266976 351236 267028
rect 121552 266432 121604 266484
rect 312544 266432 312596 266484
rect 3056 266364 3108 266416
rect 25504 266364 25556 266416
rect 59176 266364 59228 266416
rect 67640 266364 67692 266416
rect 121644 266364 121696 266416
rect 349252 266364 349304 266416
rect 59268 266296 59320 266348
rect 67824 266296 67876 266348
rect 123576 265616 123628 265668
rect 489920 265616 489972 265668
rect 60556 264936 60608 264988
rect 67732 264936 67784 264988
rect 121552 264936 121604 264988
rect 300124 264936 300176 264988
rect 48228 264868 48280 264920
rect 67640 264868 67692 264920
rect 36636 264188 36688 264240
rect 48228 264188 48280 264240
rect 121644 264188 121696 264240
rect 321560 264188 321612 264240
rect 121552 263644 121604 263696
rect 270500 263644 270552 263696
rect 50712 263576 50764 263628
rect 67640 263576 67692 263628
rect 137284 263576 137336 263628
rect 388444 263576 388496 263628
rect 121552 263508 121604 263560
rect 140780 263508 140832 263560
rect 121736 263440 121788 263492
rect 128636 263440 128688 263492
rect 128912 263440 128964 263492
rect 43996 262896 44048 262948
rect 52460 262896 52512 262948
rect 128912 262896 128964 262948
rect 414664 262896 414716 262948
rect 53564 262828 53616 262880
rect 65524 262828 65576 262880
rect 140780 262828 140832 262880
rect 471244 262828 471296 262880
rect 52460 262284 52512 262336
rect 53656 262284 53708 262336
rect 67732 262284 67784 262336
rect 48228 262216 48280 262268
rect 67640 262216 67692 262268
rect 121552 262216 121604 262268
rect 327080 262216 327132 262268
rect 121644 262148 121696 262200
rect 137284 262148 137336 262200
rect 66168 260924 66220 260976
rect 67640 260924 67692 260976
rect 57888 260856 57940 260908
rect 67732 260856 67784 260908
rect 134616 260856 134668 260908
rect 134892 260856 134944 260908
rect 232504 260856 232556 260908
rect 60648 260788 60700 260840
rect 67640 260788 67692 260840
rect 121552 260788 121604 260840
rect 146300 260788 146352 260840
rect 146760 260788 146812 260840
rect 121736 260176 121788 260228
rect 323032 260176 323084 260228
rect 146760 260108 146812 260160
rect 517612 260108 517664 260160
rect 52368 259428 52420 259480
rect 67640 259428 67692 259480
rect 121552 259428 121604 259480
rect 245016 259428 245068 259480
rect 121644 259360 121696 259412
rect 134892 259360 134944 259412
rect 126244 258680 126296 258732
rect 547880 258680 547932 258732
rect 57796 258136 57848 258188
rect 67732 258136 67784 258188
rect 56324 258068 56376 258120
rect 67640 258068 67692 258120
rect 121552 258068 121604 258120
rect 349160 258068 349212 258120
rect 547880 258068 547932 258120
rect 580172 258068 580224 258120
rect 36544 258000 36596 258052
rect 67916 258000 67968 258052
rect 15844 257320 15896 257372
rect 36544 257320 36596 257372
rect 124864 257320 124916 257372
rect 485780 257320 485832 257372
rect 59268 256708 59320 256760
rect 67640 256708 67692 256760
rect 121644 256708 121696 256760
rect 260840 256708 260892 256760
rect 121552 256640 121604 256692
rect 154580 256640 154632 256692
rect 154580 256028 154632 256080
rect 399484 256028 399536 256080
rect 159364 255960 159416 256012
rect 520924 255960 520976 256012
rect 65984 255348 66036 255400
rect 67640 255348 67692 255400
rect 53380 255280 53432 255332
rect 67732 255280 67784 255332
rect 3424 255212 3476 255264
rect 33140 255212 33192 255264
rect 57612 255212 57664 255264
rect 67640 255212 67692 255264
rect 33140 254532 33192 254584
rect 34428 254532 34480 254584
rect 58624 254532 58676 254584
rect 187056 254532 187108 254584
rect 508504 254532 508556 254584
rect 67640 253920 67692 253972
rect 121552 253920 121604 253972
rect 284300 253920 284352 253972
rect 53748 253852 53800 253904
rect 60004 253852 60056 253904
rect 17224 253172 17276 253224
rect 35716 253172 35768 253224
rect 56232 253172 56284 253224
rect 121644 253172 121696 253224
rect 400864 253172 400916 253224
rect 121552 252628 121604 252680
rect 258080 252628 258132 252680
rect 56232 252560 56284 252612
rect 67640 252560 67692 252612
rect 121644 252560 121696 252612
rect 316776 252560 316828 252612
rect 121552 252492 121604 252544
rect 143724 252492 143776 252544
rect 144828 252492 144880 252544
rect 144828 251812 144880 251864
rect 472624 251812 472676 251864
rect 61844 251268 61896 251320
rect 67640 251268 67692 251320
rect 53472 251200 53524 251252
rect 67732 251200 67784 251252
rect 121552 251200 121604 251252
rect 327264 251200 327316 251252
rect 129648 250452 129700 250504
rect 478880 250452 478932 250504
rect 122104 249840 122156 249892
rect 124312 249840 124364 249892
rect 60464 249772 60516 249824
rect 67640 249772 67692 249824
rect 121552 249772 121604 249824
rect 243544 249772 243596 249824
rect 41144 249024 41196 249076
rect 57704 249024 57756 249076
rect 169024 249024 169076 249076
rect 517520 249024 517572 249076
rect 57704 248480 57756 248532
rect 67732 248480 67784 248532
rect 54852 248412 54904 248464
rect 67640 248412 67692 248464
rect 121552 248412 121604 248464
rect 345204 248412 345256 248464
rect 121460 248344 121512 248396
rect 121736 248344 121788 248396
rect 63224 247120 63276 247172
rect 67640 247120 67692 247172
rect 121460 247120 121512 247172
rect 235264 247120 235316 247172
rect 60648 247052 60700 247104
rect 67732 247052 67784 247104
rect 124036 247052 124088 247104
rect 494244 247052 494296 247104
rect 124312 246372 124364 246424
rect 443000 246372 443052 246424
rect 121644 246304 121696 246356
rect 499672 246304 499724 246356
rect 63408 245692 63460 245744
rect 67640 245692 67692 245744
rect 121552 245692 121604 245744
rect 159364 245692 159416 245744
rect 55036 245556 55088 245608
rect 61384 245624 61436 245676
rect 67732 245624 67784 245676
rect 121460 245624 121512 245676
rect 269120 245624 269172 245676
rect 135904 244944 135956 244996
rect 227076 244944 227128 244996
rect 122288 244876 122340 244928
rect 328552 244876 328604 244928
rect 263600 244264 263652 244316
rect 579620 244264 579672 244316
rect 579988 244264 580040 244316
rect 62028 244196 62080 244248
rect 65892 244196 65944 244248
rect 231216 243652 231268 243704
rect 318156 243652 318208 243704
rect 232596 243584 232648 243636
rect 370504 243584 370556 243636
rect 121736 243516 121788 243568
rect 498292 243516 498344 243568
rect 48044 242836 48096 242888
rect 54484 242836 54536 242888
rect 67640 242972 67692 243024
rect 121460 242972 121512 243024
rect 206376 242972 206428 243024
rect 127624 242904 127676 242956
rect 231308 242904 231360 242956
rect 121460 242836 121512 242888
rect 147680 242836 147732 242888
rect 263600 242836 263652 242888
rect 121552 242768 121604 242820
rect 140780 242768 140832 242820
rect 140780 242156 140832 242208
rect 413284 242156 413336 242208
rect 62028 241476 62080 241528
rect 67640 241476 67692 241528
rect 121644 240728 121696 240780
rect 321652 240728 321704 240780
rect 121460 240184 121512 240236
rect 238116 240184 238168 240236
rect 119896 240116 119948 240168
rect 331220 240116 331272 240168
rect 3148 240048 3200 240100
rect 33600 240048 33652 240100
rect 75920 239776 75972 239828
rect 77104 239776 77156 239828
rect 80060 239776 80112 239828
rect 80968 239776 81020 239828
rect 92480 239776 92532 239828
rect 93204 239776 93256 239828
rect 95240 239776 95292 239828
rect 96424 239776 96476 239828
rect 96620 239776 96672 239828
rect 97712 239776 97764 239828
rect 100760 239776 100812 239828
rect 101576 239776 101628 239828
rect 104900 239776 104952 239828
rect 106084 239776 106136 239828
rect 114560 239776 114612 239828
rect 115744 239776 115796 239828
rect 117320 239776 117372 239828
rect 118332 239776 118384 239828
rect 124220 239776 124272 239828
rect 63408 239504 63460 239556
rect 72424 239504 72476 239556
rect 61936 239436 61988 239488
rect 98644 239436 98696 239488
rect 33600 239368 33652 239420
rect 34336 239368 34388 239420
rect 92664 239368 92716 239420
rect 113180 239300 113232 239352
rect 114468 239300 114520 239352
rect 65892 238824 65944 238876
rect 76012 238824 76064 238876
rect 76472 238824 76524 238876
rect 58624 238756 58676 238808
rect 112536 238756 112588 238808
rect 121460 238756 121512 238808
rect 346400 238756 346452 238808
rect 50896 238688 50948 238740
rect 98368 238688 98420 238740
rect 25504 238620 25556 238672
rect 56416 238620 56468 238672
rect 86776 238620 86828 238672
rect 91928 238620 91980 238672
rect 123484 238620 123536 238672
rect 92664 238552 92716 238604
rect 103520 238552 103572 238604
rect 105452 238212 105504 238264
rect 181444 238212 181496 238264
rect 251916 238212 251968 238264
rect 381544 238212 381596 238264
rect 67456 238144 67508 238196
rect 259460 238144 259512 238196
rect 69940 238076 69992 238128
rect 77944 238076 77996 238128
rect 102232 238076 102284 238128
rect 339592 238076 339644 238128
rect 73896 238008 73948 238060
rect 332600 238008 332652 238060
rect 86224 237464 86276 237516
rect 86776 237464 86828 237516
rect 85488 237396 85540 237448
rect 86316 237396 86368 237448
rect 89996 237396 90048 237448
rect 91744 237396 91796 237448
rect 103520 237396 103572 237448
rect 104164 237396 104216 237448
rect 116584 237396 116636 237448
rect 117688 237396 117740 237448
rect 69204 237328 69256 237380
rect 150532 237328 150584 237380
rect 52276 237260 52328 237312
rect 116584 237260 116636 237312
rect 50988 237192 51040 237244
rect 81624 237192 81676 237244
rect 110604 237192 110656 237244
rect 132500 237192 132552 237244
rect 58992 237124 59044 237176
rect 86132 237124 86184 237176
rect 150532 236648 150584 236700
rect 452660 236648 452712 236700
rect 81624 235968 81676 236020
rect 82084 235968 82136 236020
rect 110604 235968 110656 236020
rect 111064 235968 111116 236020
rect 89628 235900 89680 235952
rect 125600 235900 125652 235952
rect 63224 235356 63276 235408
rect 239404 235356 239456 235408
rect 251824 235356 251876 235408
rect 277400 235356 277452 235408
rect 60464 235288 60516 235340
rect 278780 235288 278832 235340
rect 113272 235220 113324 235272
rect 340972 235220 341024 235272
rect 46848 234540 46900 234592
rect 109684 234540 109736 234592
rect 61844 234064 61896 234116
rect 182824 234064 182876 234116
rect 65984 233996 66036 234048
rect 251272 233996 251324 234048
rect 112536 233928 112588 233980
rect 445760 233928 445812 233980
rect 86132 233860 86184 233912
rect 502340 233860 502392 233912
rect 93860 233724 93912 233776
rect 94044 233724 94096 233776
rect 77760 232568 77812 232620
rect 352012 232568 352064 232620
rect 56232 232500 56284 232552
rect 403624 232500 403676 232552
rect 515404 232500 515456 232552
rect 579620 232500 579672 232552
rect 49608 231752 49660 231804
rect 107292 231752 107344 231804
rect 95332 231684 95384 231736
rect 126980 231684 127032 231736
rect 127440 231684 127492 231736
rect 95056 231140 95108 231192
rect 347872 231140 347924 231192
rect 127440 231072 127492 231124
rect 393964 231072 394016 231124
rect 84200 229916 84252 229968
rect 84476 229916 84528 229968
rect 66076 229848 66128 229900
rect 251364 229848 251416 229900
rect 108580 229780 108632 229832
rect 331312 229780 331364 229832
rect 60004 229712 60056 229764
rect 468484 229712 468536 229764
rect 83464 229032 83516 229084
rect 149060 229032 149112 229084
rect 82820 228964 82872 229016
rect 128360 228964 128412 229016
rect 149060 228556 149112 228608
rect 171784 228556 171836 228608
rect 57888 228488 57940 228540
rect 314016 228488 314068 228540
rect 53472 228420 53524 228472
rect 339500 228420 339552 228472
rect 128360 228352 128412 228404
rect 513380 228352 513432 228404
rect 91100 227672 91152 227724
rect 131212 227672 131264 227724
rect 131764 227672 131816 227724
rect 71228 227060 71280 227112
rect 255412 227060 255464 227112
rect 131212 226992 131264 227044
rect 342996 226992 343048 227044
rect 64512 225632 64564 225684
rect 251180 225632 251232 225684
rect 80060 225564 80112 225616
rect 328644 225564 328696 225616
rect 75736 224884 75788 224936
rect 142252 224884 142304 224936
rect 143448 224884 143500 224936
rect 55128 224340 55180 224392
rect 151084 224340 151136 224392
rect 90088 224272 90140 224324
rect 255596 224272 255648 224324
rect 143448 224204 143500 224256
rect 333336 224204 333388 224256
rect 109684 223592 109736 223644
rect 457444 223592 457496 223644
rect 47952 222844 48004 222896
rect 276112 222844 276164 222896
rect 103612 221552 103664 221604
rect 327172 221552 327224 221604
rect 61384 221484 61436 221536
rect 371884 221484 371936 221536
rect 4804 221416 4856 221468
rect 83464 221416 83516 221468
rect 104164 221416 104216 221468
rect 466460 221416 466512 221468
rect 74632 220056 74684 220108
rect 281540 220056 281592 220108
rect 57704 218764 57756 218816
rect 489184 218764 489236 218816
rect 54944 218696 54996 218748
rect 503720 218696 503772 218748
rect 520924 218696 520976 218748
rect 580172 218696 580224 218748
rect 54852 217336 54904 217388
rect 246488 217336 246540 217388
rect 59084 217268 59136 217320
rect 488540 217268 488592 217320
rect 81532 216588 81584 216640
rect 151820 216588 151872 216640
rect 153108 216588 153160 216640
rect 77944 215976 77996 216028
rect 315396 215976 315448 216028
rect 153108 215908 153160 215960
rect 473360 215908 473412 215960
rect 113180 215228 113232 215280
rect 147772 215228 147824 215280
rect 78772 214684 78824 214736
rect 314108 214684 314160 214736
rect 147772 214616 147824 214668
rect 501052 214616 501104 214668
rect 3424 214548 3476 214600
rect 36636 214548 36688 214600
rect 396724 214548 396776 214600
rect 71780 213324 71832 213376
rect 329932 213324 329984 213376
rect 42708 213256 42760 213308
rect 304356 213256 304408 213308
rect 93952 213188 94004 213240
rect 232596 213188 232648 213240
rect 238024 213188 238076 213240
rect 512092 213188 512144 213240
rect 62028 211896 62080 211948
rect 267832 211896 267884 211948
rect 76012 211828 76064 211880
rect 336096 211828 336148 211880
rect 52368 211760 52420 211812
rect 338212 211760 338264 211812
rect 114560 210536 114612 210588
rect 325884 210536 325936 210588
rect 53564 210468 53616 210520
rect 273260 210468 273312 210520
rect 75920 210400 75972 210452
rect 330116 210400 330168 210452
rect 100852 209176 100904 209228
rect 252652 209176 252704 209228
rect 74540 209108 74592 209160
rect 323124 209108 323176 209160
rect 53656 209040 53708 209092
rect 480260 209040 480312 209092
rect 106280 208292 106332 208344
rect 138020 208292 138072 208344
rect 87052 207748 87104 207800
rect 249892 207748 249944 207800
rect 60648 207680 60700 207732
rect 263600 207680 263652 207732
rect 138020 207612 138072 207664
rect 354036 207612 354088 207664
rect 86316 206320 86368 206372
rect 264980 206320 265032 206372
rect 86224 206252 86276 206304
rect 498384 206252 498436 206304
rect 508504 206252 508556 206304
rect 580172 206252 580224 206304
rect 98092 205572 98144 205624
rect 143540 205572 143592 205624
rect 144828 205572 144880 205624
rect 3240 204960 3292 205012
rect 120172 204960 120224 205012
rect 144828 204960 144880 205012
rect 392584 204960 392636 205012
rect 50712 204892 50764 204944
rect 312636 204892 312688 204944
rect 100760 203736 100812 203788
rect 254216 203736 254268 203788
rect 91744 203668 91796 203720
rect 263692 203668 263744 203720
rect 90364 203600 90416 203652
rect 349344 203600 349396 203652
rect 195336 203532 195388 203584
rect 501236 203532 501288 203584
rect 99472 202240 99524 202292
rect 255504 202240 255556 202292
rect 98644 202172 98696 202224
rect 269212 202172 269264 202224
rect 7564 202104 7616 202156
rect 125692 202104 125744 202156
rect 465080 202104 465132 202156
rect 50804 200880 50856 200932
rect 259644 200880 259696 200932
rect 117320 200812 117372 200864
rect 337476 200812 337528 200864
rect 70400 200744 70452 200796
rect 334164 200744 334216 200796
rect 133144 199656 133196 199708
rect 262312 199656 262364 199708
rect 115940 199588 115992 199640
rect 249984 199588 250036 199640
rect 77300 199520 77352 199572
rect 266452 199520 266504 199572
rect 45376 199452 45428 199504
rect 318248 199452 318300 199504
rect 403624 199452 403676 199504
rect 459560 199452 459612 199504
rect 233884 199384 233936 199436
rect 509240 199384 509292 199436
rect 92572 198092 92624 198144
rect 259552 198092 259604 198144
rect 52184 198024 52236 198076
rect 238024 198024 238076 198076
rect 231308 197956 231360 198008
rect 510620 197956 510672 198008
rect 111800 196800 111852 196852
rect 254032 196800 254084 196852
rect 57796 196732 57848 196784
rect 271880 196732 271932 196784
rect 92480 196664 92532 196716
rect 328736 196664 328788 196716
rect 69020 196596 69072 196648
rect 496912 196596 496964 196648
rect 56324 195440 56376 195492
rect 260932 195440 260984 195492
rect 103704 195372 103756 195424
rect 321744 195372 321796 195424
rect 49516 195304 49568 195356
rect 273352 195304 273404 195356
rect 89628 195236 89680 195288
rect 506572 195236 506624 195288
rect 102140 193876 102192 193928
rect 252836 193876 252888 193928
rect 93860 193808 93912 193860
rect 352104 193808 352156 193860
rect 3424 193196 3476 193248
rect 4068 193196 4120 193248
rect 509332 193196 509384 193248
rect 221464 192720 221516 192772
rect 280160 192720 280212 192772
rect 43904 192652 43956 192704
rect 199384 192652 199436 192704
rect 214656 192652 214708 192704
rect 277492 192652 277544 192704
rect 196716 192584 196768 192636
rect 471980 192584 472032 192636
rect 53380 192516 53432 192568
rect 346492 192516 346544 192568
rect 54484 192448 54536 192500
rect 469220 192448 469272 192500
rect 224316 191292 224368 191344
rect 276204 191292 276256 191344
rect 48136 191224 48188 191276
rect 267924 191224 267976 191276
rect 46756 191156 46808 191208
rect 343640 191156 343692 191208
rect 419632 191156 419684 191208
rect 580172 191156 580224 191208
rect 119344 191088 119396 191140
rect 494336 191088 494388 191140
rect 100668 190544 100720 190596
rect 170496 190544 170548 190596
rect 106188 190476 106240 190528
rect 195336 190476 195388 190528
rect 249064 190000 249116 190052
rect 271972 190000 272024 190052
rect 155224 189932 155276 189984
rect 265164 189932 265216 189984
rect 78680 189864 78732 189916
rect 258172 189864 258224 189916
rect 59268 189796 59320 189848
rect 350632 189796 350684 189848
rect 116584 189728 116636 189780
rect 505284 189728 505336 189780
rect 102048 189048 102100 189100
rect 173164 189048 173216 189100
rect 3516 188844 3568 188896
rect 7564 188844 7616 188896
rect 213276 188504 213328 188556
rect 274640 188504 274692 188556
rect 130384 188436 130436 188488
rect 249340 188436 249392 188488
rect 99380 188368 99432 188420
rect 327356 188368 327408 188420
rect 63316 188300 63368 188352
rect 324320 188300 324372 188352
rect 135904 187688 135956 187740
rect 214656 187688 214708 187740
rect 229744 187280 229796 187332
rect 256700 187280 256752 187332
rect 222936 187212 222988 187264
rect 274732 187212 274784 187264
rect 88340 187144 88392 187196
rect 325976 187144 326028 187196
rect 73160 187076 73212 187128
rect 321836 187076 321888 187128
rect 104900 187008 104952 187060
rect 354680 187008 354732 187060
rect 72424 186940 72476 186992
rect 345296 186940 345348 186992
rect 419264 186940 419316 186992
rect 580264 186940 580316 186992
rect 133144 186328 133196 186380
rect 209228 186328 209280 186380
rect 227076 185784 227128 185836
rect 270684 185784 270736 185836
rect 151084 185716 151136 185768
rect 336740 185716 336792 185768
rect 48228 185648 48280 185700
rect 247684 185648 247736 185700
rect 67548 185580 67600 185632
rect 318340 185580 318392 185632
rect 422944 185580 422996 185632
rect 450544 185580 450596 185632
rect 124128 184968 124180 185020
rect 167828 184968 167880 185020
rect 126888 184900 126940 184952
rect 214748 184900 214800 184952
rect 429936 184832 429988 184884
rect 430580 184832 430632 184884
rect 152464 184424 152516 184476
rect 187056 184424 187108 184476
rect 225604 184424 225656 184476
rect 269304 184424 269356 184476
rect 86960 184356 87012 184408
rect 196808 184356 196860 184408
rect 206376 184356 206428 184408
rect 335452 184356 335504 184408
rect 96712 184288 96764 184340
rect 263784 184288 263836 184340
rect 467104 184288 467156 184340
rect 499764 184288 499816 184340
rect 95240 184220 95292 184272
rect 321284 184220 321336 184272
rect 472624 184220 472676 184272
rect 506664 184220 506716 184272
rect 107660 184152 107712 184204
rect 338304 184152 338356 184204
rect 464344 184152 464396 184204
rect 512184 184152 512236 184204
rect 345020 184016 345072 184068
rect 345664 184016 345716 184068
rect 121368 183540 121420 183592
rect 166356 183540 166408 183592
rect 345664 183540 345716 183592
rect 499856 183540 499908 183592
rect 240784 183132 240836 183184
rect 261116 183132 261168 183184
rect 220176 183064 220228 183116
rect 268016 183064 268068 183116
rect 142804 182996 142856 183048
rect 245384 182996 245436 183048
rect 110420 182928 110472 182980
rect 252744 182928 252796 182980
rect 45468 182860 45520 182912
rect 265072 182860 265124 182912
rect 316684 182860 316736 182912
rect 339684 182860 339736 182912
rect 96620 182792 96672 182844
rect 206376 182792 206428 182844
rect 232504 182792 232556 182844
rect 502524 182792 502576 182844
rect 130752 182248 130804 182300
rect 166540 182248 166592 182300
rect 110696 182180 110748 182232
rect 169024 182180 169076 182232
rect 457444 182112 457496 182164
rect 458180 182112 458232 182164
rect 475384 182112 475436 182164
rect 476580 182112 476632 182164
rect 160744 181704 160796 181756
rect 203524 181704 203576 181756
rect 233976 181704 234028 181756
rect 256884 181704 256936 181756
rect 489184 181704 489236 181756
rect 492864 181704 492916 181756
rect 202236 181636 202288 181688
rect 334072 181636 334124 181688
rect 483664 181636 483716 181688
rect 502432 181636 502484 181688
rect 171784 181568 171836 181620
rect 439412 181568 439464 181620
rect 482284 181568 482336 181620
rect 502616 181568 502668 181620
rect 56508 181500 56560 181552
rect 343732 181500 343784 181552
rect 471244 181500 471296 181552
rect 508044 181500 508096 181552
rect 166264 181432 166316 181484
rect 483572 181432 483624 181484
rect 485044 181432 485096 181484
rect 505192 181432 505244 181484
rect 447784 181296 447836 181348
rect 451372 181296 451424 181348
rect 132408 181024 132460 181076
rect 164976 181024 165028 181076
rect 118516 180956 118568 181008
rect 171876 180956 171928 181008
rect 114376 180888 114428 180940
rect 167736 180888 167788 180940
rect 97080 180820 97132 180872
rect 170588 180820 170640 180872
rect 385684 180820 385736 180872
rect 491300 180820 491352 180872
rect 246396 180412 246448 180464
rect 249064 180412 249116 180464
rect 314016 180412 314068 180464
rect 331496 180412 331548 180464
rect 236644 180344 236696 180396
rect 249432 180344 249484 180396
rect 316776 180344 316828 180396
rect 341156 180344 341208 180396
rect 232596 180276 232648 180328
rect 256792 180276 256844 180328
rect 305736 180276 305788 180328
rect 333244 180276 333296 180328
rect 159364 180208 159416 180260
rect 259736 180208 259788 180260
rect 311164 180208 311216 180260
rect 343824 180208 343876 180260
rect 493324 180208 493376 180260
rect 507952 180208 508004 180260
rect 29644 180140 29696 180192
rect 109684 180140 109736 180192
rect 226984 180140 227036 180192
rect 389824 180140 389876 180192
rect 468484 180140 468536 180192
rect 503904 180140 503956 180192
rect 82084 180072 82136 180124
rect 495624 180072 495676 180124
rect 407764 180004 407816 180056
rect 408408 180004 408460 180056
rect 114008 179528 114060 179580
rect 166264 179528 166316 179580
rect 115848 179460 115900 179512
rect 167920 179460 167972 179512
rect 108120 179392 108172 179444
rect 169208 179392 169260 179444
rect 408408 179392 408460 179444
rect 574744 179392 574796 179444
rect 235264 178984 235316 179036
rect 250076 178984 250128 179036
rect 238116 178916 238168 178968
rect 258356 178916 258408 178968
rect 84200 178848 84252 178900
rect 323216 178848 323268 178900
rect 69112 178780 69164 178832
rect 324412 178780 324464 178832
rect 66168 178712 66220 178764
rect 324504 178712 324556 178764
rect 331864 178712 331916 178764
rect 342444 178712 342496 178764
rect 100760 178644 100812 178696
rect 133880 178644 133932 178696
rect 505100 178644 505152 178696
rect 122104 178032 122156 178084
rect 166448 178032 166500 178084
rect 360936 178032 360988 178084
rect 416780 178032 416832 178084
rect 119528 177964 119580 178016
rect 135904 177964 135956 178016
rect 243544 177964 243596 178016
rect 249156 177964 249208 178016
rect 109960 177896 110012 177948
rect 121460 177896 121512 177948
rect 127900 177896 127952 177948
rect 133144 177896 133196 177948
rect 245384 177896 245436 177948
rect 249248 177896 249300 177948
rect 318340 177556 318392 177608
rect 329840 177556 329892 177608
rect 246304 177488 246356 177540
rect 261024 177488 261076 177540
rect 314108 177488 314160 177540
rect 332692 177488 332744 177540
rect 240876 177420 240928 177472
rect 262496 177420 262548 177472
rect 318156 177420 318208 177472
rect 336832 177420 336884 177472
rect 231124 177352 231176 177404
rect 258264 177352 258316 177404
rect 313924 177352 313976 177404
rect 341064 177352 341116 177404
rect 7564 177284 7616 177336
rect 100760 177284 100812 177336
rect 214564 177284 214616 177336
rect 270592 177284 270644 177336
rect 289084 177284 289136 177336
rect 338764 177284 338816 177336
rect 134432 177012 134484 177064
rect 165528 177012 165580 177064
rect 124496 176944 124548 176996
rect 170680 176944 170732 176996
rect 497004 176944 497056 176996
rect 498476 176944 498528 176996
rect 107016 176876 107068 176928
rect 165252 176876 165304 176928
rect 103336 176808 103388 176860
rect 169116 176808 169168 176860
rect 136088 176740 136140 176792
rect 213920 176740 213972 176792
rect 133144 176672 133196 176724
rect 356704 176672 356756 176724
rect 416780 176672 416832 176724
rect 497004 176672 497056 176724
rect 500960 176672 501012 176724
rect 214012 176604 214064 176656
rect 128176 176264 128228 176316
rect 167000 176264 167052 176316
rect 158904 176196 158956 176248
rect 211896 176196 211948 176248
rect 148232 176128 148284 176180
rect 209136 176128 209188 176180
rect 104624 176060 104676 176112
rect 169300 176060 169352 176112
rect 244924 176060 244976 176112
rect 254124 176060 254176 176112
rect 315396 176060 315448 176112
rect 330024 176060 330076 176112
rect 129464 175992 129516 176044
rect 214104 175992 214156 176044
rect 245016 175992 245068 176044
rect 262404 175992 262456 176044
rect 315304 175992 315356 176044
rect 334256 175992 334308 176044
rect 14464 175924 14516 175976
rect 111064 175924 111116 175976
rect 116952 175924 117004 175976
rect 213368 175924 213420 175976
rect 239404 175924 239456 175976
rect 262220 175924 262272 175976
rect 312544 175924 312596 175976
rect 331404 175924 331456 175976
rect 319444 175584 319496 175636
rect 321468 175584 321520 175636
rect 165528 175176 165580 175228
rect 213920 175176 213972 175228
rect 165252 174496 165304 174548
rect 214564 174496 214616 174548
rect 497004 174224 497056 174276
rect 501144 174224 501196 174276
rect 267004 174088 267056 174140
rect 307668 174088 307720 174140
rect 302884 174020 302936 174072
rect 307576 174020 307628 174072
rect 297456 173952 297508 174004
rect 307484 173952 307536 174004
rect 355324 173884 355376 173936
rect 416780 173884 416832 173936
rect 164976 173816 165028 173868
rect 213920 173816 213972 173868
rect 324320 173816 324372 173868
rect 333980 173816 334032 173868
rect 166540 173748 166592 173800
rect 214012 173748 214064 173800
rect 285036 172660 285088 172712
rect 307576 172660 307628 172712
rect 271144 172592 271196 172644
rect 307484 172592 307536 172644
rect 264244 172524 264296 172576
rect 307668 172524 307720 172576
rect 167000 172456 167052 172508
rect 213920 172456 213972 172508
rect 252468 172456 252520 172508
rect 267740 172456 267792 172508
rect 252376 172388 252428 172440
rect 256884 172388 256936 172440
rect 304448 171232 304500 171284
rect 307668 171232 307720 171284
rect 286416 171164 286468 171216
rect 306564 171164 306616 171216
rect 273996 171096 274048 171148
rect 307300 171096 307352 171148
rect 353944 171096 353996 171148
rect 416780 171096 416832 171148
rect 209228 171028 209280 171080
rect 213920 171028 213972 171080
rect 252376 171028 252428 171080
rect 262220 171028 262272 171080
rect 324320 171028 324372 171080
rect 334256 171028 334308 171080
rect 252468 170960 252520 171012
rect 261116 170960 261168 171012
rect 497004 170756 497056 170808
rect 499856 170756 499908 170808
rect 252468 170076 252520 170128
rect 259644 170076 259696 170128
rect 307024 170076 307076 170128
rect 308588 170076 308640 170128
rect 289268 169872 289320 169924
rect 307300 169872 307352 169924
rect 268568 169804 268620 169856
rect 307576 169804 307628 169856
rect 262864 169736 262916 169788
rect 307668 169736 307720 169788
rect 334624 169736 334676 169788
rect 416780 169736 416832 169788
rect 167828 169668 167880 169720
rect 214012 169668 214064 169720
rect 170680 169600 170732 169652
rect 213920 169600 213972 169652
rect 252468 169600 252520 169652
rect 263784 169600 263836 169652
rect 252376 169532 252428 169584
rect 265164 169532 265216 169584
rect 290556 168988 290608 169040
rect 307116 168988 307168 169040
rect 278228 168444 278280 168496
rect 307668 168444 307720 168496
rect 267096 168376 267148 168428
rect 307484 168376 307536 168428
rect 166448 168308 166500 168360
rect 213920 168308 213972 168360
rect 252376 168308 252428 168360
rect 262312 168308 262364 168360
rect 324320 168308 324372 168360
rect 329840 168308 329892 168360
rect 497004 168308 497056 168360
rect 502340 168308 502392 168360
rect 503628 168308 503680 168360
rect 166356 168240 166408 168292
rect 214012 168240 214064 168292
rect 252468 167900 252520 167952
rect 258080 167900 258132 167952
rect 265808 167628 265860 167680
rect 307576 167628 307628 167680
rect 503628 167628 503680 167680
rect 543004 167628 543056 167680
rect 287888 167084 287940 167136
rect 307668 167084 307720 167136
rect 257344 167016 257396 167068
rect 307484 167016 307536 167068
rect 171876 166948 171928 167000
rect 213920 166948 213972 167000
rect 324320 166948 324372 167000
rect 335544 166948 335596 167000
rect 497004 166948 497056 167000
rect 505284 166948 505336 167000
rect 252468 166336 252520 166388
rect 258356 166336 258408 166388
rect 269764 166268 269816 166320
rect 307576 166268 307628 166320
rect 505284 166268 505336 166320
rect 544384 166268 544436 166320
rect 252468 166064 252520 166116
rect 259552 166064 259604 166116
rect 258724 165588 258776 165640
rect 306748 165588 306800 165640
rect 546500 165588 546552 165640
rect 580172 165588 580224 165640
rect 167920 165520 167972 165572
rect 213920 165520 213972 165572
rect 252284 165520 252336 165572
rect 276112 165520 276164 165572
rect 324412 165520 324464 165572
rect 339592 165520 339644 165572
rect 497096 165520 497148 165572
rect 507860 165520 507912 165572
rect 167736 165452 167788 165504
rect 214012 165452 214064 165504
rect 252468 165452 252520 165504
rect 266360 165452 266412 165504
rect 324320 165452 324372 165504
rect 330024 165452 330076 165504
rect 252376 165384 252428 165436
rect 263692 165384 263744 165436
rect 264428 164840 264480 164892
rect 307668 164840 307720 164892
rect 497004 164840 497056 164892
rect 503904 164840 503956 164892
rect 507860 164840 507912 164892
rect 536104 164840 536156 164892
rect 503904 164432 503956 164484
rect 504456 164432 504508 164484
rect 294696 164296 294748 164348
rect 307576 164296 307628 164348
rect 260288 164228 260340 164280
rect 307668 164228 307720 164280
rect 340236 164228 340288 164280
rect 416780 164228 416832 164280
rect 166264 164160 166316 164212
rect 213920 164160 213972 164212
rect 252376 164160 252428 164212
rect 273260 164160 273312 164212
rect 324412 164160 324464 164212
rect 338212 164160 338264 164212
rect 497004 164160 497056 164212
rect 517612 164160 517664 164212
rect 546500 164160 546552 164212
rect 252284 164092 252336 164144
rect 270500 164092 270552 164144
rect 324320 164092 324372 164144
rect 331496 164092 331548 164144
rect 252468 164024 252520 164076
rect 269304 164024 269356 164076
rect 253296 163480 253348 163532
rect 267924 163480 267976 163532
rect 268384 163480 268436 163532
rect 307484 163480 307536 163532
rect 304356 163004 304408 163056
rect 307668 163004 307720 163056
rect 298928 162936 298980 162988
rect 307576 162936 307628 162988
rect 261668 162868 261720 162920
rect 307116 162868 307168 162920
rect 169024 162800 169076 162852
rect 213920 162800 213972 162852
rect 252376 162800 252428 162852
rect 266452 162800 266504 162852
rect 324320 162800 324372 162852
rect 342444 162800 342496 162852
rect 497004 162800 497056 162852
rect 508504 162800 508556 162852
rect 252468 162732 252520 162784
rect 265072 162732 265124 162784
rect 324412 162732 324464 162784
rect 335452 162732 335504 162784
rect 250444 162188 250496 162240
rect 258264 162188 258316 162240
rect 250536 162120 250588 162172
rect 260932 162120 260984 162172
rect 296076 161576 296128 161628
rect 307576 161576 307628 161628
rect 272708 161508 272760 161560
rect 307668 161508 307720 161560
rect 261484 161440 261536 161492
rect 307300 161440 307352 161492
rect 342904 161440 342956 161492
rect 416780 161440 416832 161492
rect 169208 161372 169260 161424
rect 213920 161372 213972 161424
rect 252468 161372 252520 161424
rect 271972 161372 272024 161424
rect 324320 161372 324372 161424
rect 340880 161372 340932 161424
rect 497004 161372 497056 161424
rect 515404 161372 515456 161424
rect 283748 160692 283800 160744
rect 307392 160692 307444 160744
rect 263048 160148 263100 160200
rect 307576 160148 307628 160200
rect 259000 160080 259052 160132
rect 307668 160080 307720 160132
rect 169300 160012 169352 160064
rect 214012 160012 214064 160064
rect 252468 160012 252520 160064
rect 269212 160012 269264 160064
rect 324320 160012 324372 160064
rect 334164 160012 334216 160064
rect 497004 160012 497056 160064
rect 512000 160012 512052 160064
rect 195336 159944 195388 159996
rect 213920 159944 213972 159996
rect 251732 159944 251784 159996
rect 254124 159944 254176 159996
rect 497096 159944 497148 159996
rect 504364 159944 504416 159996
rect 250628 159400 250680 159452
rect 259736 159400 259788 159452
rect 253480 159332 253532 159384
rect 258172 159332 258224 159384
rect 292028 158856 292080 158908
rect 307116 158856 307168 158908
rect 265716 158788 265768 158840
rect 307668 158788 307720 158840
rect 260196 158720 260248 158772
rect 306748 158720 306800 158772
rect 336004 158720 336056 158772
rect 416780 158720 416832 158772
rect 169116 158652 169168 158704
rect 213920 158652 213972 158704
rect 252468 158652 252520 158704
rect 261024 158652 261076 158704
rect 324412 158652 324464 158704
rect 343824 158652 343876 158704
rect 497004 158652 497056 158704
rect 519544 158652 519596 158704
rect 324320 158584 324372 158636
rect 331404 158584 331456 158636
rect 251824 158040 251876 158092
rect 259460 158040 259512 158092
rect 300216 157496 300268 157548
rect 306564 157496 306616 157548
rect 276756 157428 276808 157480
rect 307668 157428 307720 157480
rect 258816 157360 258868 157412
rect 307576 157360 307628 157412
rect 341524 157360 341576 157412
rect 416780 157360 416832 157412
rect 170496 157292 170548 157344
rect 214012 157292 214064 157344
rect 252468 157292 252520 157344
rect 262404 157292 262456 157344
rect 324320 157292 324372 157344
rect 336832 157292 336884 157344
rect 497004 157292 497056 157344
rect 582380 157292 582432 157344
rect 173164 157224 173216 157276
rect 213920 157224 213972 157276
rect 324320 156816 324372 156868
rect 327356 156816 327408 156868
rect 285220 156068 285272 156120
rect 307668 156068 307720 156120
rect 271236 156000 271288 156052
rect 307484 156000 307536 156052
rect 261576 155932 261628 155984
rect 307576 155932 307628 155984
rect 352564 155932 352616 155984
rect 416780 155932 416832 155984
rect 170588 155864 170640 155916
rect 213920 155864 213972 155916
rect 252376 155864 252428 155916
rect 270684 155864 270736 155916
rect 324412 155864 324464 155916
rect 345296 155864 345348 155916
rect 497004 155864 497056 155916
rect 511264 155864 511316 155916
rect 252468 155796 252520 155848
rect 264980 155796 265032 155848
rect 324320 155796 324372 155848
rect 339684 155796 339736 155848
rect 253940 155184 253992 155236
rect 268016 155184 268068 155236
rect 274088 155184 274140 155236
rect 307392 155184 307444 155236
rect 286600 154640 286652 154692
rect 307668 154640 307720 154692
rect 264336 154572 264388 154624
rect 306564 154572 306616 154624
rect 356796 154572 356848 154624
rect 416780 154572 416832 154624
rect 252468 154504 252520 154556
rect 273352 154504 273404 154556
rect 497004 154504 497056 154556
rect 502524 154504 502576 154556
rect 252100 154436 252152 154488
rect 255412 154436 255464 154488
rect 324412 154436 324464 154488
rect 328644 154436 328696 154488
rect 497096 154436 497148 154488
rect 502616 154436 502668 154488
rect 324320 154300 324372 154352
rect 325976 154300 326028 154352
rect 256240 153824 256292 153876
rect 307300 153824 307352 153876
rect 191288 153280 191340 153332
rect 213920 153280 213972 153332
rect 301596 153280 301648 153332
rect 307668 153280 307720 153332
rect 178868 153212 178920 153264
rect 214012 153212 214064 153264
rect 268476 153212 268528 153264
rect 306932 153212 306984 153264
rect 359464 153212 359516 153264
rect 416780 153212 416832 153264
rect 252284 153144 252336 153196
rect 253940 153144 253992 153196
rect 324320 153144 324372 153196
rect 341156 153144 341208 153196
rect 497004 153144 497056 153196
rect 505192 153144 505244 153196
rect 574744 153144 574796 153196
rect 579804 153144 579856 153196
rect 252376 153076 252428 153128
rect 274732 153076 274784 153128
rect 252468 153008 252520 153060
rect 276204 153008 276256 153060
rect 299112 152532 299164 152584
rect 307668 152532 307720 152584
rect 253204 152464 253256 152516
rect 307484 152464 307536 152516
rect 173164 151920 173216 151972
rect 214012 151920 214064 151972
rect 189724 151852 189776 151904
rect 213920 151852 213972 151904
rect 257436 151784 257488 151836
rect 307116 151784 307168 151836
rect 252468 151716 252520 151768
rect 254032 151716 254084 151768
rect 324320 151716 324372 151768
rect 338304 151716 338356 151768
rect 497004 151716 497056 151768
rect 508044 151716 508096 151768
rect 324412 151648 324464 151700
rect 332600 151648 332652 151700
rect 252468 151444 252520 151496
rect 255596 151444 255648 151496
rect 252284 151240 252336 151292
rect 255504 151240 255556 151292
rect 167644 151036 167696 151088
rect 184572 151036 184624 151088
rect 293408 150560 293460 150612
rect 307668 150560 307720 150612
rect 255964 150492 256016 150544
rect 307484 150492 307536 150544
rect 176016 150424 176068 150476
rect 213920 150424 213972 150476
rect 254676 150424 254728 150476
rect 307576 150424 307628 150476
rect 331864 150424 331916 150476
rect 416780 150424 416832 150476
rect 3424 150356 3476 150408
rect 22744 150356 22796 150408
rect 184572 150356 184624 150408
rect 214012 150356 214064 150408
rect 252376 150356 252428 150408
rect 284300 150356 284352 150408
rect 324320 150356 324372 150408
rect 336740 150356 336792 150408
rect 497004 150356 497056 150408
rect 501236 150356 501288 150408
rect 209136 150288 209188 150340
rect 213920 150288 213972 150340
rect 252468 150288 252520 150340
rect 280160 150288 280212 150340
rect 252284 150220 252336 150272
rect 256792 150220 256844 150272
rect 324320 149744 324372 149796
rect 327264 149744 327316 149796
rect 281080 149676 281132 149728
rect 306656 149676 306708 149728
rect 275560 149132 275612 149184
rect 307576 149132 307628 149184
rect 267280 149064 267332 149116
rect 307668 149064 307720 149116
rect 363604 149064 363656 149116
rect 416780 149064 416832 149116
rect 211896 148996 211948 149048
rect 213920 148996 213972 149048
rect 252468 148996 252520 149048
rect 281540 148996 281592 149048
rect 324320 148996 324372 149048
rect 349252 148996 349304 149048
rect 497004 148996 497056 149048
rect 509332 148996 509384 149048
rect 252376 148928 252428 148980
rect 256700 148928 256752 148980
rect 256148 148316 256200 148368
rect 306748 148316 306800 148368
rect 182916 147636 182968 147688
rect 213920 147636 213972 147688
rect 256056 147636 256108 147688
rect 307116 147636 307168 147688
rect 374644 147636 374696 147688
rect 416780 147636 416832 147688
rect 252376 147568 252428 147620
rect 278780 147568 278832 147620
rect 324320 147568 324372 147620
rect 350540 147568 350592 147620
rect 497004 147568 497056 147620
rect 505100 147568 505152 147620
rect 252468 147500 252520 147552
rect 274640 147500 274692 147552
rect 251456 147432 251508 147484
rect 254216 147432 254268 147484
rect 325792 147024 325844 147076
rect 325700 146820 325752 146872
rect 254860 146480 254912 146532
rect 307668 146480 307720 146532
rect 276848 146412 276900 146464
rect 307576 146412 307628 146464
rect 185584 146344 185636 146396
rect 214012 146344 214064 146396
rect 257528 146344 257580 146396
rect 307668 146344 307720 146396
rect 171784 146276 171836 146328
rect 213920 146276 213972 146328
rect 303620 146276 303672 146328
rect 307484 146276 307536 146328
rect 334716 146276 334768 146328
rect 416780 146276 416832 146328
rect 252468 146208 252520 146260
rect 271880 146208 271932 146260
rect 324320 146208 324372 146260
rect 353392 146208 353444 146260
rect 525800 146208 525852 146260
rect 580264 146208 580316 146260
rect 252376 146140 252428 146192
rect 267832 146140 267884 146192
rect 324412 146140 324464 146192
rect 346492 146140 346544 146192
rect 251180 146072 251232 146124
rect 253480 146072 253532 146124
rect 213368 145664 213420 145716
rect 215024 145664 215076 145716
rect 253388 145528 253440 145580
rect 306840 145528 306892 145580
rect 502984 145528 503036 145580
rect 525800 145528 525852 145580
rect 292120 144916 292172 144968
rect 306564 144916 306616 144968
rect 497004 144916 497056 144968
rect 502340 144916 502392 144968
rect 252468 144848 252520 144900
rect 260840 144848 260892 144900
rect 324320 144848 324372 144900
rect 335360 144848 335412 144900
rect 252100 144304 252152 144356
rect 268568 144304 268620 144356
rect 267188 144236 267240 144288
rect 307392 144236 307444 144288
rect 250720 144168 250772 144220
rect 303620 144168 303672 144220
rect 508044 144168 508096 144220
rect 509148 144168 509200 144220
rect 512092 144168 512144 144220
rect 307024 144100 307076 144152
rect 307392 144100 307444 144152
rect 170496 143624 170548 143676
rect 213920 143624 213972 143676
rect 302976 143624 303028 143676
rect 306564 143624 306616 143676
rect 169024 143556 169076 143608
rect 214012 143556 214064 143608
rect 290648 143556 290700 143608
rect 307668 143556 307720 143608
rect 358084 143556 358136 143608
rect 416780 143556 416832 143608
rect 497096 143556 497148 143608
rect 508044 143556 508096 143608
rect 252468 143488 252520 143540
rect 270592 143488 270644 143540
rect 497004 143488 497056 143540
rect 513380 143488 513432 143540
rect 252376 143420 252428 143472
rect 269120 143420 269172 143472
rect 324320 143420 324372 143472
rect 343732 143420 343784 143472
rect 513380 143352 513432 143404
rect 515404 143352 515456 143404
rect 167644 142808 167696 142860
rect 213460 142808 213512 142860
rect 274180 142808 274232 142860
rect 307484 142808 307536 142860
rect 289360 142196 289412 142248
rect 307668 142196 307720 142248
rect 181536 142128 181588 142180
rect 213920 142128 213972 142180
rect 254768 142128 254820 142180
rect 307576 142128 307628 142180
rect 345664 142128 345716 142180
rect 416780 142128 416832 142180
rect 252468 142060 252520 142112
rect 262496 142060 262548 142112
rect 324320 142060 324372 142112
rect 356060 142060 356112 142112
rect 497004 142060 497056 142112
rect 507952 142060 508004 142112
rect 251180 141516 251232 141568
rect 253296 141516 253348 141568
rect 287980 141448 288032 141500
rect 306564 141448 306616 141500
rect 252008 141380 252060 141432
rect 294696 141380 294748 141432
rect 496820 141380 496872 141432
rect 503260 141380 503312 141432
rect 301872 140904 301924 140956
rect 306932 140904 306984 140956
rect 209136 140836 209188 140888
rect 214012 140836 214064 140888
rect 303252 140836 303304 140888
rect 307576 140836 307628 140888
rect 174544 140768 174596 140820
rect 213920 140768 213972 140820
rect 262956 140768 263008 140820
rect 307668 140768 307720 140820
rect 333428 140768 333480 140820
rect 416780 140768 416832 140820
rect 507952 140768 508004 140820
rect 511264 140768 511316 140820
rect 252468 140700 252520 140752
rect 277492 140700 277544 140752
rect 324320 140700 324372 140752
rect 328460 140700 328512 140752
rect 496820 140700 496872 140752
rect 502984 140700 503036 140752
rect 252376 140632 252428 140684
rect 276020 140632 276072 140684
rect 177396 140020 177448 140072
rect 214656 140020 214708 140072
rect 503260 140020 503312 140072
rect 580172 140020 580224 140072
rect 251916 139952 251968 140004
rect 259000 139952 259052 140004
rect 271420 139476 271472 139528
rect 306564 139476 306616 139528
rect 184388 139408 184440 139460
rect 213920 139408 213972 139460
rect 254584 139408 254636 139460
rect 307668 139408 307720 139460
rect 411904 139408 411956 139460
rect 416780 139408 416832 139460
rect 252468 139340 252520 139392
rect 263600 139340 263652 139392
rect 324412 139340 324464 139392
rect 339500 139340 339552 139392
rect 496820 139340 496872 139392
rect 520924 139340 520976 139392
rect 324320 139272 324372 139324
rect 334072 139272 334124 139324
rect 294880 138116 294932 138168
rect 306932 138116 306984 138168
rect 195336 138048 195388 138100
rect 213920 138048 213972 138100
rect 253296 138048 253348 138100
rect 307668 138048 307720 138100
rect 174636 137980 174688 138032
rect 214012 137980 214064 138032
rect 249064 137980 249116 138032
rect 306564 137980 306616 138032
rect 3240 137912 3292 137964
rect 15844 137912 15896 137964
rect 252468 137912 252520 137964
rect 277400 137912 277452 137964
rect 324320 137912 324372 137964
rect 332692 137912 332744 137964
rect 496820 137912 496872 137964
rect 547880 137912 547932 137964
rect 252192 137232 252244 137284
rect 260288 137232 260340 137284
rect 210424 136688 210476 136740
rect 214012 136688 214064 136740
rect 260104 136688 260156 136740
rect 307116 136688 307168 136740
rect 166264 136620 166316 136672
rect 213920 136620 213972 136672
rect 250628 136620 250680 136672
rect 307668 136620 307720 136672
rect 376024 136620 376076 136672
rect 416780 136620 416832 136672
rect 252284 136552 252336 136604
rect 302884 136552 302936 136604
rect 324320 136552 324372 136604
rect 329932 136552 329984 136604
rect 496820 136552 496872 136604
rect 538220 136552 538272 136604
rect 252468 136484 252520 136536
rect 297456 136484 297508 136536
rect 497004 136484 497056 136536
rect 506480 136484 506532 136536
rect 252376 136416 252428 136468
rect 267004 136416 267056 136468
rect 268568 135872 268620 135924
rect 307024 135872 307076 135924
rect 304264 135396 304316 135448
rect 307484 135396 307536 135448
rect 206468 135328 206520 135380
rect 213920 135328 213972 135380
rect 298836 135328 298888 135380
rect 307668 135328 307720 135380
rect 171968 135260 172020 135312
rect 214012 135260 214064 135312
rect 250444 135260 250496 135312
rect 306564 135260 306616 135312
rect 403624 135260 403676 135312
rect 416780 135260 416832 135312
rect 252468 135192 252520 135244
rect 285036 135192 285088 135244
rect 336096 135192 336148 135244
rect 417332 135192 417384 135244
rect 496820 135192 496872 135244
rect 525064 135192 525116 135244
rect 252376 135124 252428 135176
rect 271144 135124 271196 135176
rect 297456 134512 297508 134564
rect 307208 134512 307260 134564
rect 282460 133968 282512 134020
rect 307576 133968 307628 134020
rect 175924 133900 175976 133952
rect 213920 133900 213972 133952
rect 275376 133900 275428 133952
rect 307668 133900 307720 133952
rect 252284 133832 252336 133884
rect 304448 133832 304500 133884
rect 324320 133832 324372 133884
rect 346400 133832 346452 133884
rect 378784 133832 378836 133884
rect 419356 133832 419408 133884
rect 252376 133764 252428 133816
rect 286416 133764 286468 133816
rect 252468 133696 252520 133748
rect 264244 133696 264296 133748
rect 259000 133152 259052 133204
rect 307392 133152 307444 133204
rect 286508 132540 286560 132592
rect 306932 132540 306984 132592
rect 187148 132472 187200 132524
rect 213920 132472 213972 132524
rect 285128 132472 285180 132524
rect 306564 132472 306616 132524
rect 324964 132472 325016 132524
rect 327080 132472 327132 132524
rect 252376 132404 252428 132456
rect 289268 132404 289320 132456
rect 324412 132404 324464 132456
rect 357532 132404 357584 132456
rect 410524 132404 410576 132456
rect 417608 132404 417660 132456
rect 252468 132336 252520 132388
rect 273996 132336 274048 132388
rect 324320 132336 324372 132388
rect 342352 132336 342404 132388
rect 294696 131248 294748 131300
rect 307484 131248 307536 131300
rect 289084 131180 289136 131232
rect 307576 131180 307628 131232
rect 173256 131112 173308 131164
rect 213920 131112 213972 131164
rect 278136 131112 278188 131164
rect 307668 131112 307720 131164
rect 252376 131044 252428 131096
rect 290556 131044 290608 131096
rect 324320 131044 324372 131096
rect 349160 131044 349212 131096
rect 252284 130976 252336 131028
rect 267096 130976 267148 131028
rect 324412 130976 324464 131028
rect 328736 130976 328788 131028
rect 252468 130908 252520 130960
rect 262864 130908 262916 130960
rect 202236 130364 202288 130416
rect 214748 130364 214800 130416
rect 267372 130364 267424 130416
rect 305736 130364 305788 130416
rect 291936 129888 291988 129940
rect 307668 129888 307720 129940
rect 290464 129820 290516 129872
rect 307484 129820 307536 129872
rect 171876 129752 171928 129804
rect 213920 129752 213972 129804
rect 273996 129752 274048 129804
rect 307576 129752 307628 129804
rect 252468 129684 252520 129736
rect 278228 129684 278280 129736
rect 324320 129684 324372 129736
rect 352012 129684 352064 129736
rect 408408 129684 408460 129736
rect 416780 129684 416832 129736
rect 496820 129684 496872 129736
rect 510620 129684 510672 129736
rect 252376 129616 252428 129668
rect 265808 129616 265860 129668
rect 324412 129616 324464 129668
rect 331220 129616 331272 129668
rect 496912 129616 496964 129668
rect 506664 129616 506716 129668
rect 252284 129548 252336 129600
rect 257344 129548 257396 129600
rect 276756 128392 276808 128444
rect 306932 128392 306984 128444
rect 188528 128324 188580 128376
rect 213920 128324 213972 128376
rect 264244 128324 264296 128376
rect 307668 128324 307720 128376
rect 252468 128256 252520 128308
rect 287888 128256 287940 128308
rect 324320 128256 324372 128308
rect 331312 128256 331364 128308
rect 377404 128256 377456 128308
rect 419632 128256 419684 128308
rect 419816 128256 419868 128308
rect 252284 128188 252336 128240
rect 269764 128188 269816 128240
rect 324412 128188 324464 128240
rect 330116 128188 330168 128240
rect 252376 128120 252428 128172
rect 258724 128120 258776 128172
rect 536104 127576 536156 127628
rect 580172 127576 580224 127628
rect 287796 127100 287848 127152
rect 307668 127100 307720 127152
rect 285036 127032 285088 127084
rect 307484 127032 307536 127084
rect 59268 126964 59320 127016
rect 65524 126964 65576 127016
rect 180156 126964 180208 127016
rect 213920 126964 213972 127016
rect 269856 126964 269908 127016
rect 307576 126964 307628 127016
rect 496912 126964 496964 127016
rect 498292 126964 498344 127016
rect 252284 126896 252336 126948
rect 283748 126896 283800 126948
rect 406384 126896 406436 126948
rect 418528 126896 418580 126948
rect 419264 126896 419316 126948
rect 496820 126896 496872 126948
rect 514760 126896 514812 126948
rect 252468 126828 252520 126880
rect 268384 126828 268436 126880
rect 252376 126760 252428 126812
rect 264428 126760 264480 126812
rect 202328 125672 202380 125724
rect 213920 125672 213972 125724
rect 283656 125672 283708 125724
rect 307576 125672 307628 125724
rect 169116 125604 169168 125656
rect 214012 125604 214064 125656
rect 276940 125604 276992 125656
rect 307668 125604 307720 125656
rect 252468 125536 252520 125588
rect 297456 125536 297508 125588
rect 324320 125536 324372 125588
rect 328552 125536 328604 125588
rect 342996 125536 343048 125588
rect 418528 125536 418580 125588
rect 419448 125536 419500 125588
rect 496820 125536 496872 125588
rect 521660 125536 521712 125588
rect 324412 125468 324464 125520
rect 345112 125468 345164 125520
rect 252100 124924 252152 124976
rect 263048 124924 263100 124976
rect 251824 124856 251876 124908
rect 302976 124856 303028 124908
rect 303068 124380 303120 124432
rect 307668 124380 307720 124432
rect 297548 124312 297600 124364
rect 307576 124312 307628 124364
rect 199476 124244 199528 124296
rect 213920 124244 213972 124296
rect 286416 124244 286468 124296
rect 307484 124244 307536 124296
rect 170588 124176 170640 124228
rect 214012 124176 214064 124228
rect 278228 124176 278280 124228
rect 307668 124176 307720 124228
rect 252376 124108 252428 124160
rect 304356 124108 304408 124160
rect 324320 124108 324372 124160
rect 353300 124108 353352 124160
rect 496820 124108 496872 124160
rect 499580 124108 499632 124160
rect 252468 124040 252520 124092
rect 298928 124040 298980 124092
rect 252284 123972 252336 124024
rect 261668 123972 261720 124024
rect 178960 122884 179012 122936
rect 213920 122884 213972 122936
rect 298744 122884 298796 122936
rect 307668 122884 307720 122936
rect 167828 122816 167880 122868
rect 214012 122816 214064 122868
rect 297640 122816 297692 122868
rect 307576 122816 307628 122868
rect 252468 122748 252520 122800
rect 296076 122748 296128 122800
rect 324320 122748 324372 122800
rect 342260 122748 342312 122800
rect 399484 122748 399536 122800
rect 419540 122748 419592 122800
rect 252376 122680 252428 122732
rect 272708 122680 272760 122732
rect 252284 122612 252336 122664
rect 261484 122612 261536 122664
rect 170404 122068 170456 122120
rect 196716 122068 196768 122120
rect 300400 121592 300452 121644
rect 307576 121592 307628 121644
rect 198188 121524 198240 121576
rect 214012 121524 214064 121576
rect 296260 121524 296312 121576
rect 307668 121524 307720 121576
rect 180248 121456 180300 121508
rect 213920 121456 213972 121508
rect 272616 121456 272668 121508
rect 306748 121456 306800 121508
rect 252468 121388 252520 121440
rect 256240 121388 256292 121440
rect 324320 121388 324372 121440
rect 352104 121388 352156 121440
rect 496820 121388 496872 121440
rect 517520 121388 517572 121440
rect 324412 121320 324464 121372
rect 347780 121320 347832 121372
rect 258724 120232 258776 120284
rect 307300 120232 307352 120284
rect 210516 120164 210568 120216
rect 214012 120164 214064 120216
rect 250536 120164 250588 120216
rect 176108 120096 176160 120148
rect 213920 120096 213972 120148
rect 252008 120096 252060 120148
rect 254860 120096 254912 120148
rect 257344 120164 257396 120216
rect 307668 120164 307720 120216
rect 307576 120096 307628 120148
rect 252284 120028 252336 120080
rect 292028 120028 292080 120080
rect 400864 120028 400916 120080
rect 416780 120028 416832 120080
rect 252468 119960 252520 120012
rect 265716 119960 265768 120012
rect 252376 119824 252428 119876
rect 260196 119824 260248 119876
rect 496820 119756 496872 119808
rect 499764 119756 499816 119808
rect 271512 119348 271564 119400
rect 307208 119348 307260 119400
rect 193956 118804 194008 118856
rect 214012 118804 214064 118856
rect 279608 118804 279660 118856
rect 306564 118804 306616 118856
rect 185676 118736 185728 118788
rect 213920 118736 213972 118788
rect 299020 118736 299072 118788
rect 307668 118736 307720 118788
rect 177488 118668 177540 118720
rect 214104 118668 214156 118720
rect 252376 118600 252428 118652
rect 300216 118600 300268 118652
rect 324320 118600 324372 118652
rect 354680 118600 354732 118652
rect 414664 118600 414716 118652
rect 416964 118600 417016 118652
rect 496820 118600 496872 118652
rect 512184 118600 512236 118652
rect 252284 118532 252336 118584
rect 274088 118532 274140 118584
rect 324412 118532 324464 118584
rect 347872 118532 347924 118584
rect 496912 118532 496964 118584
rect 509240 118532 509292 118584
rect 252468 117648 252520 117700
rect 258816 117648 258868 117700
rect 265716 117512 265768 117564
rect 307668 117512 307720 117564
rect 196900 117376 196952 117428
rect 214012 117376 214064 117428
rect 283748 117376 283800 117428
rect 307576 117376 307628 117428
rect 170404 117308 170456 117360
rect 213920 117308 213972 117360
rect 304356 117308 304408 117360
rect 307300 117308 307352 117360
rect 252468 117240 252520 117292
rect 271236 117240 271288 117292
rect 324320 117240 324372 117292
rect 340972 117240 341024 117292
rect 252376 117172 252428 117224
rect 261576 117172 261628 117224
rect 251916 116560 251968 116612
rect 267280 116560 267332 116612
rect 293316 116084 293368 116136
rect 307668 116084 307720 116136
rect 174820 116016 174872 116068
rect 214012 116016 214064 116068
rect 271144 116016 271196 116068
rect 307576 116016 307628 116068
rect 169208 115948 169260 116000
rect 213920 115948 213972 116000
rect 267004 115948 267056 116000
rect 307484 115948 307536 116000
rect 252468 115880 252520 115932
rect 285220 115880 285272 115932
rect 324320 115880 324372 115932
rect 350632 115880 350684 115932
rect 496820 115880 496872 115932
rect 503720 115880 503772 115932
rect 252376 115812 252428 115864
rect 264336 115812 264388 115864
rect 324412 115812 324464 115864
rect 343640 115812 343692 115864
rect 252284 115200 252336 115252
rect 268476 115200 268528 115252
rect 296076 114656 296128 114708
rect 307576 114656 307628 114708
rect 211896 114588 211948 114640
rect 214012 114588 214064 114640
rect 280988 114588 281040 114640
rect 307668 114588 307720 114640
rect 167736 114520 167788 114572
rect 213920 114520 213972 114572
rect 268384 114520 268436 114572
rect 307300 114520 307352 114572
rect 252468 114452 252520 114504
rect 286600 114452 286652 114504
rect 333336 114452 333388 114504
rect 416780 114452 416832 114504
rect 496820 114452 496872 114504
rect 499672 114452 499724 114504
rect 324320 114384 324372 114436
rect 349344 114384 349396 114436
rect 252376 113772 252428 113824
rect 301596 113772 301648 113824
rect 195428 113228 195480 113280
rect 214012 113228 214064 113280
rect 301688 113228 301740 113280
rect 306564 113228 306616 113280
rect 167920 113160 167972 113212
rect 213920 113160 213972 113212
rect 290556 113160 290608 113212
rect 307668 113160 307720 113212
rect 252468 113092 252520 113144
rect 299112 113092 299164 113144
rect 324320 113092 324372 113144
rect 338120 113092 338172 113144
rect 496820 113092 496872 113144
rect 501052 113092 501104 113144
rect 252284 113024 252336 113076
rect 256148 113024 256200 113076
rect 337476 113024 337528 113076
rect 416780 113024 416832 113076
rect 252284 112412 252336 112464
rect 276848 112412 276900 112464
rect 298928 111936 298980 111988
rect 307668 111936 307720 111988
rect 297456 111868 297508 111920
rect 307576 111868 307628 111920
rect 166356 111800 166408 111852
rect 213920 111800 213972 111852
rect 269764 111800 269816 111852
rect 307484 111800 307536 111852
rect 168012 111732 168064 111784
rect 176016 111732 176068 111784
rect 251180 111732 251232 111784
rect 253388 111732 253440 111784
rect 367744 111732 367796 111784
rect 416780 111732 416832 111784
rect 496912 111732 496964 111784
rect 503812 111732 503864 111784
rect 252376 111664 252428 111716
rect 257436 111664 257488 111716
rect 496820 111664 496872 111716
rect 502432 111664 502484 111716
rect 252468 111596 252520 111648
rect 281080 111596 281132 111648
rect 3700 111052 3752 111104
rect 4068 111052 4120 111104
rect 14464 111052 14516 111104
rect 294788 110576 294840 110628
rect 306748 110576 306800 110628
rect 184480 110508 184532 110560
rect 213920 110508 213972 110560
rect 292028 110508 292080 110560
rect 307300 110508 307352 110560
rect 169300 110440 169352 110492
rect 214012 110440 214064 110492
rect 279516 110440 279568 110492
rect 307668 110440 307720 110492
rect 168104 110372 168156 110424
rect 213368 110372 213420 110424
rect 251732 110372 251784 110424
rect 254676 110372 254728 110424
rect 324320 110372 324372 110424
rect 341064 110372 341116 110424
rect 496820 110372 496872 110424
rect 506572 110372 506624 110424
rect 252468 110304 252520 110356
rect 255964 110304 256016 110356
rect 302884 109148 302936 109200
rect 307576 109148 307628 109200
rect 257436 109080 257488 109132
rect 306932 109080 306984 109132
rect 172060 109012 172112 109064
rect 213920 109012 213972 109064
rect 253204 109012 253256 109064
rect 307668 109012 307720 109064
rect 252376 108944 252428 108996
rect 278320 108944 278372 108996
rect 324320 108944 324372 108996
rect 345204 108944 345256 108996
rect 252468 108876 252520 108928
rect 275560 108876 275612 108928
rect 268476 107856 268528 107908
rect 307484 107856 307536 107908
rect 174728 107720 174780 107772
rect 214012 107720 214064 107772
rect 275468 107720 275520 107772
rect 307668 107720 307720 107772
rect 170680 107652 170732 107704
rect 213920 107652 213972 107704
rect 300308 107652 300360 107704
rect 307576 107652 307628 107704
rect 252468 107584 252520 107636
rect 267188 107584 267240 107636
rect 413284 107584 413336 107636
rect 416780 107584 416832 107636
rect 252376 107516 252428 107568
rect 256056 107516 256108 107568
rect 252468 106904 252520 106956
rect 259000 106904 259052 106956
rect 301596 106428 301648 106480
rect 307668 106428 307720 106480
rect 176016 106360 176068 106412
rect 213920 106360 213972 106412
rect 264336 106360 264388 106412
rect 307484 106360 307536 106412
rect 167644 106292 167696 106344
rect 214012 106292 214064 106344
rect 256148 106292 256200 106344
rect 306748 106292 306800 106344
rect 371884 106224 371936 106276
rect 416780 106224 416832 106276
rect 324320 105816 324372 105868
rect 327172 105816 327224 105868
rect 251364 105612 251416 105664
rect 262956 105612 263008 105664
rect 252376 105544 252428 105596
rect 292120 105544 292172 105596
rect 203616 105000 203668 105052
rect 213920 105000 213972 105052
rect 303160 105000 303212 105052
rect 307576 105000 307628 105052
rect 188620 104932 188672 104984
rect 214012 104932 214064 104984
rect 282368 104932 282420 104984
rect 307668 104932 307720 104984
rect 173440 104864 173492 104916
rect 214104 104864 214156 104916
rect 261484 104864 261536 104916
rect 306748 104864 306800 104916
rect 252468 104796 252520 104848
rect 271512 104796 271564 104848
rect 395344 104796 395396 104848
rect 416780 104796 416832 104848
rect 252284 104728 252336 104780
rect 257528 104728 257580 104780
rect 330484 104116 330536 104168
rect 403624 104116 403676 104168
rect 286600 103640 286652 103692
rect 307484 103640 307536 103692
rect 271328 103572 271380 103624
rect 306932 103572 306984 103624
rect 206560 103504 206612 103556
rect 213920 103504 213972 103556
rect 255964 103504 256016 103556
rect 306748 103504 306800 103556
rect 252376 103436 252428 103488
rect 274180 103436 274232 103488
rect 354036 103436 354088 103488
rect 416780 103436 416832 103488
rect 251732 102824 251784 102876
rect 254768 102824 254820 102876
rect 495440 102824 495492 102876
rect 495624 102824 495676 102876
rect 173348 102756 173400 102808
rect 214656 102756 214708 102808
rect 252468 102552 252520 102604
rect 258908 102552 258960 102604
rect 289268 102280 289320 102332
rect 306564 102280 306616 102332
rect 274088 102212 274140 102264
rect 307668 102212 307720 102264
rect 209228 102144 209280 102196
rect 213920 102144 213972 102196
rect 258816 102144 258868 102196
rect 307576 102144 307628 102196
rect 252468 102076 252520 102128
rect 290648 102076 290700 102128
rect 382924 102076 382976 102128
rect 416780 102076 416832 102128
rect 252376 102008 252428 102060
rect 287980 102008 288032 102060
rect 252192 101396 252244 101448
rect 271420 101396 271472 101448
rect 326344 101396 326396 101448
rect 376024 101396 376076 101448
rect 511264 101396 511316 101448
rect 580172 101396 580224 101448
rect 271236 100920 271288 100972
rect 307668 100920 307720 100972
rect 300216 100852 300268 100904
rect 306564 100852 306616 100904
rect 287888 100784 287940 100836
rect 307576 100784 307628 100836
rect 177580 100716 177632 100768
rect 213920 100716 213972 100768
rect 304448 100716 304500 100768
rect 307484 100716 307536 100768
rect 252284 100648 252336 100700
rect 301872 100648 301924 100700
rect 419724 100648 419776 100700
rect 580264 100648 580316 100700
rect 252468 100580 252520 100632
rect 289360 100580 289412 100632
rect 389824 100580 389876 100632
rect 496820 100580 496872 100632
rect 252376 100512 252428 100564
rect 268568 100512 268620 100564
rect 323584 99968 323636 100020
rect 411904 99968 411956 100020
rect 301780 99492 301832 99544
rect 307484 99492 307536 99544
rect 296168 99424 296220 99476
rect 307576 99424 307628 99476
rect 211988 99356 212040 99408
rect 214288 99356 214340 99408
rect 285220 99356 285272 99408
rect 307668 99356 307720 99408
rect 252376 99288 252428 99340
rect 303252 99288 303304 99340
rect 388444 99288 388496 99340
rect 497096 99288 497148 99340
rect 252468 99220 252520 99272
rect 267372 99220 267424 99272
rect 393964 99220 394016 99272
rect 497004 99220 497056 99272
rect 396724 99152 396776 99204
rect 494060 99152 494112 99204
rect 302976 98132 303028 98184
rect 307668 98132 307720 98184
rect 199568 98064 199620 98116
rect 213920 98064 213972 98116
rect 281080 98064 281132 98116
rect 307576 98064 307628 98116
rect 166448 97996 166500 98048
rect 214012 97996 214064 98048
rect 249248 97996 249300 98048
rect 307300 97996 307352 98048
rect 370504 97928 370556 97980
rect 495440 97928 495492 97980
rect 392584 97860 392636 97912
rect 496912 97860 496964 97912
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 421012 97316 421064 97368
rect 426532 97316 426584 97368
rect 421564 97248 421616 97300
rect 456524 97248 456576 97300
rect 461584 97248 461636 97300
rect 474556 97248 474608 97300
rect 475384 97248 475436 97300
rect 492496 97248 492548 97300
rect 414664 96908 414716 96960
rect 420552 96908 420604 96960
rect 439504 96908 439556 96960
rect 440884 96908 440936 96960
rect 454040 96908 454092 96960
rect 455052 96908 455104 96960
rect 481640 96908 481692 96960
rect 482652 96908 482704 96960
rect 486424 96908 486476 96960
rect 487712 96908 487764 96960
rect 457444 96772 457496 96824
rect 460112 96772 460164 96824
rect 278320 96704 278372 96756
rect 307668 96704 307720 96756
rect 267096 96636 267148 96688
rect 307576 96636 307628 96688
rect 191196 96568 191248 96620
rect 323032 96568 323084 96620
rect 381544 96568 381596 96620
rect 495624 96568 495676 96620
rect 300124 96500 300176 96552
rect 321468 96500 321520 96552
rect 351920 96500 351972 96552
rect 421012 96500 421064 96552
rect 166908 95888 166960 95940
rect 214104 95888 214156 95940
rect 324320 95888 324372 95940
rect 351920 95888 351972 95940
rect 419172 95888 419224 95940
rect 580264 95888 580316 95940
rect 164884 95616 164936 95668
rect 165620 95616 165672 95668
rect 251824 95208 251876 95260
rect 307668 95208 307720 95260
rect 178776 95140 178828 95192
rect 321560 95140 321612 95192
rect 337384 95140 337436 95192
rect 498476 95140 498528 95192
rect 181444 95072 181496 95124
rect 321376 95072 321428 95124
rect 193864 95004 193916 95056
rect 322940 95004 322992 95056
rect 199384 94936 199436 94988
rect 321652 94936 321704 94988
rect 206376 94868 206428 94920
rect 321836 94868 321888 94920
rect 336740 94664 336792 94716
rect 337384 94664 337436 94716
rect 320824 94460 320876 94512
rect 427728 94460 427780 94512
rect 152096 94120 152148 94172
rect 189724 94120 189776 94172
rect 126520 94052 126572 94104
rect 169116 94052 169168 94104
rect 126704 93984 126756 94036
rect 181536 93984 181588 94036
rect 112352 93916 112404 93968
rect 185676 93916 185728 93968
rect 96160 93848 96212 93900
rect 172060 93848 172112 93900
rect 133144 93440 133196 93492
rect 171784 93440 171836 93492
rect 151728 93372 151780 93424
rect 191288 93372 191340 93424
rect 121736 93304 121788 93356
rect 167828 93304 167880 93356
rect 116768 93236 116820 93288
rect 166264 93236 166316 93288
rect 109224 93168 109276 93220
rect 174820 93168 174872 93220
rect 100944 93100 100996 93152
rect 188528 93100 188580 93152
rect 232504 93100 232556 93152
rect 278228 93100 278280 93152
rect 88984 92420 89036 92472
rect 166908 92420 166960 92472
rect 187056 92420 187108 92472
rect 321744 92420 321796 92472
rect 118056 92352 118108 92404
rect 195336 92352 195388 92404
rect 196808 92352 196860 92404
rect 321928 92352 321980 92404
rect 115480 92284 115532 92336
rect 210424 92284 210476 92336
rect 114468 92216 114520 92268
rect 202236 92216 202288 92268
rect 103336 92148 103388 92200
rect 173348 92148 173400 92200
rect 132408 92080 132460 92132
rect 177396 92080 177448 92132
rect 238024 91808 238076 91860
rect 251180 91808 251232 91860
rect 200764 91740 200816 91792
rect 253388 91740 253440 91792
rect 277400 91740 277452 91792
rect 481732 91740 481784 91792
rect 74816 91128 74868 91180
rect 88984 91128 89036 91180
rect 97540 91128 97592 91180
rect 116124 91128 116176 91180
rect 85856 91060 85908 91112
rect 122104 91060 122156 91112
rect 88064 90992 88116 91044
rect 211988 90992 212040 91044
rect 252468 90992 252520 91044
rect 420920 90992 420972 91044
rect 98828 90924 98880 90976
rect 184480 90924 184532 90976
rect 114928 90856 114980 90908
rect 193956 90856 194008 90908
rect 103244 90788 103296 90840
rect 167920 90788 167972 90840
rect 151544 90720 151596 90772
rect 178868 90720 178920 90772
rect 151636 90652 151688 90704
rect 173164 90652 173216 90704
rect 311900 90380 311952 90432
rect 358084 90380 358136 90432
rect 352656 90312 352708 90364
rect 456800 90312 456852 90364
rect 251916 89700 251968 89752
rect 252468 89700 252520 89752
rect 67640 89632 67692 89684
rect 214840 89632 214892 89684
rect 348424 89632 348476 89684
rect 501144 89632 501196 89684
rect 110144 89564 110196 89616
rect 170404 89564 170456 89616
rect 182824 89564 182876 89616
rect 324412 89564 324464 89616
rect 90732 89496 90784 89548
rect 188620 89496 188672 89548
rect 122840 89428 122892 89480
rect 199476 89428 199528 89480
rect 119804 89360 119856 89412
rect 174636 89360 174688 89412
rect 136456 89292 136508 89344
rect 182916 89292 182968 89344
rect 347780 89224 347832 89276
rect 348424 89224 348476 89276
rect 295984 88952 296036 89004
rect 315304 88952 315356 89004
rect 316684 88952 316736 89004
rect 345664 88952 345716 89004
rect 67732 88272 67784 88324
rect 214656 88272 214708 88324
rect 116124 88204 116176 88256
rect 214748 88204 214800 88256
rect 104256 88136 104308 88188
rect 195428 88136 195480 88188
rect 120724 88068 120776 88120
rect 178960 88068 179012 88120
rect 129464 88000 129516 88052
rect 169024 88000 169076 88052
rect 308496 87660 308548 87712
rect 324964 87660 325016 87712
rect 213184 87592 213236 87644
rect 276020 87592 276072 87644
rect 278044 87592 278096 87644
rect 331956 87592 332008 87644
rect 342352 87592 342404 87644
rect 458180 87592 458232 87644
rect 276020 86980 276072 87032
rect 276848 86980 276900 87032
rect 277400 86980 277452 87032
rect 88984 86912 89036 86964
rect 214564 86912 214616 86964
rect 339500 86912 339552 86964
rect 340144 86912 340196 86964
rect 457444 86912 457496 86964
rect 504456 86912 504508 86964
rect 580172 86912 580224 86964
rect 126520 86844 126572 86896
rect 213276 86844 213328 86896
rect 86776 86776 86828 86828
rect 166448 86776 166500 86828
rect 100576 86708 100628 86760
rect 166356 86708 166408 86760
rect 107936 86640 107988 86692
rect 169208 86640 169260 86692
rect 117136 86572 117188 86624
rect 176108 86572 176160 86624
rect 211804 86232 211856 86284
rect 322204 86232 322256 86284
rect 3148 85484 3200 85536
rect 17224 85484 17276 85536
rect 65984 85484 66036 85536
rect 216680 85484 216732 85536
rect 101864 85416 101916 85468
rect 213460 85416 213512 85468
rect 113364 85348 113416 85400
rect 177488 85348 177540 85400
rect 114376 85280 114428 85332
rect 171968 85280 172020 85332
rect 124036 85212 124088 85264
rect 170588 85212 170640 85264
rect 319444 84804 319496 84856
rect 333428 84804 333480 84856
rect 336096 84804 336148 84856
rect 460940 84804 460992 84856
rect 107476 84124 107528 84176
rect 187148 84124 187200 84176
rect 100668 84056 100720 84108
rect 169300 84056 169352 84108
rect 106096 83988 106148 84040
rect 167736 83988 167788 84040
rect 118608 83920 118660 83972
rect 180248 83920 180300 83972
rect 124128 83852 124180 83904
rect 174544 83852 174596 83904
rect 308496 83580 308548 83632
rect 334716 83580 334768 83632
rect 207664 83512 207716 83564
rect 331220 83512 331272 83564
rect 178776 83444 178828 83496
rect 307116 83444 307168 83496
rect 463792 83444 463844 83496
rect 107568 82764 107620 82816
rect 211896 82764 211948 82816
rect 119988 82696 120040 82748
rect 198188 82696 198240 82748
rect 95056 82628 95108 82680
rect 170680 82628 170732 82680
rect 104808 82560 104860 82612
rect 173256 82560 173308 82612
rect 135168 82492 135220 82544
rect 185584 82492 185636 82544
rect 206284 82084 206336 82136
rect 261576 82084 261628 82136
rect 289176 82084 289228 82136
rect 317420 82084 317472 82136
rect 466460 82084 466512 82136
rect 111708 81336 111760 81388
rect 196900 81336 196952 81388
rect 125416 81268 125468 81320
rect 209136 81268 209188 81320
rect 97816 81200 97868 81252
rect 180156 81200 180208 81252
rect 93768 81132 93820 81184
rect 167644 81132 167696 81184
rect 209044 80656 209096 80708
rect 278044 80656 278096 80708
rect 309876 80656 309928 80708
rect 470600 80656 470652 80708
rect 204904 79976 204956 80028
rect 325700 79976 325752 80028
rect 326344 79976 326396 80028
rect 92388 79908 92440 79960
rect 176016 79908 176068 79960
rect 125508 79840 125560 79892
rect 202328 79840 202380 79892
rect 113088 79772 113140 79824
rect 206468 79772 206520 79824
rect 202144 79364 202196 79416
rect 246304 79364 246356 79416
rect 184204 79296 184256 79348
rect 303620 79296 303672 79348
rect 471980 79296 472032 79348
rect 115756 78616 115808 78668
rect 210516 78616 210568 78668
rect 95148 78548 95200 78600
rect 174728 78548 174780 78600
rect 102048 78480 102100 78532
rect 171876 78480 171928 78532
rect 121368 78412 121420 78464
rect 184388 78412 184440 78464
rect 249156 78004 249208 78056
rect 355324 78004 355376 78056
rect 310520 77936 310572 77988
rect 469220 77936 469272 77988
rect 85488 77188 85540 77240
rect 177580 77188 177632 77240
rect 297364 77188 297416 77240
rect 329840 77188 329892 77240
rect 330484 77188 330536 77240
rect 110328 77120 110380 77172
rect 175924 77120 175976 77172
rect 177304 76508 177356 76560
rect 254676 76508 254728 76560
rect 324964 76508 325016 76560
rect 463884 76508 463936 76560
rect 122104 75828 122156 75880
rect 199568 75828 199620 75880
rect 93860 75216 93912 75268
rect 300400 75216 300452 75268
rect 69020 75148 69072 75200
rect 299020 75148 299072 75200
rect 300124 75148 300176 75200
rect 473360 75148 473412 75200
rect 51724 74468 51776 74520
rect 502340 74468 502392 74520
rect 104900 73856 104952 73908
rect 246488 73856 246540 73908
rect 102140 73788 102192 73840
rect 297640 73788 297692 73840
rect 63132 73108 63184 73160
rect 335360 73108 335412 73160
rect 336096 73108 336148 73160
rect 419356 73108 419408 73160
rect 579988 73108 580040 73160
rect 338764 73040 338816 73092
rect 422300 73040 422352 73092
rect 33140 72428 33192 72480
rect 304448 72428 304500 72480
rect 338120 71748 338172 71800
rect 338764 71748 338816 71800
rect 3424 71612 3476 71664
rect 7564 71612 7616 71664
rect 297364 71136 297416 71188
rect 461584 71136 461636 71188
rect 115940 71068 115992 71120
rect 297548 71068 297600 71120
rect 89720 71000 89772 71052
rect 305920 71000 305972 71052
rect 293224 69708 293276 69760
rect 474740 69708 474792 69760
rect 86960 69640 87012 69692
rect 296260 69640 296312 69692
rect 122840 68416 122892 68468
rect 276940 68416 276992 68468
rect 75920 68348 75972 68400
rect 256148 68348 256200 68400
rect 291108 68348 291160 68400
rect 476120 68348 476172 68400
rect 88984 68280 89036 68332
rect 307024 68280 307076 68332
rect 203524 67532 203576 67584
rect 289820 67532 289872 67584
rect 291108 67532 291160 67584
rect 22100 66852 22152 66904
rect 290556 66852 290608 66904
rect 20 66172 72 66224
rect 1308 66172 1360 66224
rect 251916 66172 251968 66224
rect 279424 66172 279476 66224
rect 480260 66172 480312 66224
rect 332600 66104 332652 66156
rect 385684 66104 385736 66156
rect 106280 65560 106332 65612
rect 260104 65628 260156 65680
rect 259552 65560 259604 65612
rect 334624 65560 334676 65612
rect 73160 65492 73212 65544
rect 279608 65492 279660 65544
rect 278780 65424 278832 65476
rect 279424 65424 279476 65476
rect 272524 64812 272576 64864
rect 481640 64812 481692 64864
rect 6920 64132 6972 64184
rect 281080 64132 281132 64184
rect 271880 63520 271932 63572
rect 272524 63520 272576 63572
rect 46940 62840 46992 62892
rect 258816 62840 258868 62892
rect 267740 62840 267792 62892
rect 483020 62840 483072 62892
rect 70400 62772 70452 62824
rect 285128 62772 285180 62824
rect 264980 62024 265032 62076
rect 265624 62024 265676 62076
rect 484400 62024 484452 62076
rect 74540 61412 74592 61464
rect 286508 61412 286560 61464
rect 53840 61344 53892 61396
rect 271328 61344 271380 61396
rect 261576 60664 261628 60716
rect 485780 60664 485832 60716
rect 515404 60664 515456 60716
rect 580172 60664 580224 60716
rect 260840 60256 260892 60308
rect 261576 60256 261628 60308
rect 111800 60120 111852 60172
rect 303068 60120 303120 60172
rect 64880 60052 64932 60104
rect 261484 60052 261536 60104
rect 4160 59984 4212 60036
rect 251824 59984 251876 60036
rect 3056 59304 3108 59356
rect 21364 59304 21416 59356
rect 85580 58760 85632 58812
rect 282460 58760 282512 58812
rect 259368 58692 259420 58744
rect 488540 58692 488592 58744
rect 69112 58624 69164 58676
rect 303160 58624 303212 58676
rect 254676 57944 254728 57996
rect 259368 57944 259420 57996
rect 71780 57264 71832 57316
rect 264336 57264 264388 57316
rect 246396 57196 246448 57248
rect 251272 57196 251324 57248
rect 489920 57196 489972 57248
rect 93952 55972 94004 56024
rect 268476 55972 268528 56024
rect 263600 55904 263652 55956
rect 491300 55904 491352 55956
rect 18604 55836 18656 55888
rect 307392 55836 307444 55888
rect 110420 54680 110472 54732
rect 250628 54680 250680 54732
rect 82820 54612 82872 54664
rect 275468 54612 275520 54664
rect 243544 54544 243596 54596
rect 475384 54544 475436 54596
rect 15200 54476 15252 54528
rect 307208 54476 307260 54528
rect 117320 53184 117372 53236
rect 294880 53184 294932 53236
rect 35808 53116 35860 53168
rect 132500 53116 132552 53168
rect 240784 53116 240836 53168
rect 492680 53116 492732 53168
rect 11060 53048 11112 53100
rect 267096 53048 267148 53100
rect 349804 52368 349856 52420
rect 495532 52368 495584 52420
rect 204996 51824 205048 51876
rect 241520 51824 241572 51876
rect 360936 51824 360988 51876
rect 120080 51756 120132 51808
rect 249064 51756 249116 51808
rect 114560 51688 114612 51740
rect 292028 51688 292080 51740
rect 349160 51076 349212 51128
rect 349804 51076 349856 51128
rect 244280 50532 244332 50584
rect 356704 50532 356756 50584
rect 113180 50464 113232 50516
rect 253296 50464 253348 50516
rect 85672 50396 85724 50448
rect 300308 50396 300360 50448
rect 19340 50328 19392 50380
rect 249248 50328 249300 50380
rect 192484 49648 192536 49700
rect 244280 49648 244332 49700
rect 358820 49648 358872 49700
rect 359280 49648 359332 49700
rect 494152 49648 494204 49700
rect 99380 49036 99432 49088
rect 304264 49036 304316 49088
rect 340880 49036 340932 49088
rect 359280 49036 359332 49088
rect 11152 48968 11204 49020
rect 284392 48968 284444 49020
rect 341524 48968 341576 49020
rect 285220 48900 285272 48952
rect 343640 48220 343692 48272
rect 344284 48220 344336 48272
rect 498200 48220 498252 48272
rect 118700 47608 118752 47660
rect 298928 47608 298980 47660
rect 23480 47540 23532 47592
rect 269856 47540 269908 47592
rect 269120 47472 269172 47524
rect 340236 47540 340288 47592
rect 544384 46860 544436 46912
rect 580172 46860 580224 46912
rect 284944 46248 284996 46300
rect 352564 46248 352616 46300
rect 26240 46180 26292 46232
rect 271236 46180 271288 46232
rect 334072 46180 334124 46232
rect 494428 46180 494480 46232
rect 3424 45500 3476 45552
rect 29644 45500 29696 45552
rect 280896 45500 280948 45552
rect 336004 45500 336056 45552
rect 95240 44956 95292 45008
rect 250444 44956 250496 45008
rect 121460 44888 121512 44940
rect 297456 44888 297508 44940
rect 27620 44820 27672 44872
rect 285036 44820 285088 44872
rect 316776 44820 316828 44872
rect 427820 44820 427872 44872
rect 280160 44140 280212 44192
rect 280896 44140 280948 44192
rect 92480 43460 92532 43512
rect 298836 43460 298888 43512
rect 320088 43460 320140 43512
rect 429200 43460 429252 43512
rect 57980 43392 58032 43444
rect 286600 43392 286652 43444
rect 298192 43392 298244 43444
rect 331864 43392 331916 43444
rect 342996 43392 343048 43444
rect 462320 43392 462372 43444
rect 322204 42712 322256 42764
rect 465080 42712 465132 42764
rect 276020 42644 276072 42696
rect 276664 42644 276716 42696
rect 342904 42644 342956 42696
rect 38660 42100 38712 42152
rect 264244 42100 264296 42152
rect 20720 42032 20772 42084
rect 301780 42032 301832 42084
rect 321560 41420 321612 41472
rect 322204 41420 322256 41472
rect 45560 40740 45612 40792
rect 273996 40740 274048 40792
rect 35900 40672 35952 40724
rect 300216 40672 300268 40724
rect 302240 40672 302292 40724
rect 433340 40672 433392 40724
rect 280804 39992 280856 40044
rect 296720 39992 296772 40044
rect 297364 39992 297416 40044
rect 59360 39380 59412 39432
rect 304356 39380 304408 39432
rect 2780 39312 2832 39364
rect 278320 39312 278372 39364
rect 299664 39312 299716 39364
rect 434720 39312 434772 39364
rect 196624 38020 196676 38072
rect 295340 38020 295392 38072
rect 91100 37952 91152 38004
rect 272616 37952 272668 38004
rect 436192 37952 436244 38004
rect 16580 37884 16632 37936
rect 296168 37884 296220 37936
rect 64696 37204 64748 37256
rect 307760 37204 307812 37256
rect 308496 37204 308548 37256
rect 195244 36592 195296 36644
rect 292580 36592 292632 36644
rect 436284 36592 436336 36644
rect 41420 36524 41472 36576
rect 293316 36524 293368 36576
rect 37188 35232 37240 35284
rect 135260 35232 135312 35284
rect 178684 35232 178736 35284
rect 256056 35232 256108 35284
rect 29000 35164 29052 35216
rect 287888 35164 287940 35216
rect 289728 35164 289780 35216
rect 437480 35164 437532 35216
rect 184296 34416 184348 34468
rect 288440 34416 288492 34468
rect 289728 34416 289780 34468
rect 60740 33736 60792 33788
rect 289084 33736 289136 33788
rect 3516 33056 3568 33108
rect 51724 33056 51776 33108
rect 180064 33056 180116 33108
rect 316132 33056 316184 33108
rect 316776 33056 316828 33108
rect 357440 33056 357492 33108
rect 425060 33056 425112 33108
rect 291844 32988 291896 33040
rect 356796 32988 356848 33040
rect 80060 32444 80112 32496
rect 250536 32444 250588 32496
rect 62120 32376 62172 32428
rect 283748 32376 283800 32428
rect 327080 32376 327132 32428
rect 357440 32376 357492 32428
rect 291200 31764 291252 31816
rect 291844 31764 291896 31816
rect 44180 31084 44232 31136
rect 274088 31084 274140 31136
rect 282184 31084 282236 31136
rect 438860 31084 438912 31136
rect 24860 31016 24912 31068
rect 302976 31016 303028 31068
rect 277400 30268 277452 30320
rect 278044 30268 278096 30320
rect 441620 30268 441672 30320
rect 52460 29656 52512 29708
rect 265716 29656 265768 29708
rect 64788 29588 64840 29640
rect 309968 29588 310020 29640
rect 81440 28228 81492 28280
rect 275376 28228 275428 28280
rect 280804 28228 280856 28280
rect 443000 28228 443052 28280
rect 51080 26868 51132 26920
rect 255964 26868 256016 26920
rect 270592 26868 270644 26920
rect 444380 26868 444432 26920
rect 196716 25644 196768 25696
rect 274640 25644 274692 25696
rect 445852 25644 445904 25696
rect 35992 25576 36044 25628
rect 276756 25576 276808 25628
rect 40040 25508 40092 25560
rect 289268 25508 289320 25560
rect 118792 24216 118844 24268
rect 286416 24216 286468 24268
rect 263692 24148 263744 24200
rect 445944 24148 445996 24200
rect 48320 24080 48372 24132
rect 267004 24080 267056 24132
rect 43444 23400 43496 23452
rect 44088 23400 44140 23452
rect 249800 23400 249852 23452
rect 186964 22788 187016 22840
rect 259460 22788 259512 22840
rect 447140 22788 447192 22840
rect 52552 22720 52604 22772
rect 290464 22720 290516 22772
rect 253388 22040 253440 22092
rect 449900 22040 449952 22092
rect 252560 21564 252612 21616
rect 253388 21564 253440 21616
rect 30380 21360 30432 21412
rect 280988 21360 281040 21412
rect 3424 20612 3476 20664
rect 57244 20612 57296 20664
rect 64604 20612 64656 20664
rect 246304 20612 246356 20664
rect 249800 20612 249852 20664
rect 250812 20612 250864 20664
rect 509148 20612 509200 20664
rect 579988 20612 580040 20664
rect 248420 20544 248472 20596
rect 249156 20544 249208 20596
rect 250812 20000 250864 20052
rect 451280 20000 451332 20052
rect 56600 19932 56652 19984
rect 278136 19932 278188 19984
rect 100760 18708 100812 18760
rect 257436 18708 257488 18760
rect 246304 18640 246356 18692
rect 452660 18640 452712 18692
rect 27712 18572 27764 18624
rect 301688 18572 301740 18624
rect 103520 17280 103572 17332
rect 302884 17280 302936 17332
rect 37280 17212 37332 17264
rect 268384 17212 268436 17264
rect 271236 17212 271288 17264
rect 454132 17212 454184 17264
rect 301504 16532 301556 16584
rect 363604 16532 363656 16584
rect 108120 15920 108172 15972
rect 279516 15920 279568 15972
rect 286416 15920 286468 15972
rect 454040 15920 454092 15972
rect 19432 15852 19484 15904
rect 287796 15852 287848 15904
rect 84200 14560 84252 14612
rect 258724 14560 258776 14612
rect 66720 14492 66772 14544
rect 305736 14492 305788 14544
rect 164424 14424 164476 14476
rect 414664 14424 414716 14476
rect 314660 13744 314712 13796
rect 315304 13744 315356 13796
rect 467840 13744 467892 13796
rect 255872 13676 255924 13728
rect 256056 13676 256108 13728
rect 353944 13676 353996 13728
rect 191104 13200 191156 13252
rect 257436 13200 257488 13252
rect 97448 13132 97500 13184
rect 253204 13132 253256 13184
rect 56048 13064 56100 13116
rect 305828 13064 305880 13116
rect 283104 12384 283156 12436
rect 283564 12384 283616 12436
rect 478880 12384 478932 12436
rect 77392 11772 77444 11824
rect 257344 11772 257396 11824
rect 98184 11704 98236 11756
rect 298744 11704 298796 11756
rect 360844 10956 360896 11008
rect 421564 10956 421616 11008
rect 258448 10888 258500 10940
rect 259368 10888 259420 10940
rect 124680 10276 124732 10328
rect 254584 10276 254636 10328
rect 259368 10276 259420 10328
rect 486424 10276 486476 10328
rect 284944 9596 284996 9648
rect 287796 9596 287848 9648
rect 305644 9596 305696 9648
rect 374644 9596 374696 9648
rect 3424 8984 3476 9036
rect 35164 8984 35216 9036
rect 62028 8984 62080 9036
rect 282368 8984 282420 9036
rect 34796 8916 34848 8968
rect 296076 8916 296128 8968
rect 339868 8916 339920 8968
rect 423680 8916 423732 8968
rect 188344 7692 188396 7744
rect 109316 7624 109368 7676
rect 232504 7624 232556 7676
rect 1676 7556 1728 7608
rect 43444 7556 43496 7608
rect 45468 7556 45520 7608
rect 271144 7556 271196 7608
rect 306748 7556 306800 7608
rect 431960 7556 432012 7608
rect 282276 6808 282328 6860
rect 439504 6808 439556 6860
rect 543004 6808 543056 6860
rect 580172 6808 580224 6860
rect 308588 6740 308640 6792
rect 309876 6740 309928 6792
rect 309968 6740 310020 6792
rect 430580 6740 430632 6792
rect 79692 6196 79744 6248
rect 301596 6196 301648 6248
rect 14740 6128 14792 6180
rect 283656 6128 283708 6180
rect 257068 5448 257120 5500
rect 257436 5448 257488 5500
rect 448520 5448 448572 5500
rect 43076 4836 43128 4888
rect 291936 4836 291988 4888
rect 8760 4768 8812 4820
rect 269764 4768 269816 4820
rect 293960 4768 294012 4820
rect 294880 4768 294932 4820
rect 359464 4768 359516 4820
rect 198004 4088 198056 4140
rect 246396 4088 246448 4140
rect 332692 4088 332744 4140
rect 333244 4088 333296 4140
rect 342996 4088 343048 4140
rect 351184 4088 351236 4140
rect 351644 4088 351696 4140
rect 374000 4088 374052 4140
rect 216036 4020 216088 4072
rect 240508 4020 240560 4072
rect 240784 4020 240836 4072
rect 294604 4020 294656 4072
rect 323308 4020 323360 4072
rect 331588 4020 331640 4072
rect 339868 4020 339920 4072
rect 346952 4020 347004 4072
rect 352656 4020 352708 4072
rect 274824 3952 274876 4004
rect 275284 3952 275336 4004
rect 280804 3952 280856 4004
rect 309784 3952 309836 4004
rect 320916 3952 320968 4004
rect 273904 3884 273956 3936
rect 293960 3884 294012 3936
rect 308404 3884 308456 3936
rect 319720 3884 319772 3936
rect 287704 3816 287756 3868
rect 316224 3816 316276 3868
rect 316684 3816 316736 3868
rect 125876 3612 125928 3664
rect 164884 3612 164936 3664
rect 251180 3612 251232 3664
rect 252376 3612 252428 3664
rect 78588 3544 78640 3596
rect 88984 3544 89036 3596
rect 93860 3544 93912 3596
rect 94780 3544 94832 3596
rect 103336 3544 103388 3596
rect 170404 3544 170456 3596
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 6460 3476 6512 3528
rect 18604 3476 18656 3528
rect 19340 3476 19392 3528
rect 20260 3476 20312 3528
rect 27620 3476 27672 3528
rect 28540 3476 28592 3528
rect 35900 3476 35952 3528
rect 36820 3476 36872 3528
rect 69020 3476 69072 3528
rect 69940 3476 69992 3528
rect 89168 3476 89220 3528
rect 178776 3476 178828 3528
rect 217324 3476 217376 3528
rect 242992 3544 243044 3596
rect 242900 3476 242952 3528
rect 244096 3476 244148 3528
rect 247592 3544 247644 3596
rect 263600 3612 263652 3664
rect 259460 3544 259512 3596
rect 260656 3544 260708 3596
rect 271236 3544 271288 3596
rect 276020 3476 276072 3528
rect 276848 3476 276900 3528
rect 307760 3476 307812 3528
rect 309048 3476 309100 3528
rect 316132 3476 316184 3528
rect 317328 3476 317380 3528
rect 324964 3476 325016 3528
rect 325608 3476 325660 3528
rect 329196 3476 329248 3528
rect 331220 3476 331272 3528
rect 332600 3476 332652 3528
rect 333888 3476 333940 3528
rect 340880 3476 340932 3528
rect 342168 3476 342220 3528
rect 350448 3476 350500 3528
rect 360844 3476 360896 3528
rect 18236 3408 18288 3460
rect 202236 3408 202288 3460
rect 215944 3408 215996 3460
rect 239312 3408 239364 3460
rect 286416 3408 286468 3460
rect 313832 3408 313884 3460
rect 318892 3408 318944 3460
rect 342076 3408 342128 3460
rect 500960 3408 501012 3460
rect 135260 3340 135312 3392
rect 136456 3340 136508 3392
rect 267740 3340 267792 3392
rect 274640 3340 274692 3392
rect 282184 3272 282236 3324
rect 285404 3272 285456 3324
rect 235816 3000 235868 3052
rect 238024 3000 238076 3052
rect 41328 2184 41380 2236
rect 129372 2184 129424 2236
rect 111616 2116 111668 2168
rect 294788 2116 294840 2168
rect 64328 2048 64380 2100
rect 294696 2048 294748 2100
<< metal2 >>
rect 6932 703582 7972 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 595474 3464 684247
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3516 632120 3568 632126
rect 3514 632088 3516 632097
rect 3568 632088 3570 632097
rect 3514 632023 3570 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618322 3556 619103
rect 3516 618316 3568 618322
rect 3516 618258 3568 618264
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3424 595468 3476 595474
rect 3424 595410 3476 595416
rect 3528 594114 3556 606047
rect 6932 598262 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 698970 24348 703520
rect 24308 698964 24360 698970
rect 24308 698906 24360 698912
rect 15844 670744 15896 670750
rect 15844 670686 15896 670692
rect 11704 656940 11756 656946
rect 11704 656882 11756 656888
rect 6920 598256 6972 598262
rect 6920 598198 6972 598204
rect 3516 594108 3568 594114
rect 3516 594050 3568 594056
rect 11716 588606 11744 656882
rect 11704 588600 11756 588606
rect 11704 588542 11756 588548
rect 14464 582412 14516 582418
rect 14464 582354 14516 582360
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3436 539578 3464 579935
rect 14476 554742 14504 582354
rect 3516 554736 3568 554742
rect 3516 554678 3568 554684
rect 14464 554736 14516 554742
rect 14464 554678 14516 554684
rect 3528 553897 3556 554678
rect 3514 553888 3570 553897
rect 3514 553823 3570 553832
rect 3424 539572 3476 539578
rect 3424 539514 3476 539520
rect 15856 537538 15884 670686
rect 40052 590714 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 77944 703316 77996 703322
rect 77944 703258 77996 703264
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 76564 703044 76616 703050
rect 76564 702986 76616 702992
rect 68928 702500 68980 702506
rect 68928 702442 68980 702448
rect 62028 700324 62080 700330
rect 62028 700266 62080 700272
rect 57888 697604 57940 697610
rect 57888 697546 57940 697552
rect 46848 598256 46900 598262
rect 46848 598198 46900 598204
rect 46860 597582 46888 598198
rect 46848 597576 46900 597582
rect 46848 597518 46900 597524
rect 42800 595468 42852 595474
rect 42800 595410 42852 595416
rect 42812 594862 42840 595410
rect 42800 594856 42852 594862
rect 42800 594798 42852 594804
rect 44088 594856 44140 594862
rect 44088 594798 44140 594804
rect 40040 590708 40092 590714
rect 40040 590650 40092 590656
rect 39856 584044 39908 584050
rect 39856 583986 39908 583992
rect 35808 581052 35860 581058
rect 35808 580994 35860 581000
rect 34428 572824 34480 572830
rect 34428 572766 34480 572772
rect 25504 565888 25556 565894
rect 25504 565830 25556 565836
rect 25516 544406 25544 565830
rect 30288 557592 30340 557598
rect 30288 557534 30340 557540
rect 25504 544400 25556 544406
rect 25504 544342 25556 544348
rect 15844 537532 15896 537538
rect 15844 537474 15896 537480
rect 3148 528556 3200 528562
rect 3148 528498 3200 528504
rect 3160 527921 3188 528498
rect 3146 527912 3202 527921
rect 3146 527847 3202 527856
rect 2778 514856 2834 514865
rect 2778 514791 2780 514800
rect 2832 514791 2834 514800
rect 4804 514820 4856 514826
rect 2780 514762 2832 514768
rect 4804 514762 4856 514768
rect 3422 501800 3478 501809
rect 3422 501735 3478 501744
rect 3436 495446 3464 501735
rect 4816 498166 4844 514762
rect 4804 498160 4856 498166
rect 4804 498102 4856 498108
rect 3424 495440 3476 495446
rect 3424 495382 3476 495388
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 25504 474768 25556 474774
rect 25504 474710 25556 474716
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 4804 462596 4856 462602
rect 2780 462538 2832 462544
rect 4804 462538 4856 462544
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 4816 438870 4844 462538
rect 25516 438938 25544 474710
rect 30300 458182 30328 557534
rect 33048 545148 33100 545154
rect 33048 545090 33100 545096
rect 30288 458176 30340 458182
rect 30288 458118 30340 458124
rect 33060 446418 33088 545090
rect 34336 488572 34388 488578
rect 34336 488514 34388 488520
rect 33784 458312 33836 458318
rect 33784 458254 33836 458260
rect 33048 446412 33100 446418
rect 33048 446354 33100 446360
rect 25504 438932 25556 438938
rect 25504 438874 25556 438880
rect 4804 438864 4856 438870
rect 4804 438806 4856 438812
rect 3424 429888 3476 429894
rect 3424 429830 3476 429836
rect 3436 410553 3464 429830
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3148 398132 3200 398138
rect 3148 398074 3200 398080
rect 3160 397497 3188 398074
rect 3146 397488 3202 397497
rect 3146 397423 3202 397432
rect 4804 388476 4856 388482
rect 4804 388418 4856 388424
rect 3240 372564 3292 372570
rect 3240 372506 3292 372512
rect 3252 371385 3280 372506
rect 3238 371376 3294 371385
rect 3238 371311 3294 371320
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 4816 346322 4844 388418
rect 7564 351960 7616 351966
rect 7564 351902 7616 351908
rect 2780 346316 2832 346322
rect 2780 346258 2832 346264
rect 4804 346316 4856 346322
rect 4804 346258 4856 346264
rect 2792 345409 2820 346258
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 310486 3464 319223
rect 3424 310480 3476 310486
rect 3424 310422 3476 310428
rect 7576 306270 7604 351902
rect 33060 347721 33088 446354
rect 33796 360097 33824 458254
rect 34348 390726 34376 488514
rect 34440 474706 34468 572766
rect 35716 554804 35768 554810
rect 35716 554746 35768 554752
rect 34428 474700 34480 474706
rect 34428 474642 34480 474648
rect 35164 458924 35216 458930
rect 35164 458866 35216 458872
rect 34336 390720 34388 390726
rect 34336 390662 34388 390668
rect 34428 383716 34480 383722
rect 34428 383658 34480 383664
rect 34336 365628 34388 365634
rect 34336 365570 34388 365576
rect 34348 363662 34376 365570
rect 34336 363656 34388 363662
rect 34336 363598 34388 363604
rect 33782 360088 33838 360097
rect 33782 360023 33838 360032
rect 33046 347712 33102 347721
rect 33046 347647 33102 347656
rect 14464 324352 14516 324358
rect 14464 324294 14516 324300
rect 3424 306264 3476 306270
rect 3422 306232 3424 306241
rect 7564 306264 7616 306270
rect 3476 306232 3478 306241
rect 7564 306206 7616 306212
rect 3422 306167 3478 306176
rect 14476 293962 14504 324294
rect 3056 293956 3108 293962
rect 3056 293898 3108 293904
rect 14464 293956 14516 293962
rect 14464 293898 14516 293904
rect 3068 293185 3096 293898
rect 21364 293276 21416 293282
rect 21364 293218 21416 293224
rect 3054 293176 3110 293185
rect 3054 293111 3110 293120
rect 4068 291848 4120 291854
rect 4068 291790 4120 291796
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3424 255264 3476 255270
rect 3424 255206 3476 255212
rect 3436 254153 3464 255206
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3146 241088 3202 241097
rect 3146 241023 3202 241032
rect 3160 240106 3188 241023
rect 3148 240100 3200 240106
rect 3148 240042 3200 240048
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 214606 3464 214911
rect 3424 214600 3476 214606
rect 3424 214542 3476 214548
rect 3240 205012 3292 205018
rect 3240 204954 3292 204960
rect 3252 201929 3280 204954
rect 3238 201920 3294 201929
rect 3238 201855 3294 201864
rect 4080 193254 4108 291790
rect 15844 257372 15896 257378
rect 15844 257314 15896 257320
rect 4804 221468 4856 221474
rect 4804 221410 4856 221416
rect 3424 193248 3476 193254
rect 3424 193190 3476 193196
rect 4068 193248 4120 193254
rect 4068 193190 4120 193196
rect 1306 181384 1362 181393
rect 1306 181319 1362 181328
rect 1320 66230 1348 181319
rect 3436 162897 3464 193190
rect 3516 188896 3568 188902
rect 3514 188864 3516 188873
rect 3568 188864 3570 188873
rect 3514 188799 3570 188808
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3700 111104 3752 111110
rect 3700 111046 3752 111052
rect 4068 111104 4120 111110
rect 4068 111046 4120 111052
rect 3712 110673 3740 111046
rect 3698 110664 3754 110673
rect 3698 110599 3754 110608
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 4080 93809 4108 111046
rect 4816 97782 4844 221410
rect 7564 202156 7616 202162
rect 7564 202098 7616 202104
rect 7576 188902 7604 202098
rect 7564 188896 7616 188902
rect 7564 188838 7616 188844
rect 7564 177336 7616 177342
rect 7564 177278 7616 177284
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 4066 93800 4122 93809
rect 4066 93735 4122 93744
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 7576 71670 7604 177278
rect 14464 175976 14516 175982
rect 14464 175918 14516 175924
rect 14476 111110 14504 175918
rect 15856 137970 15884 257314
rect 17224 253224 17276 253230
rect 17224 253166 17276 253172
rect 15844 137964 15896 137970
rect 15844 137906 15896 137912
rect 14464 111104 14516 111110
rect 14464 111046 14516 111052
rect 17236 85542 17264 253166
rect 17224 85536 17276 85542
rect 17224 85478 17276 85484
rect 12438 76528 12494 76537
rect 12438 76463 12494 76472
rect 3424 71664 3476 71670
rect 3422 71632 3424 71641
rect 7564 71664 7616 71670
rect 3476 71632 3478 71641
rect 7564 71606 7616 71612
rect 3422 71567 3478 71576
rect 20 66224 72 66230
rect 20 66166 72 66172
rect 1308 66224 1360 66230
rect 1308 66166 1360 66172
rect 32 16574 60 66166
rect 6920 64184 6972 64190
rect 6920 64126 6972 64132
rect 4160 60036 4212 60042
rect 4160 59978 4212 59984
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2780 39364 2832 39370
rect 2780 39306 2832 39312
rect 32 16546 152 16574
rect 124 354 152 16546
rect 1676 7608 1728 7614
rect 1676 7550 1728 7556
rect 1688 480 1716 7550
rect 2792 3534 2820 39306
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 2870 28248 2926 28257
rect 2870 28183 2926 28192
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 480 2912 28183
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 59978
rect 6932 16574 6960 64126
rect 11060 53100 11112 53106
rect 11060 53042 11112 53048
rect 9678 26888 9734 26897
rect 9678 26823 9734 26832
rect 4172 16546 5304 16574
rect 6932 16546 7696 16574
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3436 6497 3464 8978
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 5276 480 5304 16546
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6472 480 6500 3470
rect 7668 480 7696 16546
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8772 480 8800 4762
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 26823
rect 11072 6914 11100 53042
rect 11152 49020 11204 49026
rect 11152 48962 11204 48968
rect 11164 16574 11192 48962
rect 12452 16574 12480 76463
rect 21376 59362 21404 293218
rect 22744 290488 22796 290494
rect 22744 290430 22796 290436
rect 22756 150414 22784 290430
rect 25504 266416 25556 266422
rect 25504 266358 25556 266364
rect 25516 238678 25544 266358
rect 33140 255264 33192 255270
rect 33140 255206 33192 255212
rect 33152 254590 33180 255206
rect 33140 254584 33192 254590
rect 33140 254526 33192 254532
rect 33600 240100 33652 240106
rect 33600 240042 33652 240048
rect 33612 239426 33640 240042
rect 34348 239426 34376 363598
rect 34440 254590 34468 383658
rect 35176 365634 35204 458866
rect 35728 456074 35756 554746
rect 35820 489870 35848 580994
rect 37188 575544 37240 575550
rect 37188 575486 37240 575492
rect 37096 558204 37148 558210
rect 37096 558146 37148 558152
rect 35808 489864 35860 489870
rect 35808 489806 35860 489812
rect 35820 488578 35848 489806
rect 35808 488572 35860 488578
rect 35808 488514 35860 488520
rect 37004 483064 37056 483070
rect 37004 483006 37056 483012
rect 35808 476128 35860 476134
rect 35808 476070 35860 476076
rect 35716 456068 35768 456074
rect 35716 456010 35768 456016
rect 35728 455394 35756 456010
rect 35716 455388 35768 455394
rect 35716 455330 35768 455336
rect 35164 365628 35216 365634
rect 35164 365570 35216 365576
rect 35716 362228 35768 362234
rect 35716 362170 35768 362176
rect 35164 279472 35216 279478
rect 35164 279414 35216 279420
rect 34428 254584 34480 254590
rect 34428 254526 34480 254532
rect 33600 239420 33652 239426
rect 33600 239362 33652 239368
rect 34336 239420 34388 239426
rect 34336 239362 34388 239368
rect 25504 238672 25556 238678
rect 25504 238614 25556 238620
rect 29644 180192 29696 180198
rect 29644 180134 29696 180140
rect 22744 150408 22796 150414
rect 22744 150350 22796 150356
rect 22100 66904 22152 66910
rect 22100 66846 22152 66852
rect 21364 59356 21416 59362
rect 21364 59298 21416 59304
rect 18604 55888 18656 55894
rect 18604 55830 18656 55836
rect 15200 54528 15252 54534
rect 15200 54470 15252 54476
rect 15212 16574 15240 54470
rect 16580 37936 16632 37942
rect 16580 37878 16632 37884
rect 16592 16574 16620 37878
rect 11164 16546 11928 16574
rect 12452 16546 13584 16574
rect 15212 16546 15976 16574
rect 16592 16546 17080 16574
rect 11072 6886 11192 6914
rect 11164 480 11192 6886
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13556 480 13584 16546
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 14752 480 14780 6122
rect 15948 480 15976 16546
rect 17052 480 17080 16546
rect 18616 3534 18644 55830
rect 19340 50380 19392 50386
rect 19340 50322 19392 50328
rect 19352 3534 19380 50322
rect 20720 42084 20772 42090
rect 20720 42026 20772 42032
rect 20732 16574 20760 42026
rect 22112 16574 22140 66846
rect 23480 47592 23532 47598
rect 23480 47534 23532 47540
rect 23492 16574 23520 47534
rect 26240 46232 26292 46238
rect 26240 46174 26292 46180
rect 24860 31068 24912 31074
rect 24860 31010 24912 31016
rect 24872 16574 24900 31010
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 23492 16546 24256 16574
rect 24872 16546 25360 16574
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18248 480 18276 3402
rect 19444 480 19472 15846
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20272 354 20300 3470
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20272 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24228 480 24256 16546
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 46174
rect 29656 45558 29684 180134
rect 33140 72480 33192 72486
rect 33140 72422 33192 72428
rect 31758 46200 31814 46209
rect 31758 46135 31814 46144
rect 29644 45552 29696 45558
rect 29644 45494 29696 45500
rect 27620 44872 27672 44878
rect 27620 44814 27672 44820
rect 27632 3534 27660 44814
rect 29000 35216 29052 35222
rect 29000 35158 29052 35164
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27724 480 27752 18566
rect 29012 16574 29040 35158
rect 30380 21412 30432 21418
rect 30380 21354 30432 21360
rect 30392 16574 30420 21354
rect 31772 16574 31800 46135
rect 33152 16574 33180 72422
rect 29012 16546 30144 16574
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 33152 16546 33640 16574
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28552 354 28580 3470
rect 30116 480 30144 16546
rect 28878 354 28990 480
rect 28552 326 28990 354
rect 28878 -960 28990 326
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33612 480 33640 16546
rect 35176 9042 35204 279414
rect 35728 253230 35756 362170
rect 35716 253224 35768 253230
rect 35716 253166 35768 253172
rect 35820 53174 35848 476070
rect 36636 455388 36688 455394
rect 36636 455330 36688 455336
rect 36544 390720 36596 390726
rect 36544 390662 36596 390668
rect 36556 258058 36584 390662
rect 36648 358086 36676 455330
rect 37016 402974 37044 483006
rect 37108 458862 37136 558146
rect 37096 458856 37148 458862
rect 37096 458798 37148 458804
rect 37016 402946 37136 402974
rect 37108 389162 37136 402946
rect 37096 389156 37148 389162
rect 37096 389098 37148 389104
rect 37108 388482 37136 389098
rect 37096 388476 37148 388482
rect 37096 388418 37148 388424
rect 36636 358080 36688 358086
rect 36636 358022 36688 358028
rect 36636 264240 36688 264246
rect 36636 264182 36688 264188
rect 36544 258052 36596 258058
rect 36544 257994 36596 258000
rect 36556 257378 36584 257994
rect 36544 257372 36596 257378
rect 36544 257314 36596 257320
rect 36648 214606 36676 264182
rect 36636 214600 36688 214606
rect 36636 214542 36688 214548
rect 35808 53168 35860 53174
rect 35808 53110 35860 53116
rect 35900 40724 35952 40730
rect 35900 40666 35952 40672
rect 35164 9036 35216 9042
rect 35164 8978 35216 8984
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34808 480 34836 8910
rect 35912 3534 35940 40666
rect 37200 35290 37228 575486
rect 38476 536104 38528 536110
rect 38476 536046 38528 536052
rect 38488 437442 38516 536046
rect 39672 532024 39724 532030
rect 39672 531966 39724 531972
rect 38566 525872 38622 525881
rect 38566 525807 38622 525816
rect 38580 442270 38608 525807
rect 38568 442264 38620 442270
rect 38568 442206 38620 442212
rect 38476 437436 38528 437442
rect 38476 437378 38528 437384
rect 38476 433288 38528 433294
rect 38476 433230 38528 433236
rect 38488 338094 38516 433230
rect 38580 341562 38608 442206
rect 39684 437306 39712 531966
rect 39868 492726 39896 583986
rect 41236 583908 41288 583914
rect 41236 583850 41288 583856
rect 41144 549296 41196 549302
rect 41144 549238 41196 549244
rect 39948 534744 40000 534750
rect 39948 534686 40000 534692
rect 39856 492720 39908 492726
rect 39856 492662 39908 492668
rect 39764 492040 39816 492046
rect 39764 491982 39816 491988
rect 39672 437300 39724 437306
rect 39672 437242 39724 437248
rect 39580 394868 39632 394874
rect 39580 394810 39632 394816
rect 38568 341556 38620 341562
rect 38568 341498 38620 341504
rect 38476 338088 38528 338094
rect 38476 338030 38528 338036
rect 39592 267714 39620 394810
rect 39684 336598 39712 437242
rect 39776 391338 39804 491982
rect 39868 393990 39896 492662
rect 39960 434722 39988 534686
rect 41052 529304 41104 529310
rect 41052 529246 41104 529252
rect 40684 435396 40736 435402
rect 40684 435338 40736 435344
rect 40696 434722 40724 435338
rect 39948 434716 40000 434722
rect 39948 434658 40000 434664
rect 40684 434716 40736 434722
rect 40684 434658 40736 434664
rect 39856 393984 39908 393990
rect 39856 393926 39908 393932
rect 39764 391332 39816 391338
rect 39764 391274 39816 391280
rect 39764 386504 39816 386510
rect 39764 386446 39816 386452
rect 39672 336592 39724 336598
rect 39672 336534 39724 336540
rect 39776 274650 39804 386446
rect 40696 339386 40724 434658
rect 41064 433294 41092 529246
rect 41156 449886 41184 549238
rect 41248 486470 41276 583850
rect 42708 558952 42760 558958
rect 42708 558894 42760 558900
rect 41328 538280 41380 538286
rect 41328 538222 41380 538228
rect 41236 486464 41288 486470
rect 41236 486406 41288 486412
rect 41144 449880 41196 449886
rect 41144 449822 41196 449828
rect 41052 433288 41104 433294
rect 41052 433230 41104 433236
rect 41144 388476 41196 388482
rect 41144 388418 41196 388424
rect 40684 339380 40736 339386
rect 40684 339322 40736 339328
rect 39948 288448 40000 288454
rect 39948 288390 40000 288396
rect 39764 274644 39816 274650
rect 39764 274586 39816 274592
rect 39580 267708 39632 267714
rect 39580 267650 39632 267656
rect 39960 77217 39988 288390
rect 41156 249082 41184 388418
rect 41248 385830 41276 486406
rect 41340 437238 41368 538222
rect 42524 529236 42576 529242
rect 42524 529178 42576 529184
rect 42432 456748 42484 456754
rect 42432 456690 42484 456696
rect 41328 437232 41380 437238
rect 41328 437174 41380 437180
rect 41236 385824 41288 385830
rect 41236 385766 41288 385772
rect 41328 382288 41380 382294
rect 41328 382230 41380 382236
rect 41144 249076 41196 249082
rect 41144 249018 41196 249024
rect 39946 77208 40002 77217
rect 39946 77143 40002 77152
rect 38660 42152 38712 42158
rect 38660 42094 38712 42100
rect 37188 35284 37240 35290
rect 37188 35226 37240 35232
rect 35992 25628 36044 25634
rect 35992 25570 36044 25576
rect 35900 3528 35952 3534
rect 35900 3470 35952 3476
rect 36004 480 36032 25570
rect 37280 17264 37332 17270
rect 37280 17206 37332 17212
rect 37292 16574 37320 17206
rect 38672 16574 38700 42094
rect 40040 25560 40092 25566
rect 40040 25502 40092 25508
rect 40052 16574 40080 25502
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 40052 16546 40264 16574
rect 36820 3528 36872 3534
rect 36820 3470 36872 3476
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 36832 354 36860 3470
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36832 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41340 2242 41368 382230
rect 42444 362982 42472 456690
rect 42536 435470 42564 529178
rect 42616 490612 42668 490618
rect 42616 490554 42668 490560
rect 42524 435464 42576 435470
rect 42524 435406 42576 435412
rect 42628 395350 42656 490554
rect 42720 460222 42748 558894
rect 43904 556232 43956 556238
rect 43904 556174 43956 556180
rect 43812 469260 43864 469266
rect 43812 469202 43864 469208
rect 42708 460216 42760 460222
rect 42708 460158 42760 460164
rect 42720 458930 42748 460158
rect 42708 458924 42760 458930
rect 42708 458866 42760 458872
rect 43720 458176 43772 458182
rect 43720 458118 43772 458124
rect 42706 433256 42762 433265
rect 42706 433191 42762 433200
rect 42616 395344 42668 395350
rect 42616 395286 42668 395292
rect 42616 375420 42668 375426
rect 42616 375362 42668 375368
rect 42432 362976 42484 362982
rect 42432 362918 42484 362924
rect 42444 362234 42472 362918
rect 42432 362228 42484 362234
rect 42432 362170 42484 362176
rect 42628 302161 42656 375362
rect 42720 335238 42748 433191
rect 43732 359514 43760 458118
rect 43824 375358 43852 469202
rect 43916 457502 43944 556174
rect 43996 493332 44048 493338
rect 43996 493274 44048 493280
rect 43904 457496 43956 457502
rect 43904 457438 43956 457444
rect 44008 392630 44036 493274
rect 44100 484362 44128 594798
rect 46756 550656 46808 550662
rect 46756 550598 46808 550604
rect 45468 542428 45520 542434
rect 45468 542370 45520 542376
rect 45284 534812 45336 534818
rect 45284 534754 45336 534760
rect 44088 484356 44140 484362
rect 44088 484298 44140 484304
rect 44088 457496 44140 457502
rect 44088 457438 44140 457444
rect 44100 456754 44128 457438
rect 44088 456748 44140 456754
rect 44088 456690 44140 456696
rect 45296 440910 45324 534754
rect 45376 532092 45428 532098
rect 45376 532034 45428 532040
rect 45284 440904 45336 440910
rect 45284 440846 45336 440852
rect 44272 438252 44324 438258
rect 44272 438194 44324 438200
rect 44284 437442 44312 438194
rect 44272 437436 44324 437442
rect 44272 437378 44324 437384
rect 44824 437436 44876 437442
rect 44824 437378 44876 437384
rect 44088 435464 44140 435470
rect 44088 435406 44140 435412
rect 43996 392624 44048 392630
rect 43996 392566 44048 392572
rect 43996 385688 44048 385694
rect 43996 385630 44048 385636
rect 43812 375352 43864 375358
rect 43812 375294 43864 375300
rect 43720 359508 43772 359514
rect 43720 359450 43772 359456
rect 43444 357468 43496 357474
rect 43444 357410 43496 357416
rect 42800 352572 42852 352578
rect 42800 352514 42852 352520
rect 42812 351966 42840 352514
rect 42800 351960 42852 351966
rect 42800 351902 42852 351908
rect 43456 346390 43484 357410
rect 43904 352572 43956 352578
rect 43904 352514 43956 352520
rect 43444 346384 43496 346390
rect 43444 346326 43496 346332
rect 42708 335232 42760 335238
rect 42708 335174 42760 335180
rect 42614 302152 42670 302161
rect 42614 302087 42670 302096
rect 43916 301510 43944 352514
rect 43904 301504 43956 301510
rect 43904 301446 43956 301452
rect 42708 277432 42760 277438
rect 42708 277374 42760 277380
rect 42720 213314 42748 277374
rect 43904 270564 43956 270570
rect 43904 270506 43956 270512
rect 42708 213308 42760 213314
rect 42708 213250 42760 213256
rect 43916 192710 43944 270506
rect 44008 262954 44036 385630
rect 44100 335170 44128 435406
rect 44836 337958 44864 437378
rect 45388 436014 45416 532034
rect 45480 443698 45508 542370
rect 46664 537668 46716 537674
rect 46664 537610 46716 537616
rect 46572 492788 46624 492794
rect 46572 492730 46624 492736
rect 45468 443692 45520 443698
rect 45468 443634 45520 443640
rect 45376 436008 45428 436014
rect 45376 435950 45428 435956
rect 45374 357504 45430 357513
rect 45374 357439 45430 357448
rect 44824 337952 44876 337958
rect 44824 337894 44876 337900
rect 44088 335164 44140 335170
rect 44088 335106 44140 335112
rect 44088 294024 44140 294030
rect 44088 293966 44140 293972
rect 43996 262948 44048 262954
rect 43996 262890 44048 262896
rect 43904 192704 43956 192710
rect 43904 192646 43956 192652
rect 41420 36576 41472 36582
rect 41420 36518 41472 36524
rect 41432 16574 41460 36518
rect 44100 23458 44128 293966
rect 45388 280158 45416 357439
rect 45480 344350 45508 443634
rect 46584 395418 46612 492730
rect 46676 438802 46704 537610
rect 46768 451246 46796 550598
rect 46860 491298 46888 597518
rect 48228 590708 48280 590714
rect 48228 590650 48280 590656
rect 48044 581120 48096 581126
rect 48044 581062 48096 581068
rect 48056 492046 48084 581062
rect 48136 556300 48188 556306
rect 48136 556242 48188 556248
rect 48044 492040 48096 492046
rect 48044 491982 48096 491988
rect 46848 491292 46900 491298
rect 46848 491234 46900 491240
rect 47584 484492 47636 484498
rect 47584 484434 47636 484440
rect 46848 454028 46900 454034
rect 46848 453970 46900 453976
rect 46756 451240 46808 451246
rect 46756 451182 46808 451188
rect 46664 438796 46716 438802
rect 46664 438738 46716 438744
rect 46756 396772 46808 396778
rect 46756 396714 46808 396720
rect 46572 395412 46624 395418
rect 46572 395354 46624 395360
rect 46664 385756 46716 385762
rect 46664 385698 46716 385704
rect 45468 344344 45520 344350
rect 45468 344286 45520 344292
rect 46676 333946 46704 385698
rect 46768 336530 46796 396714
rect 46860 355978 46888 453970
rect 47596 391270 47624 484434
rect 48044 481704 48096 481710
rect 48044 481646 48096 481652
rect 47952 394052 48004 394058
rect 47952 393994 48004 394000
rect 47584 391264 47636 391270
rect 47584 391206 47636 391212
rect 46848 355972 46900 355978
rect 46848 355914 46900 355920
rect 46848 350600 46900 350606
rect 46848 350542 46900 350548
rect 46756 336524 46808 336530
rect 46756 336466 46808 336472
rect 46664 333940 46716 333946
rect 46664 333882 46716 333888
rect 45468 280220 45520 280226
rect 45468 280162 45520 280168
rect 44180 280152 44232 280158
rect 44180 280094 44232 280100
rect 45376 280152 45428 280158
rect 45376 280094 45428 280100
rect 44192 279478 44220 280094
rect 44180 279472 44232 279478
rect 44180 279414 44232 279420
rect 45376 269136 45428 269142
rect 45376 269078 45428 269084
rect 45388 199510 45416 269078
rect 45376 199504 45428 199510
rect 45376 199446 45428 199452
rect 45480 182918 45508 280162
rect 46756 269816 46808 269822
rect 46756 269758 46808 269764
rect 46768 191214 46796 269758
rect 46860 234598 46888 350542
rect 47964 339522 47992 393994
rect 48056 388482 48084 481646
rect 48148 458182 48176 556242
rect 48240 487830 48268 590650
rect 49608 586628 49660 586634
rect 49608 586570 49660 586576
rect 49516 585200 49568 585206
rect 49516 585142 49568 585148
rect 49424 496120 49476 496126
rect 49424 496062 49476 496068
rect 48964 491292 49016 491298
rect 48964 491234 49016 491240
rect 48228 487824 48280 487830
rect 48228 487766 48280 487772
rect 48228 472660 48280 472666
rect 48228 472602 48280 472608
rect 48136 458176 48188 458182
rect 48136 458118 48188 458124
rect 48044 388476 48096 388482
rect 48044 388418 48096 388424
rect 48044 387116 48096 387122
rect 48044 387058 48096 387064
rect 47952 339516 48004 339522
rect 47952 339458 48004 339464
rect 48056 338026 48084 387058
rect 48136 380316 48188 380322
rect 48136 380258 48188 380264
rect 48044 338020 48096 338026
rect 48044 337962 48096 337968
rect 48044 324964 48096 324970
rect 48044 324906 48096 324912
rect 48056 324358 48084 324906
rect 48044 324352 48096 324358
rect 48044 324294 48096 324300
rect 47952 277500 48004 277506
rect 47952 277442 48004 277448
rect 46848 234592 46900 234598
rect 46848 234534 46900 234540
rect 47964 222902 47992 277442
rect 48056 242894 48084 324294
rect 48148 310486 48176 380258
rect 48240 377466 48268 472602
rect 48976 387938 49004 491234
rect 49436 437374 49464 496062
rect 49528 493338 49556 585142
rect 49516 493332 49568 493338
rect 49516 493274 49568 493280
rect 49620 490618 49648 586570
rect 52368 586560 52420 586566
rect 52368 586502 52420 586508
rect 50712 585268 50764 585274
rect 50712 585210 50764 585216
rect 50724 492697 50752 585210
rect 50804 581188 50856 581194
rect 50804 581130 50856 581136
rect 50710 492688 50766 492697
rect 50710 492623 50766 492632
rect 50724 492114 50752 492623
rect 50712 492108 50764 492114
rect 50712 492050 50764 492056
rect 49608 490612 49660 490618
rect 49608 490554 49660 490560
rect 50816 485790 50844 581130
rect 52276 563100 52328 563106
rect 52276 563042 52328 563048
rect 52184 560992 52236 560998
rect 52184 560934 52236 560940
rect 50988 560312 51040 560318
rect 50988 560254 51040 560260
rect 50896 534880 50948 534886
rect 50896 534822 50948 534828
rect 50804 485784 50856 485790
rect 50804 485726 50856 485732
rect 49606 474736 49662 474745
rect 49606 474671 49662 474680
rect 49424 437368 49476 437374
rect 49424 437310 49476 437316
rect 49516 389836 49568 389842
rect 49516 389778 49568 389784
rect 48964 387932 49016 387938
rect 48964 387874 49016 387880
rect 48228 377460 48280 377466
rect 48228 377402 48280 377408
rect 48240 375426 48268 377402
rect 48228 375420 48280 375426
rect 48228 375362 48280 375368
rect 48228 363044 48280 363050
rect 48228 362986 48280 362992
rect 48136 310480 48188 310486
rect 48136 310422 48188 310428
rect 48148 309806 48176 310422
rect 48136 309800 48188 309806
rect 48136 309742 48188 309748
rect 48136 273284 48188 273290
rect 48136 273226 48188 273232
rect 48044 242888 48096 242894
rect 48044 242830 48096 242836
rect 47952 222896 48004 222902
rect 47952 222838 48004 222844
rect 48148 191282 48176 273226
rect 48240 264926 48268 362986
rect 49424 344344 49476 344350
rect 49424 344286 49476 344292
rect 49436 343670 49464 344286
rect 49424 343664 49476 343670
rect 49424 343606 49476 343612
rect 49436 304978 49464 343606
rect 49528 336734 49556 389778
rect 49620 380866 49648 474671
rect 50804 471300 50856 471306
rect 50804 471242 50856 471248
rect 50712 459604 50764 459610
rect 50712 459546 50764 459552
rect 50344 448588 50396 448594
rect 50344 448530 50396 448536
rect 50356 438530 50384 448530
rect 50344 438524 50396 438530
rect 50344 438466 50396 438472
rect 49608 380860 49660 380866
rect 49608 380802 49660 380808
rect 49620 380322 49648 380802
rect 49608 380316 49660 380322
rect 49608 380258 49660 380264
rect 49606 380216 49662 380225
rect 49606 380151 49662 380160
rect 49516 336728 49568 336734
rect 49516 336670 49568 336676
rect 49424 304972 49476 304978
rect 49424 304914 49476 304920
rect 49516 269204 49568 269210
rect 49516 269146 49568 269152
rect 48228 264920 48280 264926
rect 48228 264862 48280 264868
rect 48240 264246 48268 264862
rect 48228 264240 48280 264246
rect 48228 264182 48280 264188
rect 48228 262268 48280 262274
rect 48228 262210 48280 262216
rect 48136 191276 48188 191282
rect 48136 191218 48188 191224
rect 46756 191208 46808 191214
rect 46756 191150 46808 191156
rect 48240 185706 48268 262210
rect 49528 195362 49556 269146
rect 49620 231810 49648 380151
rect 50724 364342 50752 459546
rect 50816 400178 50844 471242
rect 50908 438870 50936 534822
rect 51000 460290 51028 560254
rect 52000 534948 52052 534954
rect 52000 534890 52052 534896
rect 50988 460284 51040 460290
rect 50988 460226 51040 460232
rect 51000 459610 51028 460226
rect 50988 459604 51040 459610
rect 50988 459546 51040 459552
rect 50896 438864 50948 438870
rect 50896 438806 50948 438812
rect 50908 438190 50936 438806
rect 50896 438184 50948 438190
rect 50896 438126 50948 438132
rect 52012 434722 52040 534890
rect 52092 532228 52144 532234
rect 52092 532170 52144 532176
rect 52104 440978 52132 532170
rect 52196 461650 52224 560934
rect 52288 463690 52316 563042
rect 52380 533390 52408 586502
rect 56508 583976 56560 583982
rect 56508 583918 56560 583924
rect 54942 583808 54998 583817
rect 54942 583743 54998 583752
rect 54484 582548 54536 582554
rect 54484 582490 54536 582496
rect 53104 581256 53156 581262
rect 53104 581198 53156 581204
rect 52368 533384 52420 533390
rect 52368 533326 52420 533332
rect 53116 483002 53144 581198
rect 53656 578264 53708 578270
rect 53656 578206 53708 578212
rect 53196 537600 53248 537606
rect 53196 537542 53248 537548
rect 53104 482996 53156 483002
rect 53104 482938 53156 482944
rect 52276 463684 52328 463690
rect 52276 463626 52328 463632
rect 53104 463684 53156 463690
rect 53104 463626 53156 463632
rect 52276 462324 52328 462330
rect 52276 462266 52328 462272
rect 52184 461644 52236 461650
rect 52184 461586 52236 461592
rect 52092 440972 52144 440978
rect 52092 440914 52144 440920
rect 52184 438728 52236 438734
rect 52184 438670 52236 438676
rect 52092 438184 52144 438190
rect 52092 438126 52144 438132
rect 52000 434716 52052 434722
rect 52000 434658 52052 434664
rect 50804 400172 50856 400178
rect 50804 400114 50856 400120
rect 50988 398880 51040 398886
rect 50988 398822 51040 398828
rect 50894 387696 50950 387705
rect 50894 387631 50950 387640
rect 50908 386578 50936 387631
rect 50896 386572 50948 386578
rect 50896 386514 50948 386520
rect 50804 385824 50856 385830
rect 50804 385766 50856 385772
rect 50816 385082 50844 385766
rect 50804 385076 50856 385082
rect 50804 385018 50856 385024
rect 50712 364336 50764 364342
rect 50712 364278 50764 364284
rect 50724 363050 50752 364278
rect 50712 363044 50764 363050
rect 50712 362986 50764 362992
rect 50816 284306 50844 385018
rect 50804 284300 50856 284306
rect 50804 284242 50856 284248
rect 50804 274712 50856 274718
rect 50804 274654 50856 274660
rect 50712 263628 50764 263634
rect 50712 263570 50764 263576
rect 49608 231804 49660 231810
rect 49608 231746 49660 231752
rect 50724 204950 50752 263570
rect 50712 204944 50764 204950
rect 50712 204886 50764 204892
rect 50816 200938 50844 274654
rect 50908 238746 50936 386514
rect 50896 238740 50948 238746
rect 50896 238682 50948 238688
rect 51000 237250 51028 398822
rect 51724 392012 51776 392018
rect 51724 391954 51776 391960
rect 51736 372570 51764 391954
rect 51724 372564 51776 372570
rect 51724 372506 51776 372512
rect 52104 339454 52132 438126
rect 52092 339448 52144 339454
rect 52092 339390 52144 339396
rect 52196 336666 52224 438670
rect 52288 437442 52316 462266
rect 53116 460934 53144 463626
rect 53208 462330 53236 537542
rect 53668 496806 53696 578206
rect 53748 537736 53800 537742
rect 53748 537678 53800 537684
rect 53656 496800 53708 496806
rect 53656 496742 53708 496748
rect 53656 496324 53708 496330
rect 53656 496266 53708 496272
rect 53196 462324 53248 462330
rect 53196 462266 53248 462272
rect 53116 460906 53328 460934
rect 53104 438320 53156 438326
rect 53104 438262 53156 438268
rect 52276 437436 52328 437442
rect 52276 437378 52328 437384
rect 53116 437238 53144 438262
rect 53104 437232 53156 437238
rect 53104 437174 53156 437180
rect 52460 391332 52512 391338
rect 52460 391274 52512 391280
rect 52472 390794 52500 391274
rect 52460 390788 52512 390794
rect 52460 390730 52512 390736
rect 52368 387932 52420 387938
rect 52368 387874 52420 387880
rect 52276 356108 52328 356114
rect 52276 356050 52328 356056
rect 52184 336660 52236 336666
rect 52184 336602 52236 336608
rect 52184 276072 52236 276078
rect 52184 276014 52236 276020
rect 51724 267708 51776 267714
rect 51724 267650 51776 267656
rect 50988 237244 51040 237250
rect 50988 237186 51040 237192
rect 50804 200932 50856 200938
rect 50804 200874 50856 200880
rect 49516 195356 49568 195362
rect 49516 195298 49568 195304
rect 48228 185700 48280 185706
rect 48228 185642 48280 185648
rect 45468 182912 45520 182918
rect 45468 182854 45520 182860
rect 51736 74526 51764 267650
rect 52196 198082 52224 276014
rect 52288 237318 52316 356050
rect 52380 267102 52408 387874
rect 53116 337890 53144 437174
rect 53300 402974 53328 460906
rect 53668 439550 53696 496266
rect 53656 439544 53708 439550
rect 53656 439486 53708 439492
rect 53760 438734 53788 537678
rect 54116 493400 54168 493406
rect 54114 493368 54116 493377
rect 54168 493368 54170 493377
rect 54114 493303 54170 493312
rect 53840 492788 53892 492794
rect 53840 492730 53892 492736
rect 53852 492182 53880 492730
rect 54496 492182 54524 582490
rect 54956 493406 54984 583743
rect 56324 574116 56376 574122
rect 56324 574058 56376 574064
rect 55036 552084 55088 552090
rect 55036 552026 55088 552032
rect 54944 493400 54996 493406
rect 54944 493342 54996 493348
rect 53840 492176 53892 492182
rect 53840 492118 53892 492124
rect 54484 492176 54536 492182
rect 54484 492118 54536 492124
rect 54852 491428 54904 491434
rect 54852 491370 54904 491376
rect 54864 454034 54892 491370
rect 54942 480312 54998 480321
rect 54942 480247 54998 480256
rect 54852 454028 54904 454034
rect 54852 453970 54904 453976
rect 54484 453348 54536 453354
rect 54484 453290 54536 453296
rect 53748 438728 53800 438734
rect 53748 438670 53800 438676
rect 53300 402946 53696 402974
rect 53668 393310 53696 402946
rect 53656 393304 53708 393310
rect 53656 393246 53708 393252
rect 53196 390788 53248 390794
rect 53196 390730 53248 390736
rect 53104 337884 53156 337890
rect 53104 337826 53156 337832
rect 53208 293282 53236 390730
rect 53668 369850 53696 393246
rect 53746 377768 53802 377777
rect 53746 377703 53802 377712
rect 53656 369844 53708 369850
rect 53656 369786 53708 369792
rect 53656 345092 53708 345098
rect 53656 345034 53708 345040
rect 53196 293276 53248 293282
rect 53196 293218 53248 293224
rect 53668 269074 53696 345034
rect 53760 339318 53788 377703
rect 53840 358080 53892 358086
rect 53840 358022 53892 358028
rect 53852 357474 53880 358022
rect 53840 357468 53892 357474
rect 53840 357410 53892 357416
rect 54496 356046 54524 453290
rect 54956 387870 54984 480247
rect 55048 453354 55076 552026
rect 55128 532160 55180 532166
rect 55128 532102 55180 532108
rect 55036 453348 55088 453354
rect 55036 453290 55088 453296
rect 55140 433226 55168 532102
rect 56140 491972 56192 491978
rect 56140 491914 56192 491920
rect 55956 475380 56008 475386
rect 55956 475322 56008 475328
rect 55968 474745 55996 475322
rect 55954 474736 56010 474745
rect 55954 474671 56010 474680
rect 55864 448588 55916 448594
rect 55864 448530 55916 448536
rect 55128 433220 55180 433226
rect 55128 433162 55180 433168
rect 55140 431954 55168 433162
rect 55048 431926 55168 431954
rect 54944 387864 54996 387870
rect 54944 387806 54996 387812
rect 54944 357468 54996 357474
rect 54944 357410 54996 357416
rect 54484 356040 54536 356046
rect 54484 355982 54536 355988
rect 53748 339312 53800 339318
rect 53748 339254 53800 339260
rect 53748 336660 53800 336666
rect 53748 336602 53800 336608
rect 53760 336054 53788 336602
rect 53748 336048 53800 336054
rect 53748 335990 53800 335996
rect 53656 269068 53708 269074
rect 53656 269010 53708 269016
rect 52368 267096 52420 267102
rect 52368 267038 52420 267044
rect 52460 262948 52512 262954
rect 52460 262890 52512 262896
rect 52472 262342 52500 262890
rect 53564 262880 53616 262886
rect 53564 262822 53616 262828
rect 52460 262336 52512 262342
rect 52460 262278 52512 262284
rect 52368 259480 52420 259486
rect 52368 259422 52420 259428
rect 52276 237312 52328 237318
rect 52276 237254 52328 237260
rect 52380 211818 52408 259422
rect 53380 255332 53432 255338
rect 53380 255274 53432 255280
rect 52368 211812 52420 211818
rect 52368 211754 52420 211760
rect 52184 198076 52236 198082
rect 52184 198018 52236 198024
rect 53392 192574 53420 255274
rect 53472 251252 53524 251258
rect 53472 251194 53524 251200
rect 53484 228478 53512 251194
rect 53472 228472 53524 228478
rect 53472 228414 53524 228420
rect 53576 210526 53604 262822
rect 53656 262336 53708 262342
rect 53656 262278 53708 262284
rect 53564 210520 53616 210526
rect 53564 210462 53616 210468
rect 53668 209098 53696 262278
rect 53760 253910 53788 335990
rect 54956 331906 54984 357410
rect 55048 339697 55076 431926
rect 55128 387864 55180 387870
rect 55128 387806 55180 387812
rect 55034 339688 55090 339697
rect 55034 339623 55090 339632
rect 55034 332072 55090 332081
rect 55034 332007 55036 332016
rect 55088 332007 55090 332016
rect 55036 331978 55088 331984
rect 54944 331900 54996 331906
rect 54944 331842 54996 331848
rect 54944 269068 54996 269074
rect 54944 269010 54996 269016
rect 54956 267034 54984 269010
rect 54944 267028 54996 267034
rect 54944 266970 54996 266976
rect 53748 253904 53800 253910
rect 53748 253846 53800 253852
rect 54852 248464 54904 248470
rect 54852 248406 54904 248412
rect 54484 242888 54536 242894
rect 54484 242830 54536 242836
rect 53656 209092 53708 209098
rect 53656 209034 53708 209040
rect 53380 192568 53432 192574
rect 53380 192510 53432 192516
rect 54496 192506 54524 242830
rect 54864 217394 54892 248406
rect 54956 218754 54984 266970
rect 55048 245614 55076 331978
rect 55140 280090 55168 387806
rect 55876 350538 55904 448530
rect 56152 439074 56180 491914
rect 56232 484356 56284 484362
rect 56232 484298 56284 484304
rect 56244 483682 56272 484298
rect 56232 483676 56284 483682
rect 56232 483618 56284 483624
rect 56140 439068 56192 439074
rect 56140 439010 56192 439016
rect 56244 398206 56272 483618
rect 56336 475386 56364 574058
rect 56416 547936 56468 547942
rect 56416 547878 56468 547884
rect 56324 475380 56376 475386
rect 56324 475322 56376 475328
rect 56428 449206 56456 547878
rect 56520 484362 56548 583918
rect 57796 582480 57848 582486
rect 57796 582422 57848 582428
rect 57704 564460 57756 564466
rect 57704 564402 57756 564408
rect 57520 537532 57572 537538
rect 57520 537474 57572 537480
rect 56508 484356 56560 484362
rect 56508 484298 56560 484304
rect 56508 455864 56560 455870
rect 56508 455806 56560 455812
rect 56416 449200 56468 449206
rect 56416 449142 56468 449148
rect 56428 448594 56456 449142
rect 56416 448588 56468 448594
rect 56416 448530 56468 448536
rect 56232 398200 56284 398206
rect 56232 398142 56284 398148
rect 56416 387252 56468 387258
rect 56416 387194 56468 387200
rect 56322 370560 56378 370569
rect 56322 370495 56378 370504
rect 55864 350532 55916 350538
rect 55864 350474 55916 350480
rect 56336 336462 56364 370495
rect 56428 339590 56456 387194
rect 56520 358086 56548 455806
rect 57532 436082 57560 537474
rect 57612 487212 57664 487218
rect 57612 487154 57664 487160
rect 57520 436076 57572 436082
rect 57520 436018 57572 436024
rect 57624 391338 57652 487154
rect 57716 465050 57744 564402
rect 57808 535022 57836 582422
rect 57900 554826 57928 697546
rect 58624 632120 58676 632126
rect 58624 632062 58676 632068
rect 57980 554872 58032 554878
rect 57900 554820 57980 554826
rect 57900 554814 58032 554820
rect 57900 554798 58020 554814
rect 57900 553466 57928 554798
rect 57900 553438 58020 553466
rect 57796 535016 57848 535022
rect 57796 534958 57848 534964
rect 57888 492788 57940 492794
rect 57888 492730 57940 492736
rect 57796 487824 57848 487830
rect 57796 487766 57848 487772
rect 57808 487218 57836 487766
rect 57796 487212 57848 487218
rect 57796 487154 57848 487160
rect 57704 465044 57756 465050
rect 57704 464986 57756 464992
rect 57704 394120 57756 394126
rect 57704 394062 57756 394068
rect 57612 391332 57664 391338
rect 57612 391274 57664 391280
rect 57242 390552 57298 390561
rect 57242 390487 57298 390496
rect 57256 389298 57284 390487
rect 57244 389292 57296 389298
rect 57244 389234 57296 389240
rect 57612 389292 57664 389298
rect 57612 389234 57664 389240
rect 56508 358080 56560 358086
rect 56508 358022 56560 358028
rect 56416 339584 56468 339590
rect 56416 339526 56468 339532
rect 56324 336456 56376 336462
rect 56324 336398 56376 336404
rect 56416 334008 56468 334014
rect 56416 333950 56468 333956
rect 55128 280084 55180 280090
rect 55128 280026 55180 280032
rect 55128 274780 55180 274786
rect 55128 274722 55180 274728
rect 55036 245608 55088 245614
rect 55036 245550 55088 245556
rect 55140 224398 55168 274722
rect 56324 258120 56376 258126
rect 56324 258062 56376 258068
rect 56232 253224 56284 253230
rect 56232 253166 56284 253172
rect 56244 252618 56272 253166
rect 56232 252612 56284 252618
rect 56232 252554 56284 252560
rect 56244 232558 56272 252554
rect 56232 232552 56284 232558
rect 56232 232494 56284 232500
rect 55128 224392 55180 224398
rect 55128 224334 55180 224340
rect 54944 218748 54996 218754
rect 54944 218690 54996 218696
rect 54852 217388 54904 217394
rect 54852 217330 54904 217336
rect 56336 195498 56364 258062
rect 56428 238678 56456 333950
rect 56520 303618 56548 358022
rect 56508 303612 56560 303618
rect 56508 303554 56560 303560
rect 57242 292904 57298 292913
rect 57242 292839 57298 292848
rect 56508 280288 56560 280294
rect 56508 280230 56560 280236
rect 56416 238672 56468 238678
rect 56416 238614 56468 238620
rect 56324 195492 56376 195498
rect 56324 195434 56376 195440
rect 54484 192500 54536 192506
rect 54484 192442 54536 192448
rect 56520 181558 56548 280230
rect 56508 181552 56560 181558
rect 56508 181494 56560 181500
rect 51724 74520 51776 74526
rect 51724 74462 51776 74468
rect 46940 62892 46992 62898
rect 46940 62834 46992 62840
rect 45560 40792 45612 40798
rect 45560 40734 45612 40740
rect 44180 31136 44232 31142
rect 44180 31078 44232 31084
rect 43444 23452 43496 23458
rect 43444 23394 43496 23400
rect 44088 23452 44140 23458
rect 44088 23394 44140 23400
rect 41432 16546 41920 16574
rect 41328 2236 41380 2242
rect 41328 2178 41380 2184
rect 41892 480 41920 16546
rect 43456 7614 43484 23394
rect 44192 16574 44220 31078
rect 45572 16574 45600 40734
rect 46952 16574 46980 62834
rect 49698 57216 49754 57225
rect 49698 57151 49754 57160
rect 48320 24132 48372 24138
rect 48320 24074 48372 24080
rect 48332 16574 48360 24074
rect 49712 16574 49740 57151
rect 51736 33114 51764 74462
rect 53840 61396 53892 61402
rect 53840 61338 53892 61344
rect 51724 33108 51776 33114
rect 51724 33050 51776 33056
rect 52460 29708 52512 29714
rect 52460 29650 52512 29656
rect 51080 26920 51132 26926
rect 51080 26862 51132 26868
rect 44192 16546 44312 16574
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 43444 7608 43496 7614
rect 43444 7550 43496 7556
rect 43076 4888 43128 4894
rect 43076 4830 43128 4836
rect 43088 480 43116 4830
rect 44284 480 44312 16546
rect 45468 7608 45520 7614
rect 45468 7550 45520 7556
rect 45480 480 45508 7550
rect 46676 480 46704 16546
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 26862
rect 52472 6914 52500 29650
rect 52552 22772 52604 22778
rect 52552 22714 52604 22720
rect 52564 16574 52592 22714
rect 53852 16574 53880 61338
rect 57256 20670 57284 292839
rect 57624 255270 57652 389234
rect 57716 336530 57744 394062
rect 57900 393314 57928 492730
rect 57992 455870 58020 553438
rect 58636 539510 58664 632062
rect 61936 585336 61988 585342
rect 61936 585278 61988 585284
rect 59176 583840 59228 583846
rect 59176 583782 59228 583788
rect 58624 539504 58676 539510
rect 58624 539446 58676 539452
rect 59188 498166 59216 583782
rect 60004 583024 60056 583030
rect 60004 582966 60056 582972
rect 59268 560380 59320 560386
rect 59268 560322 59320 560328
rect 59176 498160 59228 498166
rect 59176 498102 59228 498108
rect 59188 497690 59216 498102
rect 59176 497684 59228 497690
rect 59176 497626 59228 497632
rect 58072 496800 58124 496806
rect 58072 496742 58124 496748
rect 58084 481545 58112 496742
rect 58992 490680 59044 490686
rect 58992 490622 59044 490628
rect 58070 481536 58126 481545
rect 58070 481471 58126 481480
rect 57980 455864 58032 455870
rect 57980 455806 58032 455812
rect 57992 455394 58020 455806
rect 57980 455388 58032 455394
rect 57980 455330 58032 455336
rect 59004 437238 59032 490622
rect 59174 481536 59230 481545
rect 59174 481471 59230 481480
rect 59188 480321 59216 481471
rect 59174 480312 59230 480321
rect 59174 480247 59230 480256
rect 59188 480214 59216 480247
rect 59176 480208 59228 480214
rect 59176 480150 59228 480156
rect 59084 470620 59136 470626
rect 59084 470562 59136 470568
rect 58992 437232 59044 437238
rect 58992 437174 59044 437180
rect 57808 393286 57928 393314
rect 57808 389366 57836 393286
rect 57796 389360 57848 389366
rect 57796 389302 57848 389308
rect 57704 336524 57756 336530
rect 57704 336466 57756 336472
rect 57808 294098 57836 389302
rect 58530 388376 58586 388385
rect 58530 388311 58586 388320
rect 58544 388006 58572 388311
rect 58532 388000 58584 388006
rect 58532 387942 58584 387948
rect 59096 378049 59124 470562
rect 59176 462324 59228 462330
rect 59176 462266 59228 462272
rect 59188 461650 59216 462266
rect 59280 462262 59308 560322
rect 60016 538286 60044 582966
rect 61752 574184 61804 574190
rect 61752 574126 61804 574132
rect 60464 563168 60516 563174
rect 60464 563110 60516 563116
rect 60004 538280 60056 538286
rect 60004 538222 60056 538228
rect 60372 467900 60424 467906
rect 60372 467842 60424 467848
rect 59268 462256 59320 462262
rect 59268 462198 59320 462204
rect 59176 461644 59228 461650
rect 59176 461586 59228 461592
rect 59082 378040 59138 378049
rect 59082 377975 59138 377984
rect 59188 366382 59216 461586
rect 59268 439068 59320 439074
rect 59268 439010 59320 439016
rect 59176 366376 59228 366382
rect 59176 366318 59228 366324
rect 59084 362976 59136 362982
rect 59084 362918 59136 362924
rect 59096 361554 59124 362918
rect 59084 361548 59136 361554
rect 59084 361490 59136 361496
rect 59084 359508 59136 359514
rect 59084 359450 59136 359456
rect 59096 358834 59124 359450
rect 59084 358828 59136 358834
rect 59084 358770 59136 358776
rect 57888 347812 57940 347818
rect 57888 347754 57940 347760
rect 57900 347721 57928 347754
rect 57886 347712 57942 347721
rect 57886 347647 57942 347656
rect 58990 338056 59046 338065
rect 58990 337991 59046 338000
rect 59004 337482 59032 337991
rect 58992 337476 59044 337482
rect 58992 337418 59044 337424
rect 57796 294092 57848 294098
rect 57796 294034 57848 294040
rect 57808 291854 57836 294034
rect 57796 291848 57848 291854
rect 57796 291790 57848 291796
rect 57888 260908 57940 260914
rect 57888 260850 57940 260856
rect 57796 258188 57848 258194
rect 57796 258130 57848 258136
rect 57612 255264 57664 255270
rect 57612 255206 57664 255212
rect 57704 249076 57756 249082
rect 57704 249018 57756 249024
rect 57716 248538 57744 249018
rect 57704 248532 57756 248538
rect 57704 248474 57756 248480
rect 57716 218822 57744 248474
rect 57704 218816 57756 218822
rect 57704 218758 57756 218764
rect 57808 196790 57836 258130
rect 57900 228546 57928 260850
rect 58624 254584 58676 254590
rect 58624 254526 58676 254532
rect 58636 238814 58664 254526
rect 58624 238808 58676 238814
rect 58624 238750 58676 238756
rect 59004 237182 59032 337418
rect 59096 305794 59124 358770
rect 59188 334694 59216 366318
rect 59280 334762 59308 439010
rect 60384 373998 60412 467842
rect 60476 463826 60504 563110
rect 60740 562352 60792 562358
rect 60740 562294 60792 562300
rect 60752 560998 60780 562294
rect 60740 560992 60792 560998
rect 60740 560934 60792 560940
rect 61660 546576 61712 546582
rect 61660 546518 61712 546524
rect 60556 546508 60608 546514
rect 60556 546450 60608 546456
rect 60464 463820 60516 463826
rect 60464 463762 60516 463768
rect 60464 463684 60516 463690
rect 60464 463626 60516 463632
rect 60372 373992 60424 373998
rect 60372 373934 60424 373940
rect 60372 367804 60424 367810
rect 60372 367746 60424 367752
rect 60004 356108 60056 356114
rect 60004 356050 60056 356056
rect 60016 355978 60044 356050
rect 60004 355972 60056 355978
rect 60004 355914 60056 355920
rect 59268 334756 59320 334762
rect 59268 334698 59320 334704
rect 59176 334688 59228 334694
rect 59176 334630 59228 334636
rect 60016 316810 60044 355914
rect 60384 339250 60412 367746
rect 60476 367062 60504 463626
rect 60568 445806 60596 546450
rect 60648 541000 60700 541006
rect 60648 540942 60700 540948
rect 60556 445800 60608 445806
rect 60556 445742 60608 445748
rect 60660 441590 60688 540942
rect 61384 449948 61436 449954
rect 61384 449890 61436 449896
rect 60648 441584 60700 441590
rect 60648 441526 60700 441532
rect 60648 392692 60700 392698
rect 60648 392634 60700 392640
rect 60556 371884 60608 371890
rect 60556 371826 60608 371832
rect 60464 367056 60516 367062
rect 60464 366998 60516 367004
rect 60372 339244 60424 339250
rect 60372 339186 60424 339192
rect 60568 335306 60596 371826
rect 60556 335300 60608 335306
rect 60556 335242 60608 335248
rect 60568 334014 60596 335242
rect 60556 334008 60608 334014
rect 60556 333950 60608 333956
rect 60660 333878 60688 392634
rect 61396 352646 61424 449890
rect 61672 447234 61700 546518
rect 61764 477494 61792 574126
rect 61844 561740 61896 561746
rect 61844 561682 61896 561688
rect 61752 477488 61804 477494
rect 61752 477430 61804 477436
rect 61752 466812 61804 466818
rect 61752 466754 61804 466760
rect 61660 447228 61712 447234
rect 61660 447170 61712 447176
rect 61764 402974 61792 466754
rect 61856 463690 61884 561682
rect 61948 541686 61976 585278
rect 62040 562358 62068 700266
rect 68836 596828 68888 596834
rect 68836 596770 68888 596776
rect 68652 592680 68704 592686
rect 68652 592622 68704 592628
rect 66168 584044 66220 584050
rect 66168 583986 66220 583992
rect 65524 581800 65576 581806
rect 65524 581742 65576 581748
rect 65536 581058 65564 581742
rect 65524 581052 65576 581058
rect 65524 580994 65576 581000
rect 65524 579692 65576 579698
rect 65524 579634 65576 579640
rect 64604 578332 64656 578338
rect 64604 578274 64656 578280
rect 64512 576904 64564 576910
rect 64512 576846 64564 576852
rect 63224 569968 63276 569974
rect 63224 569910 63276 569916
rect 63132 565888 63184 565894
rect 63132 565830 63184 565836
rect 62028 562352 62080 562358
rect 62028 562294 62080 562300
rect 61936 541680 61988 541686
rect 61936 541622 61988 541628
rect 62028 539640 62080 539646
rect 62028 539582 62080 539588
rect 61844 463684 61896 463690
rect 61844 463626 61896 463632
rect 61936 442944 61988 442950
rect 61936 442886 61988 442892
rect 61844 403028 61896 403034
rect 61844 402974 61896 402976
rect 61764 402970 61896 402974
rect 61764 402946 61884 402970
rect 61856 372570 61884 402946
rect 61844 372564 61896 372570
rect 61844 372506 61896 372512
rect 61384 352640 61436 352646
rect 61384 352582 61436 352588
rect 61396 351966 61424 352582
rect 61384 351960 61436 351966
rect 61384 351902 61436 351908
rect 61844 351960 61896 351966
rect 61844 351902 61896 351908
rect 60648 333872 60700 333878
rect 60648 333814 60700 333820
rect 61856 333334 61884 351902
rect 61948 342310 61976 442886
rect 62040 441046 62068 539582
rect 63040 477624 63092 477630
rect 63040 477566 63092 477572
rect 63052 471306 63080 477566
rect 63040 471300 63092 471306
rect 63040 471242 63092 471248
rect 63144 466818 63172 565830
rect 63236 477630 63264 569910
rect 63316 567248 63368 567254
rect 63316 567190 63368 567196
rect 63224 477624 63276 477630
rect 63224 477566 63276 477572
rect 63224 477488 63276 477494
rect 63222 477456 63224 477465
rect 63276 477456 63278 477465
rect 63222 477391 63278 477400
rect 63328 467906 63356 567190
rect 63408 542496 63460 542502
rect 63408 542438 63460 542444
rect 63316 467900 63368 467906
rect 63316 467842 63368 467848
rect 63132 466812 63184 466818
rect 63132 466754 63184 466760
rect 63224 462256 63276 462262
rect 63224 462198 63276 462204
rect 63236 460970 63264 462198
rect 63224 460964 63276 460970
rect 63224 460906 63276 460912
rect 62764 451240 62816 451246
rect 62764 451182 62816 451188
rect 62028 441040 62080 441046
rect 62028 440982 62080 440988
rect 61936 342304 61988 342310
rect 61936 342246 61988 342252
rect 62040 340202 62068 440982
rect 62776 353326 62804 451182
rect 63132 383784 63184 383790
rect 63132 383726 63184 383732
rect 62764 353320 62816 353326
rect 62764 353262 62816 353268
rect 62028 340196 62080 340202
rect 62028 340138 62080 340144
rect 62028 334756 62080 334762
rect 62028 334698 62080 334704
rect 61844 333328 61896 333334
rect 61844 333270 61896 333276
rect 60004 316804 60056 316810
rect 60004 316746 60056 316752
rect 59084 305788 59136 305794
rect 59084 305730 59136 305736
rect 60648 304292 60700 304298
rect 60648 304234 60700 304240
rect 59268 300144 59320 300150
rect 59268 300086 59320 300092
rect 59176 267096 59228 267102
rect 59176 267038 59228 267044
rect 59188 266422 59216 267038
rect 59176 266416 59228 266422
rect 59176 266358 59228 266364
rect 59188 258074 59216 266358
rect 59280 266354 59308 300086
rect 59268 266348 59320 266354
rect 59268 266290 59320 266296
rect 60556 264988 60608 264994
rect 60556 264930 60608 264936
rect 59096 258046 59216 258074
rect 58992 237176 59044 237182
rect 58992 237118 59044 237124
rect 57888 228540 57940 228546
rect 57888 228482 57940 228488
rect 59096 217326 59124 258046
rect 59268 256760 59320 256766
rect 59268 256702 59320 256708
rect 59084 217320 59136 217326
rect 59084 217262 59136 217268
rect 57796 196784 57848 196790
rect 57796 196726 57848 196732
rect 59280 189854 59308 256702
rect 60004 253904 60056 253910
rect 60004 253846 60056 253852
rect 60016 229770 60044 253846
rect 60464 249824 60516 249830
rect 60464 249766 60516 249772
rect 60476 235346 60504 249766
rect 60568 236609 60596 264930
rect 60660 260846 60688 304234
rect 61936 267844 61988 267850
rect 61936 267786 61988 267792
rect 60648 260840 60700 260846
rect 60648 260782 60700 260788
rect 61844 251320 61896 251326
rect 61844 251262 61896 251268
rect 60648 247104 60700 247110
rect 60648 247046 60700 247052
rect 60554 236600 60610 236609
rect 60554 236535 60610 236544
rect 60464 235340 60516 235346
rect 60464 235282 60516 235288
rect 60004 229764 60056 229770
rect 60004 229706 60056 229712
rect 60660 207738 60688 247046
rect 61384 245676 61436 245682
rect 61384 245618 61436 245624
rect 61396 221542 61424 245618
rect 61856 234122 61884 251262
rect 61948 239494 61976 267786
rect 62040 244254 62068 334698
rect 62028 244248 62080 244254
rect 62028 244190 62080 244196
rect 62028 241528 62080 241534
rect 62028 241470 62080 241476
rect 61936 239488 61988 239494
rect 61936 239430 61988 239436
rect 61844 234116 61896 234122
rect 61844 234058 61896 234064
rect 61384 221536 61436 221542
rect 61384 221478 61436 221484
rect 62040 211954 62068 241470
rect 62028 211948 62080 211954
rect 62028 211890 62080 211896
rect 60648 207732 60700 207738
rect 60648 207674 60700 207680
rect 59268 189848 59320 189854
rect 59268 189790 59320 189796
rect 59268 127016 59320 127022
rect 59268 126958 59320 126964
rect 59280 93673 59308 126958
rect 59266 93664 59322 93673
rect 59266 93599 59322 93608
rect 63144 73166 63172 383726
rect 63236 365702 63264 460906
rect 63314 448624 63370 448633
rect 63314 448559 63370 448568
rect 63224 365696 63276 365702
rect 63224 365638 63276 365644
rect 63328 351218 63356 448559
rect 63420 442950 63448 542438
rect 64524 480185 64552 576846
rect 64616 481642 64644 578274
rect 64696 567316 64748 567322
rect 64696 567258 64748 567264
rect 64604 481636 64656 481642
rect 64604 481578 64656 481584
rect 64510 480176 64566 480185
rect 64510 480111 64566 480120
rect 64236 474700 64288 474706
rect 64236 474642 64288 474648
rect 64144 463820 64196 463826
rect 64144 463762 64196 463768
rect 63408 442944 63460 442950
rect 63408 442886 63460 442892
rect 64156 368393 64184 463762
rect 64248 379574 64276 474642
rect 64512 469532 64564 469538
rect 64512 469474 64564 469480
rect 64236 379568 64288 379574
rect 64236 379510 64288 379516
rect 64524 374678 64552 469474
rect 64708 469130 64736 567258
rect 64788 548004 64840 548010
rect 64788 547946 64840 547952
rect 64696 469124 64748 469130
rect 64696 469066 64748 469072
rect 64800 447166 64828 547946
rect 65536 481710 65564 579634
rect 66076 571600 66128 571606
rect 66076 571542 66128 571548
rect 65616 553444 65668 553450
rect 65616 553386 65668 553392
rect 65628 491434 65656 553386
rect 65616 491428 65668 491434
rect 65616 491370 65668 491376
rect 65984 491428 66036 491434
rect 65984 491370 66036 491376
rect 65996 490521 66024 491370
rect 65982 490512 66038 490521
rect 65982 490447 66038 490456
rect 65616 485852 65668 485858
rect 65616 485794 65668 485800
rect 65524 481704 65576 481710
rect 65524 481646 65576 481652
rect 64970 477592 65026 477601
rect 64970 477527 65026 477536
rect 64984 471646 65012 477527
rect 64972 471640 65024 471646
rect 64972 471582 65024 471588
rect 64984 470626 65012 471582
rect 64972 470620 65024 470626
rect 64972 470562 65024 470568
rect 65524 465112 65576 465118
rect 65524 465054 65576 465060
rect 64788 447160 64840 447166
rect 64788 447102 64840 447108
rect 64604 445800 64656 445806
rect 64604 445742 64656 445748
rect 64512 374672 64564 374678
rect 64512 374614 64564 374620
rect 64142 368384 64198 368393
rect 64142 368319 64198 368328
rect 63316 351212 63368 351218
rect 63316 351154 63368 351160
rect 63316 349172 63368 349178
rect 63316 349114 63368 349120
rect 63328 330585 63356 349114
rect 64616 347070 64644 445742
rect 64786 380216 64842 380225
rect 64786 380151 64842 380160
rect 64800 378185 64828 380151
rect 64786 378176 64842 378185
rect 64786 378111 64842 378120
rect 64788 374672 64840 374678
rect 64788 374614 64840 374620
rect 64696 365696 64748 365702
rect 64696 365638 64748 365644
rect 64708 364410 64736 365638
rect 64696 364404 64748 364410
rect 64696 364346 64748 364352
rect 64604 347064 64656 347070
rect 64604 347006 64656 347012
rect 63314 330576 63370 330585
rect 63314 330511 63370 330520
rect 63316 276140 63368 276146
rect 63316 276082 63368 276088
rect 63224 247172 63276 247178
rect 63224 247114 63276 247120
rect 63236 235414 63264 247114
rect 63224 235408 63276 235414
rect 63224 235350 63276 235356
rect 63328 188358 63356 276082
rect 64512 271924 64564 271930
rect 64512 271866 64564 271872
rect 63408 245744 63460 245750
rect 63408 245686 63460 245692
rect 63420 239562 63448 245686
rect 63408 239556 63460 239562
rect 63408 239498 63460 239504
rect 64524 225690 64552 271866
rect 64512 225684 64564 225690
rect 64512 225626 64564 225632
rect 63316 188352 63368 188358
rect 63316 188294 63368 188300
rect 63132 73160 63184 73166
rect 63132 73102 63184 73108
rect 57980 43444 58032 43450
rect 57980 43386 58032 43392
rect 57244 20664 57296 20670
rect 57244 20606 57296 20612
rect 56600 19984 56652 19990
rect 56600 19926 56652 19932
rect 56612 16574 56640 19926
rect 57992 16574 58020 43386
rect 59360 39432 59412 39438
rect 59360 39374 59412 39380
rect 52564 16546 53328 16574
rect 53852 16546 54984 16574
rect 56612 16546 56824 16574
rect 57992 16546 58480 16574
rect 52472 6886 52592 6914
rect 52564 480 52592 6886
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53300 354 53328 16546
rect 54956 480 54984 16546
rect 56048 13116 56100 13122
rect 56048 13058 56100 13064
rect 56060 480 56088 13058
rect 53718 354 53830 480
rect 53300 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58452 480 58480 16546
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 39374
rect 60740 33788 60792 33794
rect 60740 33730 60792 33736
rect 60752 16574 60780 33730
rect 62120 32428 62172 32434
rect 62120 32370 62172 32376
rect 62132 16574 62160 32370
rect 64616 20670 64644 347006
rect 64708 37262 64736 364346
rect 64696 37256 64748 37262
rect 64696 37198 64748 37204
rect 64800 29646 64828 374614
rect 65536 370190 65564 465054
rect 65628 436762 65656 485794
rect 65984 481704 66036 481710
rect 65984 481646 66036 481652
rect 65996 481574 66024 481646
rect 65984 481568 66036 481574
rect 65984 481510 66036 481516
rect 66088 473346 66116 571542
rect 66180 571334 66208 583986
rect 68468 582004 68520 582010
rect 68468 581946 68520 581952
rect 67638 581360 67694 581369
rect 67638 581295 67694 581304
rect 67652 581262 67680 581295
rect 67640 581256 67692 581262
rect 67640 581198 67692 581204
rect 67730 579184 67786 579193
rect 67730 579119 67786 579128
rect 67638 578504 67694 578513
rect 67638 578439 67694 578448
rect 67652 578270 67680 578439
rect 67744 578338 67772 579119
rect 67732 578332 67784 578338
rect 67732 578274 67784 578280
rect 67640 578264 67692 578270
rect 67640 578206 67692 578212
rect 67638 577824 67694 577833
rect 67638 577759 67694 577768
rect 67546 577144 67602 577153
rect 67546 577079 67602 577088
rect 67454 572792 67510 572801
rect 67454 572727 67510 572736
rect 66168 571328 66220 571334
rect 66168 571270 66220 571276
rect 66168 568608 66220 568614
rect 66168 568550 66220 568556
rect 66076 473340 66128 473346
rect 66076 473282 66128 473288
rect 66088 472666 66116 473282
rect 66076 472660 66128 472666
rect 66076 472602 66128 472608
rect 66074 470520 66130 470529
rect 66074 470455 66130 470464
rect 66088 469266 66116 470455
rect 66180 469538 66208 568550
rect 67362 564496 67418 564505
rect 67362 564431 67418 564440
rect 67272 484628 67324 484634
rect 67272 484570 67324 484576
rect 66168 469532 66220 469538
rect 66168 469474 66220 469480
rect 66076 469260 66128 469266
rect 66076 469202 66128 469208
rect 66076 469124 66128 469130
rect 66076 469066 66128 469072
rect 66088 468246 66116 469066
rect 66076 468240 66128 468246
rect 66076 468182 66128 468188
rect 65616 436756 65668 436762
rect 65616 436698 65668 436704
rect 65890 383888 65946 383897
rect 65890 383823 65946 383832
rect 65904 383790 65932 383823
rect 65892 383784 65944 383790
rect 65892 383726 65944 383732
rect 65984 379568 66036 379574
rect 65984 379510 66036 379516
rect 65892 373992 65944 373998
rect 65890 373960 65892 373969
rect 65944 373960 65946 373969
rect 65890 373895 65946 373904
rect 65524 370184 65576 370190
rect 65524 370126 65576 370132
rect 65996 326398 66024 379510
rect 66088 371958 66116 468182
rect 66260 447228 66312 447234
rect 66260 447170 66312 447176
rect 66168 447160 66220 447166
rect 66168 447102 66220 447108
rect 66076 371952 66128 371958
rect 66076 371894 66128 371900
rect 66088 331809 66116 371894
rect 66180 349790 66208 447102
rect 66168 349784 66220 349790
rect 66168 349726 66220 349732
rect 66272 349178 66300 447170
rect 67284 439618 67312 484570
rect 67376 466454 67404 564431
rect 67468 474337 67496 572727
rect 67560 478553 67588 577079
rect 67652 576910 67680 577759
rect 67640 576904 67692 576910
rect 67640 576846 67692 576852
rect 67638 575784 67694 575793
rect 67638 575719 67694 575728
rect 67652 575550 67680 575719
rect 67640 575544 67692 575550
rect 67640 575486 67692 575492
rect 67730 575104 67786 575113
rect 67730 575039 67786 575048
rect 67638 574424 67694 574433
rect 67638 574359 67694 574368
rect 67652 574122 67680 574359
rect 67744 574190 67772 575039
rect 67732 574184 67784 574190
rect 67732 574126 67784 574132
rect 67640 574116 67692 574122
rect 67640 574058 67692 574064
rect 67638 573472 67694 573481
rect 67638 573407 67694 573416
rect 67652 572830 67680 573407
rect 67640 572824 67692 572830
rect 67640 572766 67692 572772
rect 68480 571713 68508 581946
rect 68664 580689 68692 592622
rect 68650 580680 68706 580689
rect 68650 580615 68706 580624
rect 68664 579698 68692 580615
rect 68652 579692 68704 579698
rect 68652 579634 68704 579640
rect 68848 579614 68876 596770
rect 68756 579586 68876 579614
rect 68650 576464 68706 576473
rect 68650 576399 68706 576408
rect 68282 571704 68338 571713
rect 68282 571639 68338 571648
rect 68466 571704 68522 571713
rect 68466 571639 68522 571648
rect 68296 571606 68324 571639
rect 68284 571600 68336 571606
rect 68284 571542 68336 571548
rect 68284 571328 68336 571334
rect 68284 571270 68336 571276
rect 67638 570072 67694 570081
rect 67638 570007 67694 570016
rect 67652 569974 67680 570007
rect 67640 569968 67692 569974
rect 67640 569910 67692 569916
rect 67638 568712 67694 568721
rect 67638 568647 67694 568656
rect 67652 568614 67680 568647
rect 67640 568608 67692 568614
rect 67640 568550 67692 568556
rect 67730 567624 67786 567633
rect 67730 567559 67786 567568
rect 67640 567316 67692 567322
rect 67640 567258 67692 567264
rect 67652 567225 67680 567258
rect 67744 567254 67772 567559
rect 67732 567248 67784 567254
rect 67638 567216 67694 567225
rect 67732 567190 67784 567196
rect 67638 567151 67694 567160
rect 67638 566264 67694 566273
rect 67638 566199 67694 566208
rect 67652 565894 67680 566199
rect 67640 565888 67692 565894
rect 67640 565830 67692 565836
rect 67638 564904 67694 564913
rect 67638 564839 67694 564848
rect 67652 564466 67680 564839
rect 67640 564460 67692 564466
rect 67640 564402 67692 564408
rect 67730 563544 67786 563553
rect 67730 563479 67786 563488
rect 67640 563168 67692 563174
rect 67638 563136 67640 563145
rect 67692 563136 67694 563145
rect 67744 563106 67772 563479
rect 67638 563071 67694 563080
rect 67732 563100 67784 563106
rect 67732 563042 67784 563048
rect 67640 562352 67692 562358
rect 67638 562320 67640 562329
rect 67692 562320 67694 562329
rect 67638 562255 67694 562264
rect 67638 562184 67694 562193
rect 67638 562119 67694 562128
rect 67652 561746 67680 562119
rect 67640 561740 67692 561746
rect 67640 561682 67692 561688
rect 67730 560824 67786 560833
rect 67730 560759 67786 560768
rect 67638 560416 67694 560425
rect 67744 560386 67772 560759
rect 67638 560351 67694 560360
rect 67732 560380 67784 560386
rect 67652 560318 67680 560351
rect 67732 560322 67784 560328
rect 67640 560312 67692 560318
rect 67640 560254 67692 560260
rect 67638 559464 67694 559473
rect 67638 559399 67694 559408
rect 67652 558958 67680 559399
rect 67640 558952 67692 558958
rect 67640 558894 67692 558900
rect 67640 557592 67692 557598
rect 67638 557560 67640 557569
rect 67692 557560 67694 557569
rect 67638 557495 67694 557504
rect 68296 557433 68324 571270
rect 68282 557424 68338 557433
rect 68282 557359 68338 557368
rect 67730 556744 67786 556753
rect 67730 556679 67786 556688
rect 67640 556300 67692 556306
rect 67640 556242 67692 556248
rect 67652 556209 67680 556242
rect 67744 556238 67772 556679
rect 67732 556232 67784 556238
rect 67638 556200 67694 556209
rect 67732 556174 67784 556180
rect 67638 556135 67694 556144
rect 67730 555384 67786 555393
rect 67730 555319 67786 555328
rect 67640 554872 67692 554878
rect 67638 554840 67640 554849
rect 67692 554840 67694 554849
rect 67744 554810 67772 555319
rect 67638 554775 67694 554784
rect 67732 554804 67784 554810
rect 67732 554746 67784 554752
rect 67638 553480 67694 553489
rect 67638 553415 67640 553424
rect 67692 553415 67694 553424
rect 67640 553386 67692 553392
rect 67638 552120 67694 552129
rect 67638 552055 67640 552064
rect 67692 552055 67694 552064
rect 67640 552026 67692 552032
rect 67638 551304 67694 551313
rect 67638 551239 67694 551248
rect 67652 550662 67680 551239
rect 67640 550656 67692 550662
rect 67640 550598 67692 550604
rect 67638 549944 67694 549953
rect 67638 549879 67694 549888
rect 67652 549302 67680 549879
rect 67640 549296 67692 549302
rect 67640 549238 67692 549244
rect 67730 548584 67786 548593
rect 67730 548519 67786 548528
rect 67638 548040 67694 548049
rect 67638 547975 67640 547984
rect 67692 547975 67694 547984
rect 67640 547946 67692 547952
rect 67744 547942 67772 548519
rect 67732 547936 67784 547942
rect 67732 547878 67784 547884
rect 67730 547224 67786 547233
rect 67730 547159 67786 547168
rect 67744 546582 67772 547159
rect 67732 546576 67784 546582
rect 67638 546544 67694 546553
rect 67732 546518 67784 546524
rect 67638 546479 67640 546488
rect 67692 546479 67694 546488
rect 67640 546450 67692 546456
rect 68098 545320 68154 545329
rect 68098 545255 68154 545264
rect 68112 545154 68140 545255
rect 68100 545148 68152 545154
rect 68100 545090 68152 545096
rect 68008 544400 68060 544406
rect 68008 544342 68060 544348
rect 68020 543969 68048 544342
rect 68006 543960 68062 543969
rect 68006 543895 68062 543904
rect 68006 543280 68062 543289
rect 68006 543215 68062 543224
rect 67638 542600 67694 542609
rect 67638 542535 67694 542544
rect 67652 542502 67680 542535
rect 67640 542496 67692 542502
rect 67640 542438 67692 542444
rect 68020 542434 68048 543215
rect 68008 542428 68060 542434
rect 68008 542370 68060 542376
rect 67638 541240 67694 541249
rect 67638 541175 67694 541184
rect 67652 541006 67680 541175
rect 67640 541000 67692 541006
rect 67640 540942 67692 540948
rect 67638 540152 67694 540161
rect 67638 540087 67694 540096
rect 67652 539646 67680 540087
rect 67640 539640 67692 539646
rect 67640 539582 67692 539588
rect 68664 489914 68692 576399
rect 68756 569954 68784 579586
rect 68940 572529 68968 702442
rect 71044 700392 71096 700398
rect 71044 700334 71096 700340
rect 69020 696992 69072 696998
rect 69020 696934 69072 696940
rect 68926 572520 68982 572529
rect 68926 572455 68982 572464
rect 68940 571849 68968 572455
rect 68926 571840 68982 571849
rect 68926 571775 68982 571784
rect 68756 569926 68876 569954
rect 68848 558929 68876 569926
rect 68834 558920 68890 558929
rect 68834 558855 68890 558864
rect 68848 558210 68876 558855
rect 68836 558204 68888 558210
rect 68836 558146 68888 558152
rect 68834 550760 68890 550769
rect 68834 550695 68890 550704
rect 68742 544504 68798 544513
rect 68742 544439 68798 544448
rect 68572 489886 68692 489914
rect 67640 489864 67692 489870
rect 67638 489832 67640 489841
rect 67692 489832 67694 489841
rect 67638 489767 67694 489776
rect 67638 487248 67694 487257
rect 67638 487183 67640 487192
rect 67692 487183 67694 487192
rect 67640 487154 67692 487160
rect 67638 486568 67694 486577
rect 67638 486503 67694 486512
rect 67652 486470 67680 486503
rect 67640 486464 67692 486470
rect 67640 486406 67692 486412
rect 67638 485888 67694 485897
rect 67638 485823 67640 485832
rect 67692 485823 67694 485832
rect 67640 485794 67692 485800
rect 67638 485208 67694 485217
rect 67638 485143 67694 485152
rect 67652 484498 67680 485143
rect 67640 484492 67692 484498
rect 67640 484434 67692 484440
rect 67638 483984 67694 483993
rect 67638 483919 67694 483928
rect 67652 483682 67680 483919
rect 67640 483676 67692 483682
rect 67640 483618 67692 483624
rect 67640 482996 67692 483002
rect 67640 482938 67692 482944
rect 67652 482633 67680 482938
rect 67638 482624 67694 482633
rect 67638 482559 67694 482568
rect 68008 481636 68060 481642
rect 68008 481578 68060 481584
rect 67640 481568 67692 481574
rect 67640 481510 67692 481516
rect 67652 481273 67680 481510
rect 67638 481264 67694 481273
rect 67638 481199 67694 481208
rect 68020 481137 68048 481578
rect 68006 481128 68062 481137
rect 68006 481063 68062 481072
rect 67640 480208 67692 480214
rect 67638 480176 67640 480185
rect 67692 480176 67694 480185
rect 67638 480111 67694 480120
rect 67546 478544 67602 478553
rect 67546 478479 67602 478488
rect 67560 477737 67588 478479
rect 67546 477728 67602 477737
rect 67546 477663 67602 477672
rect 67732 477488 67784 477494
rect 67732 477430 67784 477436
rect 67638 476368 67694 476377
rect 67638 476303 67694 476312
rect 67652 476134 67680 476303
rect 67744 476241 67772 477430
rect 68572 477057 68600 489886
rect 68650 484664 68706 484673
rect 68650 484599 68652 484608
rect 68704 484599 68706 484608
rect 68652 484570 68704 484576
rect 68374 477048 68430 477057
rect 68374 476983 68430 476992
rect 68558 477048 68614 477057
rect 68558 476983 68614 476992
rect 67730 476232 67786 476241
rect 67730 476167 67786 476176
rect 67640 476128 67692 476134
rect 67640 476070 67692 476076
rect 67638 475688 67694 475697
rect 67638 475623 67694 475632
rect 67652 475386 67680 475623
rect 67640 475380 67692 475386
rect 67640 475322 67692 475328
rect 67638 475008 67694 475017
rect 67638 474943 67694 474952
rect 67652 474774 67680 474943
rect 67640 474768 67692 474774
rect 67640 474710 67692 474716
rect 67454 474328 67510 474337
rect 67454 474263 67510 474272
rect 67468 473385 67496 474263
rect 67454 473376 67510 473385
rect 67454 473311 67510 473320
rect 67640 473340 67692 473346
rect 67640 473282 67692 473288
rect 67652 472705 67680 473282
rect 67638 472696 67694 472705
rect 67638 472631 67694 472640
rect 67640 471640 67692 471646
rect 67638 471608 67640 471617
rect 67692 471608 67694 471617
rect 67638 471543 67694 471552
rect 67640 471300 67692 471306
rect 67640 471242 67692 471248
rect 67652 471073 67680 471242
rect 67638 471064 67694 471073
rect 67638 470999 67694 471008
rect 67638 469704 67694 469713
rect 67638 469639 67694 469648
rect 67652 469266 67680 469639
rect 67730 469568 67786 469577
rect 67730 469503 67732 469512
rect 67784 469503 67786 469512
rect 67732 469474 67784 469480
rect 67640 469260 67692 469266
rect 67640 469202 67692 469208
rect 67730 468344 67786 468353
rect 67730 468279 67786 468288
rect 67640 468240 67692 468246
rect 67638 468208 67640 468217
rect 67692 468208 67694 468217
rect 67638 468143 67694 468152
rect 67744 467906 67772 468279
rect 67732 467900 67784 467906
rect 67732 467842 67784 467848
rect 67638 466848 67694 466857
rect 67638 466783 67640 466792
rect 67692 466783 67694 466792
rect 67640 466754 67692 466760
rect 67376 466426 67588 466454
rect 67560 465610 67588 466426
rect 67730 466168 67786 466177
rect 67730 466103 67786 466112
rect 67638 465624 67694 465633
rect 67560 465582 67638 465610
rect 67560 460934 67588 465582
rect 67638 465559 67694 465568
rect 67744 465118 67772 466103
rect 67732 465112 67784 465118
rect 67732 465054 67784 465060
rect 67822 464128 67878 464137
rect 67822 464063 67878 464072
rect 67640 463820 67692 463826
rect 67640 463762 67692 463768
rect 67652 463729 67680 463762
rect 67836 463758 67864 464063
rect 67824 463752 67876 463758
rect 67638 463720 67694 463729
rect 67824 463694 67876 463700
rect 67638 463655 67694 463664
rect 67732 463684 67784 463690
rect 67732 463626 67784 463632
rect 67638 463448 67694 463457
rect 67638 463383 67694 463392
rect 67652 462398 67680 463383
rect 67744 462913 67772 463626
rect 67730 462904 67786 462913
rect 67730 462839 67786 462848
rect 67640 462392 67692 462398
rect 67640 462334 67692 462340
rect 67638 461408 67694 461417
rect 67638 461343 67694 461352
rect 67652 460970 67680 461343
rect 67376 460906 67588 460934
rect 67640 460964 67692 460970
rect 67640 460906 67692 460912
rect 67272 439612 67324 439618
rect 67272 439554 67324 439560
rect 67376 397526 67404 460906
rect 67638 460728 67694 460737
rect 67638 460663 67694 460672
rect 67652 460290 67680 460663
rect 67640 460284 67692 460290
rect 67640 460226 67692 460232
rect 67732 460216 67784 460222
rect 67730 460184 67732 460193
rect 67784 460184 67786 460193
rect 67730 460119 67786 460128
rect 67456 458856 67508 458862
rect 67640 458856 67692 458862
rect 67456 458798 67508 458804
rect 67638 458824 67640 458833
rect 67692 458824 67694 458833
rect 67364 397520 67416 397526
rect 67364 397462 67416 397468
rect 67376 369753 67404 397462
rect 67362 369744 67418 369753
rect 67362 369679 67418 369688
rect 67468 362409 67496 458798
rect 67638 458759 67694 458768
rect 67638 458688 67694 458697
rect 67638 458623 67694 458632
rect 67652 458318 67680 458623
rect 67640 458312 67692 458318
rect 67640 458254 67692 458260
rect 67732 458176 67784 458182
rect 67732 458118 67784 458124
rect 67638 458008 67694 458017
rect 67638 457943 67694 457952
rect 67652 457502 67680 457943
rect 67640 457496 67692 457502
rect 67744 457473 67772 458118
rect 67640 457438 67692 457444
rect 67730 457464 67786 457473
rect 67730 457399 67786 457408
rect 67640 456068 67692 456074
rect 67640 456010 67692 456016
rect 67652 455977 67680 456010
rect 67638 455968 67694 455977
rect 67638 455903 67694 455912
rect 67640 455388 67692 455394
rect 67640 455330 67692 455336
rect 67652 455297 67680 455330
rect 67638 455288 67694 455297
rect 67638 455223 67694 455232
rect 67640 454028 67692 454034
rect 67640 453970 67692 453976
rect 67652 453937 67680 453970
rect 67638 453928 67694 453937
rect 67638 453863 67694 453872
rect 67640 453348 67692 453354
rect 67640 453290 67692 453296
rect 67652 453257 67680 453290
rect 67638 453248 67694 453257
rect 67638 453183 67694 453192
rect 67638 449984 67694 449993
rect 67638 449919 67640 449928
rect 67692 449919 67694 449928
rect 67640 449890 67692 449896
rect 67730 449304 67786 449313
rect 67730 449239 67786 449248
rect 67640 449200 67692 449206
rect 67638 449168 67640 449177
rect 67692 449168 67694 449177
rect 67638 449103 67694 449112
rect 67744 448633 67772 449239
rect 67730 448624 67786 448633
rect 67730 448559 67786 448568
rect 67730 447808 67786 447817
rect 67730 447743 67786 447752
rect 67638 447264 67694 447273
rect 67638 447199 67640 447208
rect 67692 447199 67694 447208
rect 67640 447170 67692 447176
rect 67744 447166 67772 447743
rect 67732 447160 67784 447166
rect 67732 447102 67784 447108
rect 67730 446584 67786 446593
rect 67730 446519 67786 446528
rect 67638 446448 67694 446457
rect 67638 446383 67640 446392
rect 67692 446383 67694 446392
rect 67640 446354 67692 446360
rect 67744 445806 67772 446519
rect 67732 445800 67784 445806
rect 67732 445742 67784 445748
rect 68190 445496 68246 445505
rect 68190 445431 68246 445440
rect 67638 443728 67694 443737
rect 67638 443663 67640 443672
rect 67692 443663 67694 443672
rect 67640 443634 67692 443640
rect 67640 442944 67692 442950
rect 67640 442886 67692 442892
rect 67652 442513 67680 442886
rect 67638 442504 67694 442513
rect 67638 442439 67694 442448
rect 67638 442368 67694 442377
rect 67638 442303 67694 442312
rect 67652 442270 67680 442303
rect 67640 442264 67692 442270
rect 67640 442206 67692 442212
rect 67640 441584 67692 441590
rect 67640 441526 67692 441532
rect 67652 441153 67680 441526
rect 67638 441144 67694 441153
rect 67694 441102 67772 441130
rect 67638 441079 67694 441088
rect 67640 441040 67692 441046
rect 67638 441008 67640 441017
rect 67692 441008 67694 441017
rect 67638 440943 67694 440952
rect 67744 440314 67772 441102
rect 67560 440286 67772 440314
rect 67454 362400 67510 362409
rect 67454 362335 67510 362344
rect 67364 353320 67416 353326
rect 67364 353262 67416 353268
rect 66260 349172 66312 349178
rect 66260 349114 66312 349120
rect 67272 342304 67324 342310
rect 67272 342246 67324 342252
rect 66074 331800 66130 331809
rect 66074 331735 66130 331744
rect 65984 326392 66036 326398
rect 65984 326334 66036 326340
rect 67284 320958 67312 342246
rect 67376 330546 67404 353262
rect 67364 330540 67416 330546
rect 67364 330482 67416 330488
rect 67468 323746 67496 362335
rect 67560 341601 67588 440286
rect 67638 382528 67694 382537
rect 67638 382463 67694 382472
rect 67652 382294 67680 382463
rect 67640 382288 67692 382294
rect 67640 382230 67692 382236
rect 67640 380860 67692 380866
rect 67640 380802 67692 380808
rect 67652 380769 67680 380802
rect 67638 380760 67694 380769
rect 67638 380695 67694 380704
rect 67638 379808 67694 379817
rect 67638 379743 67694 379752
rect 67652 379574 67680 379743
rect 67640 379568 67692 379574
rect 67640 379510 67692 379516
rect 67640 377460 67692 377466
rect 67640 377402 67692 377408
rect 67652 377369 67680 377402
rect 67638 377360 67694 377369
rect 67638 377295 67694 377304
rect 67640 374672 67692 374678
rect 67640 374614 67692 374620
rect 67652 374513 67680 374614
rect 67638 374504 67694 374513
rect 67638 374439 67694 374448
rect 67640 372564 67692 372570
rect 67640 372506 67692 372512
rect 67652 371793 67680 372506
rect 67732 371952 67784 371958
rect 67730 371920 67732 371929
rect 67784 371920 67786 371929
rect 67730 371855 67786 371864
rect 67638 371784 67694 371793
rect 67638 371719 67694 371728
rect 67640 369844 67692 369850
rect 67640 369786 67692 369792
rect 67652 369073 67680 369786
rect 67638 369064 67694 369073
rect 67638 368999 67694 369008
rect 68008 367056 68060 367062
rect 68008 366998 68060 367004
rect 67638 366480 67694 366489
rect 67638 366415 67694 366424
rect 67652 366382 67680 366415
rect 67640 366376 67692 366382
rect 67640 366318 67692 366324
rect 68020 366081 68048 366998
rect 68006 366072 68062 366081
rect 68006 366007 68062 366016
rect 67638 364440 67694 364449
rect 67638 364375 67640 364384
rect 67692 364375 67694 364384
rect 67640 364346 67692 364352
rect 67732 364336 67784 364342
rect 67730 364304 67732 364313
rect 67784 364304 67786 364313
rect 67730 364239 67786 364248
rect 67640 363656 67692 363662
rect 67638 363624 67640 363633
rect 67692 363624 67694 363633
rect 67638 363559 67694 363568
rect 67640 361548 67692 361554
rect 67640 361490 67692 361496
rect 67652 360913 67680 361490
rect 67638 360904 67694 360913
rect 67638 360839 67694 360848
rect 67638 359272 67694 359281
rect 67638 359207 67694 359216
rect 67652 358834 67680 359207
rect 67640 358828 67692 358834
rect 67640 358770 67692 358776
rect 67730 358184 67786 358193
rect 67730 358119 67786 358128
rect 67640 358080 67692 358086
rect 67638 358048 67640 358057
rect 67692 358048 67694 358057
rect 67638 357983 67694 357992
rect 67744 357474 67772 358119
rect 67732 357468 67784 357474
rect 67732 357410 67784 357416
rect 67640 356040 67692 356046
rect 67640 355982 67692 355988
rect 67652 355881 67680 355982
rect 67732 355972 67784 355978
rect 67732 355914 67784 355920
rect 67638 355872 67694 355881
rect 67638 355807 67694 355816
rect 67744 355473 67772 355914
rect 67730 355464 67786 355473
rect 67730 355399 67786 355408
rect 67638 353832 67694 353841
rect 67638 353767 67694 353776
rect 67652 353326 67680 353767
rect 67640 353320 67692 353326
rect 67640 353262 67692 353268
rect 67640 352640 67692 352646
rect 67638 352608 67640 352617
rect 67692 352608 67694 352617
rect 67638 352543 67694 352552
rect 67914 351248 67970 351257
rect 67914 351183 67916 351192
rect 67968 351183 67970 351192
rect 67916 351154 67968 351160
rect 67640 350532 67692 350538
rect 67640 350474 67692 350480
rect 67652 350441 67680 350474
rect 67638 350432 67694 350441
rect 67638 350367 67694 350376
rect 67640 349104 67692 349110
rect 67638 349072 67640 349081
rect 67692 349072 67694 349081
rect 67638 349007 67694 349016
rect 67732 347744 67784 347750
rect 67732 347686 67784 347692
rect 67638 347168 67694 347177
rect 67638 347103 67694 347112
rect 67652 347070 67680 347103
rect 67640 347064 67692 347070
rect 67744 347041 67772 347686
rect 67640 347006 67692 347012
rect 67730 347032 67786 347041
rect 67730 346967 67786 346976
rect 68204 346390 68232 445431
rect 68282 444272 68338 444281
rect 68282 444207 68338 444216
rect 68296 364334 68324 444207
rect 68388 402974 68416 476983
rect 68756 460934 68784 544439
rect 68572 460906 68784 460934
rect 68572 445505 68600 460906
rect 68848 454594 68876 550695
rect 68926 543960 68982 543969
rect 68926 543895 68982 543904
rect 68756 454566 68876 454594
rect 68756 451353 68784 454566
rect 68742 451344 68798 451353
rect 68742 451279 68798 451288
rect 68558 445496 68614 445505
rect 68558 445431 68614 445440
rect 68756 441614 68784 451279
rect 68940 444281 68968 543895
rect 69032 543289 69060 696934
rect 70952 584044 71004 584050
rect 70952 583986 71004 583992
rect 70400 583976 70452 583982
rect 70400 583918 70452 583924
rect 70308 583772 70360 583778
rect 70308 583714 70360 583720
rect 69202 582448 69258 582457
rect 69202 582383 69258 582392
rect 69112 577040 69164 577046
rect 69112 576982 69164 576988
rect 69018 543280 69074 543289
rect 69018 543215 69074 543224
rect 69124 482905 69152 576982
rect 69216 545329 69244 582383
rect 69768 581318 70058 581346
rect 69768 577046 69796 581318
rect 69756 577040 69808 577046
rect 69756 576982 69808 576988
rect 69202 545320 69258 545329
rect 69202 545255 69258 545264
rect 69202 541784 69258 541793
rect 69202 541719 69258 541728
rect 69216 525774 69244 541719
rect 69664 541680 69716 541686
rect 69664 541622 69716 541628
rect 69296 533384 69348 533390
rect 69296 533326 69348 533332
rect 69204 525768 69256 525774
rect 69202 525736 69204 525745
rect 69256 525736 69258 525745
rect 69202 525671 69258 525680
rect 69110 482896 69166 482905
rect 69110 482831 69166 482840
rect 68926 444272 68982 444281
rect 68926 444207 68982 444216
rect 68756 441586 68876 441614
rect 68388 402946 68784 402974
rect 68756 383722 68784 402946
rect 68744 383716 68796 383722
rect 68744 383658 68796 383664
rect 68756 383489 68784 383658
rect 68742 383480 68798 383489
rect 68742 383415 68798 383424
rect 68376 370184 68428 370190
rect 68374 370152 68376 370161
rect 68428 370152 68430 370161
rect 68374 370087 68430 370096
rect 68848 364334 68876 441586
rect 69124 437617 69152 482831
rect 69308 460934 69336 533326
rect 69676 498846 69704 541622
rect 69768 540110 70058 540138
rect 69768 533390 69796 540110
rect 70320 539102 70348 583714
rect 70412 581890 70440 583918
rect 70964 581890 70992 583986
rect 71056 582010 71084 700334
rect 71792 583030 71820 702986
rect 75184 702840 75236 702846
rect 75184 702782 75236 702788
rect 71872 594856 71924 594862
rect 71872 594798 71924 594804
rect 71780 583024 71832 583030
rect 71780 582966 71832 582972
rect 71884 582162 71912 594798
rect 74632 590708 74684 590714
rect 74632 590650 74684 590656
rect 73344 583908 73396 583914
rect 73344 583850 73396 583856
rect 71792 582134 71912 582162
rect 71044 582004 71096 582010
rect 71044 581946 71096 581952
rect 70412 581862 70702 581890
rect 70964 581862 71300 581890
rect 71792 581754 71820 582134
rect 73356 581890 73384 583850
rect 74644 581890 74672 590650
rect 75196 586514 75224 702782
rect 75104 586486 75224 586514
rect 75104 583953 75132 586486
rect 76576 585274 76604 702986
rect 77956 596174 77984 703258
rect 79324 702636 79376 702642
rect 79324 702578 79376 702584
rect 79336 596174 79364 702578
rect 89180 702434 89208 703520
rect 95148 703248 95200 703254
rect 95148 703190 95200 703196
rect 88352 702406 89208 702434
rect 85580 597576 85632 597582
rect 85580 597518 85632 597524
rect 77956 596146 78076 596174
rect 76564 585268 76616 585274
rect 76564 585210 76616 585216
rect 75090 583944 75146 583953
rect 73278 581862 73384 581890
rect 74566 581862 74672 581890
rect 75012 583902 75090 583930
rect 75012 581754 75040 583902
rect 75090 583879 75146 583888
rect 76576 581890 76604 585210
rect 78048 585206 78076 596146
rect 79244 596146 79364 596174
rect 85592 596174 85620 597518
rect 85592 596146 85712 596174
rect 78036 585200 78088 585206
rect 78036 585142 78088 585148
rect 77852 584112 77904 584118
rect 77852 584054 77904 584060
rect 76748 582548 76800 582554
rect 76748 582490 76800 582496
rect 76498 581862 76604 581890
rect 76760 581890 76788 582490
rect 77864 581890 77892 584054
rect 76760 581862 77096 581890
rect 77786 581862 77892 581890
rect 78048 581890 78076 585142
rect 79244 584118 79272 596146
rect 82084 591320 82136 591326
rect 82084 591262 82136 591268
rect 79324 586628 79376 586634
rect 79324 586570 79376 586576
rect 79232 584112 79284 584118
rect 79232 584054 79284 584060
rect 79336 581890 79364 586570
rect 80612 585336 80664 585342
rect 80612 585278 80664 585284
rect 80624 581890 80652 585278
rect 82096 583817 82124 591262
rect 85304 586696 85356 586702
rect 85304 586638 85356 586644
rect 84292 586560 84344 586566
rect 84292 586502 84344 586508
rect 82542 583944 82598 583953
rect 82542 583879 82598 583888
rect 81438 583808 81494 583817
rect 81438 583743 81494 583752
rect 82082 583808 82138 583817
rect 82082 583743 82138 583752
rect 81452 581890 81480 583743
rect 82556 581890 82584 583879
rect 83372 583772 83424 583778
rect 83372 583714 83424 583720
rect 83280 582616 83332 582622
rect 83280 582558 83332 582564
rect 83292 581890 83320 582558
rect 78048 581862 78384 581890
rect 79336 581862 79672 581890
rect 80624 581862 80960 581890
rect 81452 581862 81604 581890
rect 82294 581862 82584 581890
rect 82938 581862 83320 581890
rect 83384 581890 83412 583714
rect 84304 581890 84332 586502
rect 84476 582480 84528 582486
rect 84476 582422 84528 582428
rect 83384 581862 83536 581890
rect 84226 581862 84332 581890
rect 84488 581890 84516 582422
rect 84488 581862 84824 581890
rect 75460 581800 75512 581806
rect 71792 581726 71944 581754
rect 72252 581738 72588 581754
rect 72240 581732 72588 581738
rect 72292 581726 72588 581732
rect 75012 581726 75164 581754
rect 85316 581754 85344 586638
rect 85684 581890 85712 596146
rect 88352 588606 88380 702406
rect 90364 670744 90416 670750
rect 90364 670686 90416 670692
rect 90376 591326 90404 670686
rect 93124 618316 93176 618322
rect 93124 618258 93176 618264
rect 90364 591320 90416 591326
rect 90364 591262 90416 591268
rect 87328 588600 87380 588606
rect 87328 588542 87380 588548
rect 88340 588600 88392 588606
rect 88340 588542 88392 588548
rect 87340 585274 87368 588542
rect 91008 586628 91060 586634
rect 91008 586570 91060 586576
rect 87328 585268 87380 585274
rect 87328 585210 87380 585216
rect 87512 585268 87564 585274
rect 87512 585210 87564 585216
rect 87524 581890 87552 585210
rect 88248 584248 88300 584254
rect 88248 584190 88300 584196
rect 88260 581890 88288 584190
rect 88984 583772 89036 583778
rect 88984 583714 89036 583720
rect 88996 581890 89024 583714
rect 89628 582480 89680 582486
rect 89628 582422 89680 582428
rect 89640 581890 89668 582422
rect 91020 581890 91048 586570
rect 91650 586392 91706 586401
rect 91650 586327 91706 586336
rect 91560 582548 91612 582554
rect 91560 582490 91612 582496
rect 91572 581890 91600 582490
rect 85684 581862 86112 581890
rect 87446 581862 87552 581890
rect 88090 581862 88288 581890
rect 88734 581862 89024 581890
rect 89378 581862 89668 581890
rect 90666 581862 91048 581890
rect 91310 581862 91600 581890
rect 91664 581890 91692 586327
rect 93136 585410 93164 618258
rect 94872 586560 94924 586566
rect 94872 586502 94924 586508
rect 94134 586392 94190 586401
rect 94134 586327 94190 586336
rect 93124 585404 93176 585410
rect 93124 585346 93176 585352
rect 92848 582684 92900 582690
rect 92848 582626 92900 582632
rect 92860 581890 92888 582626
rect 94148 581890 94176 586327
rect 94884 581890 94912 586502
rect 95160 585342 95188 703190
rect 104808 702976 104860 702982
rect 104808 702918 104860 702924
rect 104820 586770 104848 702918
rect 105464 702434 105492 703520
rect 109684 703180 109736 703186
rect 109684 703122 109736 703128
rect 108948 702568 109000 702574
rect 108948 702510 109000 702516
rect 105464 702406 105584 702434
rect 103520 586764 103572 586770
rect 103520 586706 103572 586712
rect 104808 586764 104860 586770
rect 104808 586706 104860 586712
rect 95884 585404 95936 585410
rect 95884 585346 95936 585352
rect 95148 585336 95200 585342
rect 95148 585278 95200 585284
rect 95160 582162 95188 585278
rect 91664 581862 91908 581890
rect 92598 581862 92888 581890
rect 93886 581862 94176 581890
rect 94530 581862 94912 581890
rect 94976 582134 95188 582162
rect 94976 581754 95004 582134
rect 95896 581890 95924 585346
rect 97908 585200 97960 585206
rect 97908 585142 97960 585148
rect 96528 584044 96580 584050
rect 96528 583986 96580 583992
rect 96540 581890 96568 583986
rect 96712 583840 96764 583846
rect 96712 583782 96764 583788
rect 95818 581862 95924 581890
rect 96462 581862 96568 581890
rect 96724 581890 96752 583782
rect 97920 581890 97948 585142
rect 103532 585018 103560 586706
rect 103348 584990 103560 585018
rect 101402 584352 101458 584361
rect 101402 584287 101458 584296
rect 101416 584186 101444 584287
rect 98736 584180 98788 584186
rect 98736 584122 98788 584128
rect 101404 584180 101456 584186
rect 101404 584122 101456 584128
rect 98748 581890 98776 584122
rect 99288 584112 99340 584118
rect 99288 584054 99340 584060
rect 99300 581890 99328 584054
rect 101312 583976 101364 583982
rect 101312 583918 101364 583924
rect 101324 581890 101352 583918
rect 101864 583908 101916 583914
rect 101864 583850 101916 583856
rect 101876 581890 101904 583850
rect 102140 583772 102192 583778
rect 102140 583714 102192 583720
rect 102152 583030 102180 583714
rect 102140 583024 102192 583030
rect 102140 582966 102192 582972
rect 103348 581890 103376 584990
rect 104440 583840 104492 583846
rect 103886 583808 103942 583817
rect 104440 583782 104492 583788
rect 103886 583743 103942 583752
rect 103900 581890 103928 583743
rect 104452 581890 104480 583782
rect 105268 583772 105320 583778
rect 105268 583714 105320 583720
rect 96724 581862 97060 581890
rect 97750 581862 97948 581890
rect 98394 581862 98776 581890
rect 99038 581862 99328 581890
rect 100970 581862 101352 581890
rect 101614 581862 101904 581890
rect 102902 581862 103376 581890
rect 103546 581862 103928 581890
rect 104190 581862 104480 581890
rect 102598 581768 102654 581777
rect 75512 581748 75808 581754
rect 75460 581742 75808 581748
rect 75472 581726 75808 581742
rect 78692 581738 79028 581754
rect 78680 581732 79028 581738
rect 72240 581674 72292 581680
rect 78732 581726 79028 581732
rect 85316 581726 85468 581754
rect 90022 581738 90312 581754
rect 90022 581732 90324 581738
rect 90022 581726 90272 581732
rect 78680 581674 78732 581680
rect 94976 581726 95128 581754
rect 100326 581738 100616 581754
rect 100326 581732 100628 581738
rect 100326 581726 100576 581732
rect 90272 581674 90324 581680
rect 102258 581726 102598 581754
rect 105280 581754 105308 583714
rect 104834 581738 105032 581754
rect 104834 581732 105044 581738
rect 104834 581726 104992 581732
rect 102598 581703 102654 581712
rect 100576 581674 100628 581680
rect 105280 581726 105478 581754
rect 104992 581674 105044 581680
rect 105556 572914 105584 702406
rect 106280 698964 106332 698970
rect 106280 698906 106332 698912
rect 105636 584248 105688 584254
rect 105636 584190 105688 584196
rect 105648 576162 105676 584190
rect 106186 577824 106242 577833
rect 106186 577759 106242 577768
rect 105636 576156 105688 576162
rect 105636 576098 105688 576104
rect 105556 572886 105676 572914
rect 105648 572830 105676 572886
rect 105636 572824 105688 572830
rect 105636 572766 105688 572772
rect 105726 548448 105782 548457
rect 105726 548383 105782 548392
rect 70412 540110 70702 540138
rect 70308 539096 70360 539102
rect 70308 539038 70360 539044
rect 69756 533384 69808 533390
rect 69756 533326 69808 533332
rect 70412 529310 70440 540110
rect 71332 536110 71360 540138
rect 71976 539186 72004 540138
rect 71884 539158 72004 539186
rect 71320 536104 71372 536110
rect 71320 536046 71372 536052
rect 71884 532030 71912 539158
rect 71964 539096 72016 539102
rect 71964 539038 72016 539044
rect 71872 532024 71924 532030
rect 71872 531966 71924 531972
rect 70400 529304 70452 529310
rect 70400 529246 70452 529252
rect 71976 499574 72004 539038
rect 72424 533316 72476 533322
rect 72424 533258 72476 533264
rect 71792 499546 72004 499574
rect 69664 498840 69716 498846
rect 69664 498782 69716 498788
rect 71688 493332 71740 493338
rect 71688 493274 71740 493280
rect 70952 492720 71004 492726
rect 70952 492662 71004 492668
rect 70400 492176 70452 492182
rect 70400 492118 70452 492124
rect 70032 492108 70084 492114
rect 70032 492050 70084 492056
rect 70044 489940 70072 492050
rect 70412 489954 70440 492118
rect 70964 489954 70992 492662
rect 71700 491314 71728 493274
rect 71792 491881 71820 499546
rect 72436 492658 72464 533258
rect 72620 532234 72648 540138
rect 73264 534750 73292 540138
rect 73908 538218 73936 540138
rect 73896 538212 73948 538218
rect 73896 538154 73948 538160
rect 73252 534744 73304 534750
rect 73252 534686 73304 534692
rect 72608 532228 72660 532234
rect 72608 532170 72660 532176
rect 74552 529145 74580 540138
rect 75196 538214 75224 540138
rect 76467 540110 76512 540138
rect 75104 538186 75224 538214
rect 75104 532098 75132 538186
rect 75184 535016 75236 535022
rect 75184 534958 75236 534964
rect 75092 532092 75144 532098
rect 75092 532034 75144 532040
rect 74538 529136 74594 529145
rect 74538 529071 74594 529080
rect 74540 498840 74592 498846
rect 74540 498782 74592 498788
rect 72424 492652 72476 492658
rect 72424 492594 72476 492600
rect 72240 492040 72292 492046
rect 72240 491982 72292 491988
rect 71778 491872 71834 491881
rect 71778 491807 71834 491816
rect 71792 491502 71820 491807
rect 71780 491496 71832 491502
rect 71780 491438 71832 491444
rect 71700 491286 71820 491314
rect 71792 489954 71820 491286
rect 72252 489954 72280 491982
rect 73252 490612 73304 490618
rect 73252 490554 73304 490560
rect 70412 489926 70656 489954
rect 70964 489926 71300 489954
rect 71792 489926 71944 489954
rect 72252 489926 72588 489954
rect 73264 489940 73292 490554
rect 74552 489940 74580 498782
rect 75196 495038 75224 534958
rect 76484 532166 76512 540110
rect 76472 532160 76524 532166
rect 76472 532102 76524 532108
rect 77128 529242 77156 540138
rect 77772 534818 77800 540138
rect 78416 534954 78444 540138
rect 78404 534948 78456 534954
rect 78404 534890 78456 534896
rect 77760 534812 77812 534818
rect 77760 534754 77812 534760
rect 77116 529236 77168 529242
rect 77116 529178 77168 529184
rect 78404 495508 78456 495514
rect 78404 495450 78456 495456
rect 78416 495038 78444 495450
rect 75184 495032 75236 495038
rect 75184 494974 75236 494980
rect 78404 495032 78456 495038
rect 78404 494974 78456 494980
rect 74816 493400 74868 493406
rect 74816 493342 74868 493348
rect 74828 489954 74856 493342
rect 75828 493060 75880 493066
rect 75828 493002 75880 493008
rect 74828 489926 75164 489954
rect 75840 489940 75868 493002
rect 77760 492720 77812 492726
rect 77760 492662 77812 492668
rect 76472 492040 76524 492046
rect 76472 491982 76524 491988
rect 76484 489940 76512 491982
rect 76748 491496 76800 491502
rect 76748 491438 76800 491444
rect 76760 489954 76788 491438
rect 76760 489926 77096 489954
rect 77772 489940 77800 492662
rect 78416 489940 78444 494974
rect 79060 490686 79088 540138
rect 79704 537674 79732 540138
rect 80348 538218 80376 540138
rect 80336 538212 80388 538218
rect 80336 538154 80388 538160
rect 79692 537668 79744 537674
rect 79692 537610 79744 537616
rect 80348 537577 80376 538154
rect 80334 537568 80390 537577
rect 80334 537503 80390 537512
rect 80610 499624 80666 499633
rect 80610 499559 80666 499568
rect 80624 498846 80652 499559
rect 80612 498840 80664 498846
rect 80612 498782 80664 498788
rect 79692 496188 79744 496194
rect 79692 496130 79744 496136
rect 79048 490680 79100 490686
rect 79048 490622 79100 490628
rect 79704 489940 79732 496130
rect 80992 496126 81020 540138
rect 81636 537441 81664 540138
rect 82907 540110 82952 540138
rect 82924 537742 82952 540110
rect 82912 537736 82964 537742
rect 82912 537678 82964 537684
rect 81622 537432 81678 537441
rect 81622 537367 81678 537376
rect 83464 536852 83516 536858
rect 83464 536794 83516 536800
rect 83280 497480 83332 497486
rect 83280 497422 83332 497428
rect 81532 496256 81584 496262
rect 81532 496198 81584 496204
rect 80980 496120 81032 496126
rect 80980 496062 81032 496068
rect 80980 494828 81032 494834
rect 80980 494770 81032 494776
rect 80060 491360 80112 491366
rect 80060 491302 80112 491308
rect 80072 489954 80100 491302
rect 80072 489926 80316 489954
rect 80992 489940 81020 494770
rect 81544 493066 81572 496198
rect 83292 495446 83320 497422
rect 83476 496330 83504 536794
rect 83568 534886 83596 540138
rect 84108 537668 84160 537674
rect 84108 537610 84160 537616
rect 83556 534880 83608 534886
rect 83556 534822 83608 534828
rect 84120 497554 84148 537610
rect 84108 497548 84160 497554
rect 84108 497490 84160 497496
rect 83464 496324 83516 496330
rect 83464 496266 83516 496272
rect 83280 495440 83332 495446
rect 83280 495382 83332 495388
rect 82912 494760 82964 494766
rect 82912 494702 82964 494708
rect 81532 493060 81584 493066
rect 81532 493002 81584 493008
rect 81624 492856 81676 492862
rect 81624 492798 81676 492804
rect 81636 489940 81664 492798
rect 82266 491600 82322 491609
rect 82266 491535 82322 491544
rect 82280 489940 82308 491535
rect 82924 489940 82952 494702
rect 83292 489954 83320 495382
rect 84212 494737 84240 540138
rect 84856 532098 84884 540138
rect 85500 536858 85528 540138
rect 86144 537606 86172 540138
rect 86132 537600 86184 537606
rect 86132 537542 86184 537548
rect 85488 536852 85540 536858
rect 85488 536794 85540 536800
rect 84844 532092 84896 532098
rect 84844 532034 84896 532040
rect 86788 499574 86816 540138
rect 87142 536072 87198 536081
rect 87142 536007 87198 536016
rect 86788 499546 86908 499574
rect 85580 497616 85632 497622
rect 85580 497558 85632 497564
rect 85592 495394 85620 497558
rect 85500 495366 85620 495394
rect 84198 494728 84254 494737
rect 84198 494663 84254 494672
rect 84844 492652 84896 492658
rect 84844 492594 84896 492600
rect 83292 489926 83536 489954
rect 84856 489940 84884 492594
rect 85500 489940 85528 495366
rect 86132 492108 86184 492114
rect 86132 492050 86184 492056
rect 86144 489940 86172 492050
rect 86776 491496 86828 491502
rect 86776 491438 86828 491444
rect 86788 489940 86816 491438
rect 86880 490618 86908 499546
rect 87156 492114 87184 536007
rect 87432 500177 87460 540138
rect 88076 538121 88104 540138
rect 89347 540110 89392 540138
rect 88062 538112 88118 538121
rect 88062 538047 88118 538056
rect 87418 500168 87474 500177
rect 87418 500103 87474 500112
rect 87420 499520 87472 499526
rect 87420 499462 87472 499468
rect 87144 492108 87196 492114
rect 87144 492050 87196 492056
rect 86868 490612 86920 490618
rect 86868 490554 86920 490560
rect 87432 489940 87460 499462
rect 89364 498914 89392 540110
rect 90008 537674 90036 540138
rect 89996 537668 90048 537674
rect 89996 537610 90048 537616
rect 89352 498908 89404 498914
rect 89352 498850 89404 498856
rect 88064 498840 88116 498846
rect 88064 498782 88116 498788
rect 88076 489940 88104 498782
rect 90272 493468 90324 493474
rect 90272 493410 90324 493416
rect 88708 493400 88760 493406
rect 88708 493342 88760 493348
rect 88720 489940 88748 493342
rect 90284 492794 90312 493410
rect 90272 492788 90324 492794
rect 90272 492730 90324 492736
rect 89904 492108 89956 492114
rect 89904 492050 89956 492056
rect 89916 490754 89944 492050
rect 89996 491836 90048 491842
rect 89996 491778 90048 491784
rect 89904 490748 89956 490754
rect 89904 490690 89956 490696
rect 90008 489940 90036 491778
rect 90284 489954 90312 492730
rect 90652 491978 90680 540138
rect 91296 537538 91324 540138
rect 91284 537532 91336 537538
rect 91284 537474 91336 537480
rect 91008 534812 91060 534818
rect 91008 534754 91060 534760
rect 90640 491972 90692 491978
rect 90640 491914 90692 491920
rect 91020 491842 91048 534754
rect 91940 499574 91968 540138
rect 92584 534721 92612 540138
rect 92570 534712 92626 534721
rect 92570 534647 92626 534656
rect 91940 499546 92060 499574
rect 91100 497684 91152 497690
rect 91100 497626 91152 497632
rect 91008 491836 91060 491842
rect 91008 491778 91060 491784
rect 91020 491570 91048 491778
rect 91008 491564 91060 491570
rect 91008 491506 91060 491512
rect 90284 489926 90620 489954
rect 91112 489818 91140 497626
rect 91928 493876 91980 493882
rect 91928 493818 91980 493824
rect 91940 489940 91968 493818
rect 92032 492114 92060 499546
rect 93228 497690 93256 540138
rect 93872 534750 93900 540138
rect 94516 536858 94544 540138
rect 95787 540110 95832 540138
rect 95148 539028 95200 539034
rect 95148 538970 95200 538976
rect 94504 536852 94556 536858
rect 94504 536794 94556 536800
rect 93860 534744 93912 534750
rect 93860 534686 93912 534692
rect 93768 532024 93820 532030
rect 93768 531966 93820 531972
rect 93216 497684 93268 497690
rect 93216 497626 93268 497632
rect 93780 494086 93808 531966
rect 95056 496120 95108 496126
rect 95056 496062 95108 496068
rect 94964 495032 95016 495038
rect 94964 494974 95016 494980
rect 94872 494896 94924 494902
rect 94872 494838 94924 494844
rect 92480 494080 92532 494086
rect 92480 494022 92532 494028
rect 93768 494080 93820 494086
rect 93768 494022 93820 494028
rect 92492 492658 92520 494022
rect 93216 493332 93268 493338
rect 93216 493274 93268 493280
rect 92480 492652 92532 492658
rect 92480 492594 92532 492600
rect 92020 492108 92072 492114
rect 92020 492050 92072 492056
rect 92572 491700 92624 491706
rect 92572 491642 92624 491648
rect 92584 489940 92612 491642
rect 93228 489940 93256 493274
rect 93860 491360 93912 491366
rect 93860 491302 93912 491308
rect 93872 489940 93900 491302
rect 94884 489954 94912 494838
rect 94976 491706 95004 494974
rect 95068 493882 95096 496062
rect 95056 493876 95108 493882
rect 95056 493818 95108 493824
rect 95160 491706 95188 538970
rect 95804 537606 95832 540110
rect 95792 537600 95844 537606
rect 95792 537542 95844 537548
rect 96448 499574 96476 540138
rect 97092 537742 97120 540138
rect 97080 537736 97132 537742
rect 97080 537678 97132 537684
rect 97736 500313 97764 540138
rect 98380 539578 98408 540138
rect 98368 539572 98420 539578
rect 98368 539514 98420 539520
rect 98380 538214 98408 539514
rect 99024 539510 99052 540138
rect 99012 539504 99064 539510
rect 99012 539446 99064 539452
rect 99024 538898 99052 539446
rect 99288 538960 99340 538966
rect 99288 538902 99340 538908
rect 99012 538892 99064 538898
rect 99012 538834 99064 538840
rect 98380 538186 98684 538214
rect 97722 500304 97778 500313
rect 97722 500239 97778 500248
rect 96264 499546 96476 499574
rect 95792 493536 95844 493542
rect 95792 493478 95844 493484
rect 94964 491700 95016 491706
rect 94964 491642 95016 491648
rect 95148 491700 95200 491706
rect 95148 491642 95200 491648
rect 94884 489926 95128 489954
rect 95804 489940 95832 493478
rect 96264 490686 96292 499546
rect 98656 494970 98684 538186
rect 98644 494964 98696 494970
rect 98644 494906 98696 494912
rect 96528 492856 96580 492862
rect 96528 492798 96580 492804
rect 96344 491700 96396 491706
rect 96344 491642 96396 491648
rect 96356 491314 96384 491642
rect 96436 491496 96488 491502
rect 96434 491464 96436 491473
rect 96488 491464 96490 491473
rect 96434 491399 96490 491408
rect 96434 491328 96490 491337
rect 96356 491286 96434 491314
rect 96540 491298 96568 492798
rect 99300 492658 99328 538902
rect 99668 528554 99696 540138
rect 100312 537538 100340 540138
rect 100956 538150 100984 540138
rect 102227 540110 102272 540138
rect 100944 538144 100996 538150
rect 100944 538086 100996 538092
rect 100300 537532 100352 537538
rect 100300 537474 100352 537480
rect 100956 537441 100984 538086
rect 102244 537742 102272 540110
rect 102140 537736 102192 537742
rect 102140 537678 102192 537684
rect 102232 537736 102284 537742
rect 102232 537678 102284 537684
rect 100942 537432 100998 537441
rect 100942 537367 100998 537376
rect 101956 536716 102008 536722
rect 101956 536658 102008 536664
rect 99746 535392 99802 535401
rect 99746 535327 99802 535336
rect 99484 528526 99696 528554
rect 97724 492652 97776 492658
rect 97724 492594 97776 492600
rect 99288 492652 99340 492658
rect 99288 492594 99340 492600
rect 97080 491972 97132 491978
rect 97080 491914 97132 491920
rect 96434 491263 96490 491272
rect 96528 491292 96580 491298
rect 96252 490680 96304 490686
rect 96252 490622 96304 490628
rect 96448 489940 96476 491263
rect 96528 491234 96580 491240
rect 97092 489940 97120 491914
rect 97736 489940 97764 492594
rect 99300 491881 99328 492594
rect 99286 491872 99342 491881
rect 99286 491807 99342 491816
rect 99012 491496 99064 491502
rect 99012 491438 99064 491444
rect 98368 491428 98420 491434
rect 98368 491370 98420 491376
rect 98380 489940 98408 491370
rect 99024 489940 99052 491438
rect 99288 491360 99340 491366
rect 99288 491302 99340 491308
rect 91560 489864 91612 489870
rect 91112 489812 91560 489818
rect 91112 489806 91612 489812
rect 91112 489790 91600 489806
rect 99300 489433 99328 491302
rect 99380 490748 99432 490754
rect 99380 490690 99432 490696
rect 99286 489424 99342 489433
rect 99286 489359 99342 489368
rect 69308 460906 69704 460934
rect 69202 451888 69258 451897
rect 69202 451823 69258 451832
rect 69216 451314 69244 451823
rect 69204 451308 69256 451314
rect 69204 451250 69256 451256
rect 69110 437608 69166 437617
rect 69110 437543 69166 437552
rect 69018 434752 69074 434761
rect 69018 434687 69020 434696
rect 69072 434687 69074 434696
rect 69020 434658 69072 434664
rect 69032 433809 69060 434658
rect 69018 433800 69074 433809
rect 69018 433735 69074 433744
rect 69216 428466 69244 451250
rect 69676 440042 69704 460906
rect 99286 443728 99342 443737
rect 99286 443663 99342 443672
rect 72344 440706 72634 440722
rect 93886 440706 94176 440722
rect 72148 440700 72200 440706
rect 72148 440642 72200 440648
rect 72332 440700 72634 440706
rect 72384 440694 72634 440700
rect 92388 440700 92440 440706
rect 72332 440642 72384 440648
rect 93886 440700 94188 440706
rect 93886 440694 94136 440700
rect 92388 440642 92440 440648
rect 69676 440014 70058 440042
rect 69676 431954 69704 440014
rect 70688 433294 70716 440028
rect 71042 438968 71098 438977
rect 71042 438903 71098 438912
rect 70676 433288 70728 433294
rect 70676 433230 70728 433236
rect 69400 431926 69704 431954
rect 69204 428460 69256 428466
rect 69204 428402 69256 428408
rect 69112 400240 69164 400246
rect 69112 400182 69164 400188
rect 69124 376009 69152 400182
rect 69110 376000 69166 376009
rect 69110 375935 69166 375944
rect 69112 375352 69164 375358
rect 69112 375294 69164 375300
rect 69124 374649 69152 375294
rect 69110 374640 69166 374649
rect 69110 374575 69166 374584
rect 68296 364306 68692 364334
rect 68848 364306 68968 364334
rect 68376 349784 68428 349790
rect 68374 349752 68376 349761
rect 68428 349752 68430 349761
rect 68374 349687 68430 349696
rect 68192 346384 68244 346390
rect 68190 346352 68192 346361
rect 68244 346352 68246 346361
rect 68190 346287 68246 346296
rect 68204 346261 68232 346287
rect 68664 345098 68692 364306
rect 68940 353161 68968 364306
rect 68926 353152 68982 353161
rect 68926 353087 68982 353096
rect 68940 352578 68968 353087
rect 68928 352572 68980 352578
rect 68928 352514 68980 352520
rect 68742 351248 68798 351257
rect 68742 351183 68798 351192
rect 68652 345092 68704 345098
rect 68652 345034 68704 345040
rect 68664 345001 68692 345034
rect 68650 344992 68706 345001
rect 68650 344927 68706 344936
rect 67638 343768 67694 343777
rect 67638 343703 67694 343712
rect 67652 343670 67680 343703
rect 67640 343664 67692 343670
rect 67640 343606 67692 343612
rect 67638 342952 67694 342961
rect 67638 342887 67694 342896
rect 67652 342310 67680 342887
rect 67640 342304 67692 342310
rect 67640 342246 67692 342252
rect 68650 341728 68706 341737
rect 68650 341663 68706 341672
rect 67546 341592 67602 341601
rect 68664 341562 68692 341663
rect 67546 341527 67602 341536
rect 68652 341556 68704 341562
rect 68652 341498 68704 341504
rect 67914 340232 67970 340241
rect 67914 340167 67916 340176
rect 67968 340167 67970 340176
rect 67916 340138 67968 340144
rect 68756 329089 68784 351183
rect 68834 349752 68890 349761
rect 68834 349687 68890 349696
rect 68742 329080 68798 329089
rect 68742 329015 68798 329024
rect 67456 323740 67508 323746
rect 67456 323682 67508 323688
rect 68848 322153 68876 349687
rect 68834 322144 68890 322153
rect 68834 322079 68890 322088
rect 67272 320952 67324 320958
rect 67272 320894 67324 320900
rect 65984 320884 66036 320890
rect 65984 320826 66036 320832
rect 65614 302152 65670 302161
rect 65614 302087 65670 302096
rect 65628 288386 65656 302087
rect 65996 290494 66024 320826
rect 69124 313954 69152 374575
rect 69202 370152 69258 370161
rect 69202 370087 69258 370096
rect 69216 319462 69244 370087
rect 69400 364334 69428 431926
rect 71056 401674 71084 438903
rect 71332 438258 71360 440028
rect 71320 438252 71372 438258
rect 71320 438194 71372 438200
rect 71976 437306 72004 440028
rect 72160 437306 72188 440642
rect 71964 437300 72016 437306
rect 71964 437242 72016 437248
rect 72148 437300 72200 437306
rect 72148 437242 72200 437248
rect 72344 431954 72372 440642
rect 73264 435402 73292 440028
rect 73908 438326 73936 440028
rect 73896 438320 73948 438326
rect 73896 438262 73948 438268
rect 73802 437608 73858 437617
rect 73802 437543 73858 437552
rect 73252 435396 73304 435402
rect 73252 435338 73304 435344
rect 71976 431926 72372 431954
rect 70400 401668 70452 401674
rect 70400 401610 70452 401616
rect 71044 401668 71096 401674
rect 71044 401610 71096 401616
rect 69664 396840 69716 396846
rect 69664 396782 69716 396788
rect 69676 371890 69704 396782
rect 69756 387864 69808 387870
rect 69756 387806 69808 387812
rect 69768 385914 69796 387806
rect 70124 387184 70176 387190
rect 70124 387126 70176 387132
rect 69768 385886 70058 385914
rect 70136 373994 70164 387126
rect 70412 385914 70440 401610
rect 71044 398200 71096 398206
rect 71044 398142 71096 398148
rect 71056 389162 71084 398142
rect 71044 389156 71096 389162
rect 71044 389098 71096 389104
rect 71780 388476 71832 388482
rect 71780 388418 71832 388424
rect 71792 385914 71820 388418
rect 71976 387258 72004 431926
rect 72424 396092 72476 396098
rect 72424 396034 72476 396040
rect 72436 389094 72464 396034
rect 72424 389088 72476 389094
rect 72424 389030 72476 389036
rect 71964 387252 72016 387258
rect 71964 387194 72016 387200
rect 72436 385914 72464 389030
rect 73816 387841 73844 437543
rect 74552 433265 74580 440028
rect 75184 439612 75236 439618
rect 75184 439554 75236 439560
rect 74632 436008 74684 436014
rect 74632 435950 74684 435956
rect 74538 433256 74594 433265
rect 74538 433191 74594 433200
rect 73526 387832 73582 387841
rect 73526 387767 73582 387776
rect 73802 387832 73858 387841
rect 73802 387767 73858 387776
rect 73540 385914 73568 387767
rect 74644 387122 74672 435950
rect 75196 393314 75224 439554
rect 75460 438184 75512 438190
rect 75458 438152 75460 438161
rect 75512 438152 75514 438161
rect 75458 438087 75514 438096
rect 75840 436014 75868 440028
rect 75828 436008 75880 436014
rect 75828 435950 75880 435956
rect 76484 433226 76512 440028
rect 76564 436756 76616 436762
rect 76564 436698 76616 436704
rect 76472 433220 76524 433226
rect 76472 433162 76524 433168
rect 76576 402974 76604 436698
rect 77128 435470 77156 440028
rect 77772 437306 77800 440028
rect 78430 440014 78628 440042
rect 77300 437300 77352 437306
rect 77300 437242 77352 437248
rect 77760 437300 77812 437306
rect 77760 437242 77812 437248
rect 77116 435464 77168 435470
rect 77116 435406 77168 435412
rect 76576 402946 76696 402974
rect 74920 393286 75224 393314
rect 74816 389156 74868 389162
rect 74816 389098 74868 389104
rect 74632 387116 74684 387122
rect 74632 387058 74684 387064
rect 74828 386442 74856 389098
rect 74920 388142 74948 393286
rect 75552 391264 75604 391270
rect 75552 391206 75604 391212
rect 75564 390590 75592 391206
rect 75552 390584 75604 390590
rect 75552 390526 75604 390532
rect 74908 388136 74960 388142
rect 74908 388078 74960 388084
rect 74816 386436 74868 386442
rect 74816 386378 74868 386384
rect 74828 385914 74856 386378
rect 70412 385886 70702 385914
rect 71792 385886 71990 385914
rect 72436 385886 72634 385914
rect 73278 385886 73568 385914
rect 74566 385886 74856 385914
rect 74920 385914 74948 388078
rect 75564 385914 75592 390526
rect 76668 386481 76696 402946
rect 77312 396778 77340 437242
rect 78600 434761 78628 440014
rect 78772 438796 78824 438802
rect 78772 438738 78824 438744
rect 78784 437918 78812 438738
rect 78772 437912 78824 437918
rect 78772 437854 78824 437860
rect 78586 434752 78642 434761
rect 78586 434687 78588 434696
rect 78640 434687 78642 434696
rect 78588 434658 78640 434664
rect 77300 396772 77352 396778
rect 77300 396714 77352 396720
rect 77852 394188 77904 394194
rect 77852 394130 77904 394136
rect 76654 386472 76710 386481
rect 76654 386407 76710 386416
rect 76668 385914 76696 386407
rect 77864 385914 77892 394130
rect 78784 394058 78812 437854
rect 79060 437238 79088 440028
rect 79704 437918 79732 440028
rect 79692 437912 79744 437918
rect 79692 437854 79744 437860
rect 80992 437481 81020 440028
rect 81636 437510 81664 440028
rect 82280 438190 82308 440028
rect 82924 438734 82952 440028
rect 83464 439544 83516 439550
rect 83464 439486 83516 439492
rect 82912 438728 82964 438734
rect 82912 438670 82964 438676
rect 82268 438184 82320 438190
rect 82268 438126 82320 438132
rect 81624 437504 81676 437510
rect 80978 437472 81034 437481
rect 81624 437446 81676 437452
rect 82820 437504 82872 437510
rect 82820 437446 82872 437452
rect 80978 437407 81034 437416
rect 78864 437232 78916 437238
rect 78864 437174 78916 437180
rect 79048 437232 79100 437238
rect 79048 437174 79100 437180
rect 78772 394052 78824 394058
rect 78772 393994 78824 394000
rect 78220 391332 78272 391338
rect 78220 391274 78272 391280
rect 78232 390658 78260 391274
rect 78220 390652 78272 390658
rect 78220 390594 78272 390600
rect 74920 385886 75210 385914
rect 75564 385886 75854 385914
rect 76668 385886 77142 385914
rect 77786 385886 77892 385914
rect 77864 385370 77892 385886
rect 78232 385778 78260 390594
rect 78232 385750 78430 385778
rect 78876 385762 78904 437174
rect 80992 436529 81020 437407
rect 81636 437374 81664 437446
rect 81624 437368 81676 437374
rect 81624 437310 81676 437316
rect 80058 436520 80114 436529
rect 80058 436455 80114 436464
rect 80978 436520 81034 436529
rect 80978 436455 81034 436464
rect 80072 402974 80100 436455
rect 80072 402946 80192 402974
rect 80060 390720 80112 390726
rect 80060 390662 80112 390668
rect 79324 389292 79376 389298
rect 79324 389234 79376 389240
rect 79336 385914 79364 389234
rect 80072 385914 80100 390662
rect 80164 387025 80192 402946
rect 81808 395412 81860 395418
rect 81808 395354 81860 395360
rect 81820 394806 81848 395354
rect 81808 394800 81860 394806
rect 81808 394742 81860 394748
rect 80150 387016 80206 387025
rect 80150 386951 80206 386960
rect 80612 386572 80664 386578
rect 80612 386514 80664 386520
rect 80624 385914 80652 386514
rect 81820 385914 81848 394742
rect 82832 389842 82860 437446
rect 82912 434716 82964 434722
rect 82912 434658 82964 434664
rect 82924 431934 82952 434658
rect 82912 431928 82964 431934
rect 82912 431870 82964 431876
rect 83476 394126 83504 439486
rect 83568 438258 83596 440028
rect 84212 438977 84240 440028
rect 84198 438968 84254 438977
rect 84198 438903 84254 438912
rect 83556 438252 83608 438258
rect 83556 438194 83608 438200
rect 84856 438190 84884 440028
rect 85776 440014 86158 440042
rect 85776 439550 85804 440014
rect 85764 439544 85816 439550
rect 85764 439486 85816 439492
rect 84844 438184 84896 438190
rect 84844 438126 84896 438132
rect 86788 437442 86816 440028
rect 87446 440014 87644 440042
rect 87616 438666 87644 440014
rect 87604 438660 87656 438666
rect 87604 438602 87656 438608
rect 86224 437436 86276 437442
rect 86224 437378 86276 437384
rect 86776 437436 86828 437442
rect 86776 437378 86828 437384
rect 86236 400994 86264 437378
rect 86224 400988 86276 400994
rect 86224 400930 86276 400936
rect 84844 395344 84896 395350
rect 84844 395286 84896 395292
rect 84856 394738 84884 395286
rect 84844 394732 84896 394738
rect 84844 394674 84896 394680
rect 85120 394732 85172 394738
rect 85120 394674 85172 394680
rect 83464 394120 83516 394126
rect 83464 394062 83516 394068
rect 83004 393984 83056 393990
rect 83004 393926 83056 393932
rect 83016 393446 83044 393926
rect 83004 393440 83056 393446
rect 83004 393382 83056 393388
rect 82912 392624 82964 392630
rect 82912 392566 82964 392572
rect 82924 392086 82952 392566
rect 82912 392080 82964 392086
rect 82912 392022 82964 392028
rect 82820 389836 82872 389842
rect 82820 389778 82872 389784
rect 83016 385914 83044 393382
rect 83648 392080 83700 392086
rect 83648 392022 83700 392028
rect 79336 385886 79718 385914
rect 80072 385886 80362 385914
rect 80624 385886 81006 385914
rect 81820 385886 82294 385914
rect 82938 385886 83044 385914
rect 83660 385778 83688 392022
rect 84476 390788 84528 390794
rect 84476 390730 84528 390736
rect 84488 385914 84516 390730
rect 85132 385914 85160 394674
rect 86408 388476 86460 388482
rect 86408 388418 86460 388424
rect 86420 385914 86448 388418
rect 87052 388000 87104 388006
rect 87052 387942 87104 387948
rect 84488 385886 84870 385914
rect 85132 385886 85514 385914
rect 86158 385886 86448 385914
rect 87064 385914 87092 387942
rect 87616 387190 87644 438602
rect 88076 438326 88104 440028
rect 88720 439006 88748 440028
rect 89378 440014 89852 440042
rect 89824 439618 89852 440014
rect 89812 439612 89864 439618
rect 89812 439554 89864 439560
rect 88982 439512 89038 439521
rect 88982 439447 89038 439456
rect 88708 439000 88760 439006
rect 88708 438942 88760 438948
rect 88996 438326 89024 439447
rect 88064 438320 88116 438326
rect 88064 438262 88116 438268
rect 88984 438320 89036 438326
rect 88984 438262 89036 438268
rect 87696 404388 87748 404394
rect 87696 404330 87748 404336
rect 87708 394194 87736 404330
rect 88340 395344 88392 395350
rect 88340 395286 88392 395292
rect 87696 394188 87748 394194
rect 87696 394130 87748 394136
rect 88248 392624 88300 392630
rect 88248 392566 88300 392572
rect 87604 387184 87656 387190
rect 87604 387126 87656 387132
rect 88260 385914 88288 392566
rect 87064 385886 87446 385914
rect 88090 385886 88288 385914
rect 88352 385914 88380 395286
rect 88996 387122 89024 438262
rect 89824 392698 89852 439554
rect 90008 438870 90036 440028
rect 90928 440014 91310 440042
rect 91756 440014 91954 440042
rect 90928 439074 90956 440014
rect 90916 439068 90968 439074
rect 90916 439010 90968 439016
rect 89996 438864 90048 438870
rect 89996 438806 90048 438812
rect 91756 436082 91784 440014
rect 91744 436076 91796 436082
rect 91744 436018 91796 436024
rect 91756 399498 91784 436018
rect 91744 399492 91796 399498
rect 91744 399434 91796 399440
rect 90086 398032 90142 398041
rect 90086 397967 90142 397976
rect 89812 392692 89864 392698
rect 89812 392634 89864 392640
rect 88984 387116 89036 387122
rect 88984 387058 89036 387064
rect 90100 385914 90128 397967
rect 92400 392154 92428 440642
rect 93964 440042 93992 440694
rect 94136 440642 94188 440648
rect 92584 438258 92612 440028
rect 93242 440014 93716 440042
rect 93886 440028 93992 440042
rect 92572 438252 92624 438258
rect 92572 438194 92624 438200
rect 93688 437481 93716 440014
rect 93872 440014 93992 440028
rect 93872 438546 93900 440014
rect 93780 438518 93900 438546
rect 93674 437472 93730 437481
rect 93674 437407 93730 437416
rect 93688 400926 93716 437407
rect 93780 402286 93808 438518
rect 94516 437442 94544 440028
rect 94504 437436 94556 437442
rect 94504 437378 94556 437384
rect 93768 402280 93820 402286
rect 93768 402222 93820 402228
rect 93676 400920 93728 400926
rect 93676 400862 93728 400868
rect 94136 398948 94188 398954
rect 94136 398890 94188 398896
rect 91560 392148 91612 392154
rect 91560 392090 91612 392096
rect 92388 392148 92440 392154
rect 92388 392090 92440 392096
rect 91008 388544 91060 388550
rect 91008 388486 91060 388492
rect 91020 385914 91048 388486
rect 91572 385914 91600 392090
rect 94044 390720 94096 390726
rect 94044 390662 94096 390668
rect 92940 387932 92992 387938
rect 92940 387874 92992 387880
rect 92848 387864 92900 387870
rect 92848 387806 92900 387812
rect 92860 385914 92888 387806
rect 88352 385886 88734 385914
rect 90022 385886 90312 385914
rect 90666 385886 91048 385914
rect 91310 385886 91600 385914
rect 92598 385886 92888 385914
rect 92952 385914 92980 387874
rect 94056 385914 94084 390662
rect 92952 385886 93242 385914
rect 93886 385886 94084 385914
rect 94148 385914 94176 398890
rect 94516 396846 94544 437378
rect 95160 437374 95188 440028
rect 96448 438938 96476 440028
rect 96528 439544 96580 439550
rect 96528 439486 96580 439492
rect 96436 438932 96488 438938
rect 96436 438874 96488 438880
rect 95884 438864 95936 438870
rect 95884 438806 95936 438812
rect 95148 437368 95200 437374
rect 95148 437310 95200 437316
rect 94504 396840 94556 396846
rect 94504 396782 94556 396788
rect 95160 396778 95188 437310
rect 95896 396914 95924 438806
rect 96448 438802 96476 438874
rect 96540 438870 96568 439486
rect 96618 438968 96674 438977
rect 96618 438903 96674 438912
rect 96528 438864 96580 438870
rect 96528 438806 96580 438812
rect 96436 438796 96488 438802
rect 96436 438738 96488 438744
rect 96632 403646 96660 438903
rect 97092 438598 97120 440028
rect 97736 439793 97764 440028
rect 97722 439784 97778 439793
rect 97722 439719 97778 439728
rect 97736 438977 97764 439719
rect 97722 438968 97778 438977
rect 97722 438903 97778 438912
rect 97080 438592 97132 438598
rect 97080 438534 97132 438540
rect 97908 438252 97960 438258
rect 97908 438194 97960 438200
rect 97724 438184 97776 438190
rect 97724 438126 97776 438132
rect 97736 436762 97764 438126
rect 97724 436756 97776 436762
rect 97724 436698 97776 436704
rect 96620 403640 96672 403646
rect 96620 403582 96672 403588
rect 95884 396908 95936 396914
rect 95884 396850 95936 396856
rect 95148 396772 95200 396778
rect 95148 396714 95200 396720
rect 97448 392692 97500 392698
rect 97448 392634 97500 392640
rect 96434 389872 96490 389881
rect 96434 389807 96490 389816
rect 96528 389836 96580 389842
rect 96448 389201 96476 389807
rect 96528 389778 96580 389784
rect 95882 389192 95938 389201
rect 95882 389127 95938 389136
rect 96434 389192 96490 389201
rect 96434 389127 96490 389136
rect 95896 385914 95924 389127
rect 96540 385914 96568 389778
rect 97460 385914 97488 392634
rect 97920 388618 97948 438194
rect 98380 437889 98408 440028
rect 99024 438734 99052 440028
rect 99012 438728 99064 438734
rect 99012 438670 99064 438676
rect 99300 437889 99328 443663
rect 98366 437880 98422 437889
rect 98366 437815 98422 437824
rect 99286 437880 99342 437889
rect 99286 437815 99342 437824
rect 98642 398032 98698 398041
rect 98642 397967 98698 397976
rect 98656 397594 98684 397967
rect 98644 397588 98696 397594
rect 98644 397530 98696 397536
rect 98552 393984 98604 393990
rect 98552 393926 98604 393932
rect 98460 388680 98512 388686
rect 98460 388622 98512 388628
rect 97908 388612 97960 388618
rect 97908 388554 97960 388560
rect 98472 385914 98500 388622
rect 94148 385886 94530 385914
rect 95818 385886 95924 385914
rect 96462 385886 96568 385914
rect 97106 385886 97488 385914
rect 98394 385886 98500 385914
rect 98564 385914 98592 393926
rect 98656 388482 98684 397530
rect 99300 394058 99328 437815
rect 99288 394052 99340 394058
rect 99288 393994 99340 394000
rect 98644 388476 98696 388482
rect 98644 388418 98696 388424
rect 99392 385914 99420 490690
rect 99484 444446 99512 528526
rect 99656 491360 99708 491366
rect 99656 491302 99708 491308
rect 99668 489940 99696 491302
rect 99654 484664 99710 484673
rect 99760 484650 99788 535327
rect 99932 491564 99984 491570
rect 99932 491506 99984 491512
rect 99710 484622 99788 484650
rect 99654 484599 99710 484608
rect 99668 484430 99696 484599
rect 99656 484424 99708 484430
rect 99656 484366 99708 484372
rect 99944 484362 99972 491506
rect 99932 484356 99984 484362
rect 99932 484298 99984 484304
rect 99564 472796 99616 472802
rect 99564 472738 99616 472744
rect 99472 444440 99524 444446
rect 99472 444382 99524 444388
rect 99470 443184 99526 443193
rect 99470 443119 99526 443128
rect 99484 438530 99512 443119
rect 99576 442513 99604 472738
rect 101404 464976 101456 464982
rect 101404 464918 101456 464924
rect 100668 454776 100720 454782
rect 100668 454718 100720 454724
rect 99562 442504 99618 442513
rect 99562 442439 99618 442448
rect 99668 438870 99696 440028
rect 99656 438864 99708 438870
rect 99656 438806 99708 438812
rect 99472 438524 99524 438530
rect 99472 438466 99524 438472
rect 98564 385886 99038 385914
rect 99392 385886 100064 385914
rect 78864 385756 78916 385762
rect 83582 385750 83688 385778
rect 78864 385698 78916 385704
rect 77496 385354 77892 385370
rect 90284 385354 90312 385886
rect 100036 385354 100064 385886
rect 100680 385694 100708 454718
rect 100760 444440 100812 444446
rect 100760 444382 100812 444388
rect 100772 440337 100800 444382
rect 100758 440328 100814 440337
rect 100758 440263 100814 440272
rect 101416 438258 101444 464918
rect 101494 451208 101550 451217
rect 101494 451143 101550 451152
rect 101404 438252 101456 438258
rect 101404 438194 101456 438200
rect 101508 431866 101536 451143
rect 101968 447137 101996 536658
rect 102152 495434 102180 537678
rect 102888 537674 102916 540138
rect 103532 537985 103560 540138
rect 103518 537976 103574 537985
rect 103518 537911 103574 537920
rect 102876 537668 102928 537674
rect 102876 537610 102928 537616
rect 102152 495406 102364 495434
rect 102046 491464 102102 491473
rect 102046 491399 102102 491408
rect 102060 489870 102088 491399
rect 102048 489864 102100 489870
rect 102048 489806 102100 489812
rect 101954 447128 102010 447137
rect 101954 447063 102010 447072
rect 101968 445806 101996 447063
rect 101956 445800 102008 445806
rect 101956 445742 102008 445748
rect 101496 431860 101548 431866
rect 101496 431802 101548 431808
rect 101508 429894 101536 431802
rect 101496 429888 101548 429894
rect 101496 429830 101548 429836
rect 101128 396840 101180 396846
rect 101128 396782 101180 396788
rect 101036 389292 101088 389298
rect 101036 389234 101088 389240
rect 101048 385914 101076 389234
rect 100970 385886 101076 385914
rect 101140 385914 101168 396782
rect 102060 389298 102088 489806
rect 102138 485208 102194 485217
rect 102138 485143 102194 485152
rect 102152 485110 102180 485143
rect 102140 485104 102192 485110
rect 102140 485046 102192 485052
rect 102336 484401 102364 495406
rect 102416 492108 102468 492114
rect 102416 492050 102468 492056
rect 102322 484392 102378 484401
rect 102322 484327 102378 484336
rect 102138 483848 102194 483857
rect 102138 483783 102194 483792
rect 102152 483682 102180 483783
rect 102140 483676 102192 483682
rect 102140 483618 102192 483624
rect 102140 482996 102192 483002
rect 102140 482938 102192 482944
rect 102152 482633 102180 482938
rect 102138 482624 102194 482633
rect 102138 482559 102194 482568
rect 102138 481808 102194 481817
rect 102138 481743 102194 481752
rect 102152 481710 102180 481743
rect 102140 481704 102192 481710
rect 102140 481646 102192 481652
rect 102324 481636 102376 481642
rect 102324 481578 102376 481584
rect 102138 481264 102194 481273
rect 102138 481199 102194 481208
rect 102152 480962 102180 481199
rect 102336 481137 102364 481578
rect 102322 481128 102378 481137
rect 102322 481063 102378 481072
rect 102140 480956 102192 480962
rect 102140 480898 102192 480904
rect 102428 480254 102456 492050
rect 103426 489288 103482 489297
rect 103426 489223 103482 489232
rect 103440 489190 103468 489223
rect 103428 489184 103480 489190
rect 103428 489126 103480 489132
rect 103428 488504 103480 488510
rect 103426 488472 103428 488481
rect 103480 488472 103482 488481
rect 103426 488407 103482 488416
rect 103426 487928 103482 487937
rect 103426 487863 103482 487872
rect 103440 487830 103468 487863
rect 103428 487824 103480 487830
rect 103428 487766 103480 487772
rect 103428 487144 103480 487150
rect 103428 487086 103480 487092
rect 103440 486713 103468 487086
rect 103426 486704 103482 486713
rect 103426 486639 103482 486648
rect 103426 486568 103482 486577
rect 103426 486503 103482 486512
rect 103440 486470 103468 486503
rect 103428 486464 103480 486470
rect 103428 486406 103480 486412
rect 103520 484356 103572 484362
rect 103520 484298 103572 484304
rect 102244 480226 102456 480254
rect 102140 480208 102192 480214
rect 102140 480150 102192 480156
rect 102152 479913 102180 480150
rect 102138 479904 102194 479913
rect 102138 479839 102194 479848
rect 102138 479768 102194 479777
rect 102138 479703 102140 479712
rect 102192 479703 102194 479712
rect 102140 479674 102192 479680
rect 102138 477864 102194 477873
rect 102138 477799 102194 477808
rect 102152 477562 102180 477799
rect 102140 477556 102192 477562
rect 102140 477498 102192 477504
rect 102140 477420 102192 477426
rect 102140 477362 102192 477368
rect 102152 477057 102180 477362
rect 102138 477048 102194 477057
rect 102138 476983 102194 476992
rect 102140 475924 102192 475930
rect 102140 475866 102192 475872
rect 102152 475697 102180 475866
rect 102138 475688 102194 475697
rect 102138 475623 102194 475632
rect 102140 474700 102192 474706
rect 102140 474642 102192 474648
rect 102152 474337 102180 474642
rect 102138 474328 102194 474337
rect 102138 474263 102194 474272
rect 102138 472968 102194 472977
rect 102138 472903 102194 472912
rect 102152 472666 102180 472903
rect 102140 472660 102192 472666
rect 102140 472602 102192 472608
rect 102140 471980 102192 471986
rect 102140 471922 102192 471928
rect 102152 471617 102180 471922
rect 102138 471608 102194 471617
rect 102138 471543 102194 471552
rect 102140 470552 102192 470558
rect 102140 470494 102192 470500
rect 102152 470257 102180 470494
rect 102138 470248 102194 470257
rect 102138 470183 102194 470192
rect 102138 466848 102194 466857
rect 102138 466783 102194 466792
rect 102152 466546 102180 466783
rect 102140 466540 102192 466546
rect 102140 466482 102192 466488
rect 102140 466404 102192 466410
rect 102140 466346 102192 466352
rect 102152 466177 102180 466346
rect 102138 466168 102194 466177
rect 102138 466103 102194 466112
rect 102140 465724 102192 465730
rect 102140 465666 102192 465672
rect 102152 465633 102180 465666
rect 102138 465624 102194 465633
rect 102138 465559 102194 465568
rect 102140 465044 102192 465050
rect 102140 464986 102192 464992
rect 102152 464817 102180 464986
rect 102244 464982 102272 480226
rect 102324 477488 102376 477494
rect 102324 477430 102376 477436
rect 102336 476513 102364 477430
rect 102414 477184 102470 477193
rect 102414 477119 102470 477128
rect 102322 476504 102378 476513
rect 102322 476439 102378 476448
rect 102428 476066 102456 477119
rect 102416 476060 102468 476066
rect 102416 476002 102468 476008
rect 103428 476060 103480 476066
rect 103428 476002 103480 476008
rect 102324 475992 102376 475998
rect 102324 475934 102376 475940
rect 102336 475153 102364 475934
rect 102322 475144 102378 475153
rect 102322 475079 102378 475088
rect 102324 473340 102376 473346
rect 102324 473282 102376 473288
rect 102336 472433 102364 473282
rect 102322 472424 102378 472433
rect 102322 472359 102378 472368
rect 102876 471300 102928 471306
rect 102876 471242 102928 471248
rect 102322 470928 102378 470937
rect 102322 470863 102378 470872
rect 102336 470626 102364 470863
rect 102324 470620 102376 470626
rect 102324 470562 102376 470568
rect 102888 469713 102916 471242
rect 102874 469704 102930 469713
rect 102874 469639 102930 469648
rect 103150 466984 103206 466993
rect 103150 466919 103206 466928
rect 103164 466478 103192 466919
rect 103152 466472 103204 466478
rect 103152 466414 103204 466420
rect 103336 465724 103388 465730
rect 103336 465666 103388 465672
rect 102232 464976 102284 464982
rect 102232 464918 102284 464924
rect 102138 464808 102194 464817
rect 102138 464743 102194 464752
rect 102140 464160 102192 464166
rect 102138 464128 102140 464137
rect 102192 464128 102194 464137
rect 102138 464063 102194 464072
rect 102140 463684 102192 463690
rect 102140 463626 102192 463632
rect 102152 463457 102180 463626
rect 102138 463448 102194 463457
rect 102138 463383 102194 463392
rect 102232 462324 102284 462330
rect 102232 462266 102284 462272
rect 102140 462256 102192 462262
rect 102140 462198 102192 462204
rect 102152 462097 102180 462198
rect 102138 462088 102194 462097
rect 102138 462023 102194 462032
rect 102244 461553 102272 462266
rect 102230 461544 102286 461553
rect 102230 461479 102286 461488
rect 102140 460896 102192 460902
rect 102140 460838 102192 460844
rect 102152 460193 102180 460838
rect 102230 460728 102286 460737
rect 102230 460663 102286 460672
rect 102138 460184 102194 460193
rect 102138 460119 102194 460128
rect 102244 459610 102272 460663
rect 102232 459604 102284 459610
rect 102232 459546 102284 459552
rect 102140 459468 102192 459474
rect 102140 459410 102192 459416
rect 102152 459377 102180 459410
rect 102138 459368 102194 459377
rect 102138 459303 102194 459312
rect 103242 458688 103298 458697
rect 103242 458623 103298 458632
rect 103256 458182 103284 458623
rect 103244 458176 103296 458182
rect 103244 458118 103296 458124
rect 102140 458108 102192 458114
rect 102140 458050 102192 458056
rect 102152 458017 102180 458050
rect 102138 458008 102194 458017
rect 102138 457943 102194 457952
rect 102140 456748 102192 456754
rect 102140 456690 102192 456696
rect 102152 456657 102180 456690
rect 102232 456680 102284 456686
rect 102138 456648 102194 456657
rect 102232 456622 102284 456628
rect 102138 456583 102194 456592
rect 102244 456113 102272 456622
rect 102230 456104 102286 456113
rect 102230 456039 102286 456048
rect 102140 455388 102192 455394
rect 102140 455330 102192 455336
rect 102152 455297 102180 455330
rect 102138 455288 102194 455297
rect 102138 455223 102194 455232
rect 102140 454844 102192 454850
rect 102140 454786 102192 454792
rect 102152 454617 102180 454786
rect 102138 454608 102194 454617
rect 102138 454543 102194 454552
rect 102874 453384 102930 453393
rect 102874 453319 102876 453328
rect 102928 453319 102930 453328
rect 102876 453290 102928 453296
rect 102140 453280 102192 453286
rect 102138 453248 102140 453257
rect 102192 453248 102194 453257
rect 102138 453183 102194 453192
rect 102140 452600 102192 452606
rect 102138 452568 102140 452577
rect 102192 452568 102194 452577
rect 102138 452503 102194 452512
rect 102140 449880 102192 449886
rect 102140 449822 102192 449828
rect 102152 449313 102180 449822
rect 102138 449304 102194 449313
rect 102138 449239 102194 449248
rect 102232 448520 102284 448526
rect 102138 448488 102194 448497
rect 102232 448462 102284 448468
rect 102138 448423 102140 448432
rect 102192 448423 102194 448432
rect 102140 448394 102192 448400
rect 102244 447953 102272 448462
rect 102230 447944 102286 447953
rect 102230 447879 102286 447888
rect 103152 445120 103204 445126
rect 103150 445088 103152 445097
rect 103204 445088 103206 445097
rect 102600 445052 102652 445058
rect 103150 445023 103206 445032
rect 102600 444994 102652 445000
rect 102612 443193 102640 444994
rect 102598 443184 102654 443193
rect 102598 443119 102654 443128
rect 102690 442504 102746 442513
rect 102690 442439 102746 442448
rect 102704 441726 102732 442439
rect 103150 441824 103206 441833
rect 103150 441759 103206 441768
rect 102692 441720 102744 441726
rect 102692 441662 102744 441668
rect 103164 441658 103192 441759
rect 103152 441652 103204 441658
rect 103152 441594 103204 441600
rect 103150 440872 103206 440881
rect 103150 440807 103206 440816
rect 103164 440366 103192 440807
rect 103152 440360 103204 440366
rect 102138 440328 102194 440337
rect 103152 440302 103204 440308
rect 102138 440263 102140 440272
rect 102192 440263 102194 440272
rect 102140 440234 102192 440240
rect 103256 389910 103284 458118
rect 103348 394126 103376 465666
rect 103336 394120 103388 394126
rect 103336 394062 103388 394068
rect 103440 391241 103468 476002
rect 103532 402974 103560 484298
rect 103612 469872 103664 469878
rect 103612 469814 103664 469820
rect 103624 469033 103652 469814
rect 103610 469024 103666 469033
rect 103610 468959 103666 468968
rect 103612 451920 103664 451926
rect 103612 451862 103664 451868
rect 103624 450673 103652 451862
rect 103704 451716 103756 451722
rect 103704 451658 103756 451664
rect 103610 450664 103666 450673
rect 103610 450599 103666 450608
rect 103716 449857 103744 451658
rect 103702 449848 103758 449857
rect 103702 449783 103758 449792
rect 104176 445874 104204 540138
rect 104820 538121 104848 540138
rect 105478 540110 105584 540138
rect 104806 538112 104862 538121
rect 104806 538047 104862 538056
rect 105556 536722 105584 540110
rect 105544 536716 105596 536722
rect 105544 536658 105596 536664
rect 105740 534074 105768 548383
rect 105556 534046 105768 534074
rect 104900 489932 104952 489938
rect 104900 489874 104952 489880
rect 104254 449848 104310 449857
rect 104254 449783 104310 449792
rect 104164 445868 104216 445874
rect 104164 445810 104216 445816
rect 104176 445126 104204 445810
rect 104164 445120 104216 445126
rect 104164 445062 104216 445068
rect 104162 444408 104218 444417
rect 104162 444343 104218 444352
rect 103532 402946 103836 402974
rect 103426 391232 103482 391241
rect 103426 391167 103482 391176
rect 103244 389904 103296 389910
rect 103244 389846 103296 389852
rect 102048 389292 102100 389298
rect 102048 389234 102100 389240
rect 102600 389224 102652 389230
rect 102600 389166 102652 389172
rect 102612 385914 102640 389166
rect 103808 386510 103836 402946
rect 104176 401062 104204 444343
rect 104268 403714 104296 449783
rect 104256 403708 104308 403714
rect 104256 403650 104308 403656
rect 104164 401056 104216 401062
rect 104164 400998 104216 401004
rect 104532 389360 104584 389366
rect 104532 389302 104584 389308
rect 103888 386572 103940 386578
rect 103888 386514 103940 386520
rect 103796 386504 103848 386510
rect 103796 386446 103848 386452
rect 103900 385914 103928 386514
rect 103980 386504 104032 386510
rect 103980 386446 104032 386452
rect 101140 385886 101614 385914
rect 102258 385886 102640 385914
rect 103546 385886 103928 385914
rect 103992 385914 104020 386446
rect 104544 385914 104572 389302
rect 104912 386374 104940 489874
rect 104990 479768 105046 479777
rect 104990 479703 104992 479712
rect 105044 479703 105046 479712
rect 104992 479674 105044 479680
rect 105556 456686 105584 534046
rect 106200 486470 106228 577759
rect 106292 560425 106320 698906
rect 106464 594108 106516 594114
rect 106464 594050 106516 594056
rect 106370 564496 106426 564505
rect 106370 564431 106426 564440
rect 106278 560416 106334 560425
rect 106278 560351 106334 560360
rect 106188 486464 106240 486470
rect 106188 486406 106240 486412
rect 106188 479732 106240 479738
rect 106188 479674 106240 479680
rect 106200 476814 106228 479674
rect 106188 476808 106240 476814
rect 106188 476750 106240 476756
rect 105636 474904 105688 474910
rect 105636 474846 105688 474852
rect 105648 464166 105676 474846
rect 106384 473346 106412 564431
rect 106476 540705 106504 594050
rect 108960 586514 108988 702510
rect 108776 586486 108988 586514
rect 106922 583944 106978 583953
rect 106922 583879 106978 583888
rect 106936 560998 106964 583879
rect 107660 582412 107712 582418
rect 107660 582354 107712 582360
rect 107672 573345 107700 582354
rect 108210 580136 108266 580145
rect 108210 580071 108266 580080
rect 108224 579698 108252 580071
rect 108212 579692 108264 579698
rect 108212 579634 108264 579640
rect 108776 577425 108804 586486
rect 109040 582684 109092 582690
rect 109040 582626 109092 582632
rect 108948 581732 109000 581738
rect 108948 581674 109000 581680
rect 108960 581126 108988 581674
rect 108948 581120 109000 581126
rect 108948 581062 109000 581068
rect 108854 579456 108910 579465
rect 108854 579391 108910 579400
rect 108868 578338 108896 579391
rect 108946 578776 109002 578785
rect 108946 578711 109002 578720
rect 108856 578332 108908 578338
rect 108856 578274 108908 578280
rect 108960 578270 108988 578711
rect 108948 578264 109000 578270
rect 108948 578206 109000 578212
rect 108762 577416 108818 577425
rect 108762 577351 108818 577360
rect 108946 576056 109002 576065
rect 108946 575991 109002 576000
rect 108960 575550 108988 575991
rect 108948 575544 109000 575550
rect 108948 575486 109000 575492
rect 108946 574696 109002 574705
rect 108946 574631 109002 574640
rect 108960 574122 108988 574631
rect 108948 574116 109000 574122
rect 108948 574058 109000 574064
rect 108946 574016 109002 574025
rect 108946 573951 109002 573960
rect 108960 573374 108988 573951
rect 108948 573368 109000 573374
rect 107658 573336 107714 573345
rect 107658 573271 107714 573280
rect 108670 573336 108726 573345
rect 108948 573310 109000 573316
rect 108670 573271 108726 573280
rect 108684 573034 108712 573271
rect 108672 573028 108724 573034
rect 108672 572970 108724 572976
rect 108946 572792 109002 572801
rect 108946 572727 108948 572736
rect 109000 572727 109002 572736
rect 108948 572698 109000 572704
rect 108946 571976 109002 571985
rect 108946 571911 109002 571920
rect 108960 571402 108988 571911
rect 108948 571396 109000 571402
rect 108948 571338 109000 571344
rect 108946 570072 109002 570081
rect 108946 570007 109002 570016
rect 108960 569974 108988 570007
rect 108948 569968 109000 569974
rect 108948 569910 109000 569916
rect 107658 569256 107714 569265
rect 107658 569191 107714 569200
rect 107672 568682 107700 569191
rect 107660 568676 107712 568682
rect 107660 568618 107712 568624
rect 108946 567896 109002 567905
rect 108946 567831 109002 567840
rect 108960 567594 108988 567831
rect 108948 567588 109000 567594
rect 108948 567530 109000 567536
rect 108948 567248 109000 567254
rect 108946 567216 108948 567225
rect 109000 567216 109002 567225
rect 108946 567151 109002 567160
rect 108854 566536 108910 566545
rect 108854 566471 108910 566480
rect 108868 565962 108896 566471
rect 108856 565956 108908 565962
rect 108856 565898 108908 565904
rect 108948 565888 109000 565894
rect 108946 565856 108948 565865
rect 109000 565856 109002 565865
rect 108946 565791 109002 565800
rect 108854 565176 108910 565185
rect 108854 565111 108910 565120
rect 108868 564466 108896 565111
rect 108856 564460 108908 564466
rect 108856 564402 108908 564408
rect 108948 564392 109000 564398
rect 108948 564334 109000 564340
rect 108960 563961 108988 564334
rect 108946 563952 109002 563961
rect 108946 563887 109002 563896
rect 108946 562456 109002 562465
rect 108946 562391 109002 562400
rect 108960 561746 108988 562391
rect 108948 561740 109000 561746
rect 108948 561682 109000 561688
rect 108946 561096 109002 561105
rect 108946 561031 109002 561040
rect 106924 560992 106976 560998
rect 106924 560934 106976 560940
rect 107658 560416 107714 560425
rect 107658 560351 107660 560360
rect 107712 560351 107714 560360
rect 107660 560322 107712 560328
rect 108960 560318 108988 561031
rect 108948 560312 109000 560318
rect 108948 560254 109000 560260
rect 108854 559736 108910 559745
rect 108854 559671 108910 559680
rect 108868 558958 108896 559671
rect 108946 559056 109002 559065
rect 108946 558991 108948 559000
rect 109000 558991 109002 559000
rect 108948 558962 109000 558968
rect 108856 558952 108908 558958
rect 108856 558894 108908 558900
rect 108946 558376 109002 558385
rect 108946 558311 109002 558320
rect 108960 557802 108988 558311
rect 108948 557796 109000 557802
rect 108948 557738 109000 557744
rect 107750 557696 107806 557705
rect 107750 557631 107806 557640
rect 107014 552256 107070 552265
rect 107014 552191 107070 552200
rect 106922 542056 106978 542065
rect 106922 541991 106978 542000
rect 106462 540696 106518 540705
rect 106462 540631 106518 540640
rect 106830 540696 106886 540705
rect 106830 540631 106886 540640
rect 106844 539646 106872 540631
rect 106832 539640 106884 539646
rect 106832 539582 106884 539588
rect 106372 473340 106424 473346
rect 106372 473282 106424 473288
rect 105636 464160 105688 464166
rect 105636 464102 105688 464108
rect 105544 456680 105596 456686
rect 105544 456622 105596 456628
rect 105544 456000 105596 456006
rect 105544 455942 105596 455948
rect 105556 438666 105584 455942
rect 105544 438660 105596 438666
rect 105544 438602 105596 438608
rect 105648 394194 105676 464102
rect 106188 456816 106240 456822
rect 106188 456758 106240 456764
rect 106200 456686 106228 456758
rect 106188 456680 106240 456686
rect 106188 456622 106240 456628
rect 106188 454708 106240 454714
rect 106188 454650 106240 454656
rect 106200 453286 106228 454650
rect 106188 453280 106240 453286
rect 106188 453222 106240 453228
rect 106936 449954 106964 541991
rect 107028 460970 107056 552191
rect 107658 551576 107714 551585
rect 107658 551511 107714 551520
rect 107672 550730 107700 551511
rect 107660 550724 107712 550730
rect 107660 550666 107712 550672
rect 107658 546816 107714 546825
rect 107658 546751 107714 546760
rect 107568 473340 107620 473346
rect 107568 473282 107620 473288
rect 107580 472734 107608 473282
rect 107568 472728 107620 472734
rect 107568 472670 107620 472676
rect 107566 470656 107622 470665
rect 107566 470591 107568 470600
rect 107620 470591 107622 470600
rect 107568 470562 107620 470568
rect 107568 462392 107620 462398
rect 107568 462334 107620 462340
rect 107580 462262 107608 462334
rect 107568 462256 107620 462262
rect 107568 462198 107620 462204
rect 107016 460964 107068 460970
rect 107016 460906 107068 460912
rect 107476 459604 107528 459610
rect 107476 459546 107528 459552
rect 107488 451274 107516 459546
rect 107568 458856 107620 458862
rect 107568 458798 107620 458804
rect 107580 458114 107608 458798
rect 107568 458108 107620 458114
rect 107568 458050 107620 458056
rect 107672 455394 107700 546751
rect 107764 465730 107792 557631
rect 108946 557016 109002 557025
rect 108946 556951 109002 556960
rect 107934 556336 107990 556345
rect 107934 556271 107990 556280
rect 107842 543416 107898 543425
rect 107842 543351 107898 543360
rect 107856 542434 107884 543351
rect 107844 542428 107896 542434
rect 107844 542370 107896 542376
rect 107842 542328 107898 542337
rect 107842 542263 107898 542272
rect 107752 465724 107804 465730
rect 107752 465666 107804 465672
rect 107660 455388 107712 455394
rect 107660 455330 107712 455336
rect 107672 454850 107700 455330
rect 107660 454844 107712 454850
rect 107660 454786 107712 454792
rect 107856 451722 107884 542263
rect 107948 474910 107976 556271
rect 108960 556238 108988 556951
rect 108948 556232 109000 556238
rect 108948 556174 109000 556180
rect 108856 556164 108908 556170
rect 108856 556106 108908 556112
rect 108868 555801 108896 556106
rect 108854 555792 108910 555801
rect 108854 555727 108910 555736
rect 108946 554296 109002 554305
rect 108946 554231 109002 554240
rect 108960 553450 108988 554231
rect 108948 553444 109000 553450
rect 108948 553386 109000 553392
rect 108946 552936 109002 552945
rect 108946 552871 109002 552880
rect 108960 552090 108988 552871
rect 108948 552084 109000 552090
rect 108948 552026 109000 552032
rect 108946 550896 109002 550905
rect 108946 550831 109002 550840
rect 108960 550662 108988 550831
rect 108948 550656 109000 550662
rect 108948 550598 109000 550604
rect 108854 550216 108910 550225
rect 108854 550151 108910 550160
rect 108868 549370 108896 550151
rect 108946 549536 109002 549545
rect 108946 549471 109002 549480
rect 108856 549364 108908 549370
rect 108856 549306 108908 549312
rect 108960 549302 108988 549471
rect 108948 549296 109000 549302
rect 108948 549238 109000 549244
rect 108946 547496 109002 547505
rect 108946 547431 109002 547440
rect 108960 546514 108988 547431
rect 108948 546508 109000 546514
rect 108948 546450 109000 546456
rect 108946 546136 109002 546145
rect 108946 546071 109002 546080
rect 108960 545766 108988 546071
rect 108948 545760 109000 545766
rect 108948 545702 109000 545708
rect 108946 545456 109002 545465
rect 108946 545391 109002 545400
rect 108960 545154 108988 545391
rect 108948 545148 109000 545154
rect 108948 545090 109000 545096
rect 108946 544776 109002 544785
rect 108946 544711 109002 544720
rect 108960 544406 108988 544711
rect 108948 544400 109000 544406
rect 108948 544342 109000 544348
rect 108946 544096 109002 544105
rect 108946 544031 109002 544040
rect 108960 543794 108988 544031
rect 108948 543788 109000 543794
rect 108948 543730 109000 543736
rect 108304 540796 108356 540802
rect 108304 540738 108356 540744
rect 108316 540025 108344 540738
rect 108302 540016 108358 540025
rect 108302 539951 108358 539960
rect 109052 489870 109080 582626
rect 109130 581768 109186 581777
rect 109130 581703 109186 581712
rect 109144 539034 109172 581703
rect 109696 540802 109724 703122
rect 111064 703112 111116 703118
rect 111064 703054 111116 703060
rect 110420 584044 110472 584050
rect 110420 583986 110472 583992
rect 109776 568676 109828 568682
rect 109776 568618 109828 568624
rect 109684 540796 109736 540802
rect 109684 540738 109736 540744
rect 109132 539028 109184 539034
rect 109132 538970 109184 538976
rect 109684 538280 109736 538286
rect 109684 538222 109736 538228
rect 109696 537849 109724 538222
rect 109682 537840 109738 537849
rect 109682 537775 109738 537784
rect 109314 491600 109370 491609
rect 109314 491535 109370 491544
rect 109132 490612 109184 490618
rect 109132 490554 109184 490560
rect 109040 489864 109092 489870
rect 109040 489806 109092 489812
rect 109038 489424 109094 489433
rect 109038 489359 109094 489368
rect 109052 488442 109080 489359
rect 109040 488436 109092 488442
rect 109040 488378 109092 488384
rect 107936 474904 107988 474910
rect 107936 474846 107988 474852
rect 108488 464432 108540 464438
rect 108488 464374 108540 464380
rect 108304 455388 108356 455394
rect 108304 455330 108356 455336
rect 107844 451716 107896 451722
rect 107844 451658 107896 451664
rect 107488 451246 107608 451274
rect 106924 449948 106976 449954
rect 106924 449890 106976 449896
rect 107474 449440 107530 449449
rect 107474 449375 107530 449384
rect 106188 449200 106240 449206
rect 106188 449142 106240 449148
rect 106200 448458 106228 449142
rect 107488 448633 107516 449375
rect 107474 448624 107530 448633
rect 107474 448559 107530 448568
rect 107488 448526 107516 448559
rect 107476 448520 107528 448526
rect 107476 448462 107528 448468
rect 106188 448452 106240 448458
rect 106188 448394 106240 448400
rect 107476 448112 107528 448118
rect 107476 448054 107528 448060
rect 107384 436756 107436 436762
rect 107384 436698 107436 436704
rect 107016 398880 107068 398886
rect 107016 398822 107068 398828
rect 105636 394188 105688 394194
rect 105636 394130 105688 394136
rect 106924 388476 106976 388482
rect 106924 388418 106976 388424
rect 104900 386368 104952 386374
rect 104900 386310 104952 386316
rect 105912 386368 105964 386374
rect 105912 386310 105964 386316
rect 103992 385886 104190 385914
rect 104544 385886 104834 385914
rect 105924 385778 105952 386310
rect 106936 385914 106964 388418
rect 106766 385886 106964 385914
rect 107028 385914 107056 398822
rect 107396 387190 107424 436698
rect 107488 390522 107516 448054
rect 107580 399566 107608 451246
rect 107568 399560 107620 399566
rect 107568 399502 107620 399508
rect 108316 398206 108344 455330
rect 108396 445868 108448 445874
rect 108396 445810 108448 445816
rect 108408 398274 108436 445810
rect 108500 436762 108528 464374
rect 109144 456006 109172 490554
rect 109328 489870 109356 491535
rect 109316 489864 109368 489870
rect 109316 489806 109368 489812
rect 109788 478922 109816 568618
rect 110432 493474 110460 583986
rect 110512 582616 110564 582622
rect 110512 582558 110564 582564
rect 110420 493468 110472 493474
rect 110420 493410 110472 493416
rect 110524 492046 110552 582558
rect 110604 572824 110656 572830
rect 110604 572766 110656 572772
rect 110616 556170 110644 572766
rect 110604 556164 110656 556170
rect 110604 556106 110656 556112
rect 110616 555490 110644 556106
rect 110604 555484 110656 555490
rect 110604 555426 110656 555432
rect 110696 550724 110748 550730
rect 110696 550666 110748 550672
rect 110604 537736 110656 537742
rect 110604 537678 110656 537684
rect 110512 492040 110564 492046
rect 110512 491982 110564 491988
rect 110420 491496 110472 491502
rect 110420 491438 110472 491444
rect 110432 491230 110460 491438
rect 110420 491224 110472 491230
rect 110420 491166 110472 491172
rect 110328 488436 110380 488442
rect 110328 488378 110380 488384
rect 109776 478916 109828 478922
rect 109776 478858 109828 478864
rect 109788 477426 109816 478858
rect 109776 477420 109828 477426
rect 109776 477362 109828 477368
rect 109132 456000 109184 456006
rect 109132 455942 109184 455948
rect 108488 436756 108540 436762
rect 108488 436698 108540 436704
rect 108396 398268 108448 398274
rect 108396 398210 108448 398216
rect 108304 398200 108356 398206
rect 108304 398142 108356 398148
rect 109408 391672 109460 391678
rect 109408 391614 109460 391620
rect 107476 390516 107528 390522
rect 107476 390458 107528 390464
rect 109420 388686 109448 391614
rect 109408 388680 109460 388686
rect 109408 388622 109460 388628
rect 110340 387938 110368 488378
rect 110616 472802 110644 537678
rect 110708 529242 110736 550666
rect 111076 538218 111104 703054
rect 115848 702908 115900 702914
rect 115848 702850 115900 702856
rect 113088 702704 113140 702710
rect 113088 702646 113140 702652
rect 112076 585812 112128 585818
rect 112076 585754 112128 585760
rect 112088 584361 112116 585754
rect 111890 584352 111946 584361
rect 111890 584287 111946 584296
rect 112074 584352 112130 584361
rect 112074 584287 112130 584296
rect 111800 579692 111852 579698
rect 111800 579634 111852 579640
rect 111064 538212 111116 538218
rect 111064 538154 111116 538160
rect 110696 529236 110748 529242
rect 110696 529178 110748 529184
rect 110708 528630 110736 529178
rect 110696 528624 110748 528630
rect 110696 528566 110748 528572
rect 110696 494080 110748 494086
rect 110696 494022 110748 494028
rect 110604 472796 110656 472802
rect 110604 472738 110656 472744
rect 110604 395412 110656 395418
rect 110604 395354 110656 395360
rect 110616 394874 110644 395354
rect 110604 394868 110656 394874
rect 110604 394810 110656 394816
rect 109592 387932 109644 387938
rect 109592 387874 109644 387880
rect 110328 387932 110380 387938
rect 110328 387874 110380 387880
rect 108948 387864 109000 387870
rect 108948 387806 109000 387812
rect 107384 387184 107436 387190
rect 107384 387126 107436 387132
rect 108960 385914 108988 387806
rect 109604 385914 109632 387874
rect 110328 386504 110380 386510
rect 110328 386446 110380 386452
rect 110340 385914 110368 386446
rect 110616 386050 110644 394810
rect 110708 391678 110736 494022
rect 111708 491224 111760 491230
rect 111708 491166 111760 491172
rect 110696 391672 110748 391678
rect 110696 391614 110748 391620
rect 110708 391270 110736 391614
rect 110696 391264 110748 391270
rect 110696 391206 110748 391212
rect 111720 390794 111748 491166
rect 111812 488510 111840 579634
rect 111904 495038 111932 584287
rect 112352 545760 112404 545766
rect 112350 545728 112352 545737
rect 113100 545737 113128 702646
rect 113272 586696 113324 586702
rect 113272 586638 113324 586644
rect 113180 573028 113232 573034
rect 113180 572970 113232 572976
rect 112404 545728 112406 545737
rect 112350 545663 112406 545672
rect 113086 545728 113142 545737
rect 113086 545663 113142 545672
rect 111984 532092 112036 532098
rect 111984 532034 112036 532040
rect 111892 495032 111944 495038
rect 111892 494974 111944 494980
rect 111800 488504 111852 488510
rect 111800 488446 111852 488452
rect 111812 487898 111840 488446
rect 111800 487892 111852 487898
rect 111800 487834 111852 487840
rect 111798 485752 111854 485761
rect 111798 485687 111854 485696
rect 111812 485110 111840 485687
rect 111800 485104 111852 485110
rect 111800 485046 111852 485052
rect 111996 464438 112024 532034
rect 112076 495508 112128 495514
rect 112076 495450 112128 495456
rect 111984 464432 112036 464438
rect 111984 464374 112036 464380
rect 112088 440978 112116 495450
rect 112442 488064 112498 488073
rect 112442 487999 112498 488008
rect 112076 440972 112128 440978
rect 112076 440914 112128 440920
rect 111708 390788 111760 390794
rect 111708 390730 111760 390736
rect 111800 388612 111852 388618
rect 111800 388554 111852 388560
rect 111812 387025 111840 388554
rect 112456 388074 112484 487999
rect 112628 485104 112680 485110
rect 112628 485046 112680 485052
rect 112640 484430 112668 485046
rect 112536 484424 112588 484430
rect 112536 484366 112588 484372
rect 112628 484424 112680 484430
rect 112628 484366 112680 484372
rect 112548 479534 112576 484366
rect 113192 480962 113220 572970
rect 113284 496194 113312 586638
rect 113364 583908 113416 583914
rect 113364 583850 113416 583856
rect 113272 496188 113324 496194
rect 113272 496130 113324 496136
rect 113376 493474 113404 583850
rect 114560 583772 114612 583778
rect 114560 583714 114612 583720
rect 113548 498908 113600 498914
rect 113548 498850 113600 498856
rect 113364 493468 113416 493474
rect 113364 493410 113416 493416
rect 113456 491428 113508 491434
rect 113456 491370 113508 491376
rect 113364 490680 113416 490686
rect 113364 490622 113416 490628
rect 113180 480956 113232 480962
rect 113180 480898 113232 480904
rect 112536 479528 112588 479534
rect 112536 479470 112588 479476
rect 112628 470620 112680 470626
rect 112628 470562 112680 470568
rect 112536 441720 112588 441726
rect 112536 441662 112588 441668
rect 112548 391338 112576 441662
rect 112640 402974 112668 470562
rect 113192 454782 113220 480898
rect 113180 454776 113232 454782
rect 113180 454718 113232 454724
rect 113376 438598 113404 490622
rect 113468 448118 113496 491370
rect 113456 448112 113508 448118
rect 113456 448054 113508 448060
rect 113560 439618 113588 498850
rect 114468 492108 114520 492114
rect 114468 492050 114520 492056
rect 114480 491434 114508 492050
rect 114468 491428 114520 491434
rect 114468 491370 114520 491376
rect 114572 491366 114600 583714
rect 114744 567588 114796 567594
rect 114744 567530 114796 567536
rect 114652 557796 114704 557802
rect 114652 557738 114704 557744
rect 114560 491360 114612 491366
rect 114560 491302 114612 491308
rect 114572 487558 114600 491302
rect 114560 487552 114612 487558
rect 114560 487494 114612 487500
rect 114664 466274 114692 557738
rect 114756 477494 114784 567530
rect 115860 544406 115888 702850
rect 117228 702772 117280 702778
rect 117228 702714 117280 702720
rect 115940 585404 115992 585410
rect 115940 585346 115992 585352
rect 115848 544400 115900 544406
rect 115848 544342 115900 544348
rect 115952 534818 115980 585346
rect 116032 583976 116084 583982
rect 116032 583918 116084 583924
rect 115940 534812 115992 534818
rect 115940 534754 115992 534760
rect 114834 500440 114890 500449
rect 114834 500375 114890 500384
rect 114848 499594 114876 500375
rect 114836 499588 114888 499594
rect 114836 499530 114888 499536
rect 114836 495032 114888 495038
rect 114836 494974 114888 494980
rect 114744 477488 114796 477494
rect 114744 477430 114796 477436
rect 114652 466268 114704 466274
rect 114652 466210 114704 466216
rect 113548 439612 113600 439618
rect 113548 439554 113600 439560
rect 113364 438592 113416 438598
rect 113364 438534 113416 438540
rect 114468 438592 114520 438598
rect 114468 438534 114520 438540
rect 114480 438190 114508 438534
rect 114468 438184 114520 438190
rect 114468 438126 114520 438132
rect 112640 402946 112760 402974
rect 112536 391332 112588 391338
rect 112536 391274 112588 391280
rect 112168 388068 112220 388074
rect 112168 388010 112220 388016
rect 112444 388068 112496 388074
rect 112444 388010 112496 388016
rect 111798 387016 111854 387025
rect 111798 386951 111854 386960
rect 110616 386022 110920 386050
rect 107028 385886 107410 385914
rect 108698 385886 108988 385914
rect 109342 385886 109632 385914
rect 109986 385886 110368 385914
rect 110892 385914 110920 386022
rect 112180 385914 112208 388010
rect 110892 385886 111274 385914
rect 111918 385886 112208 385914
rect 105924 385750 106228 385778
rect 112732 385762 112760 402946
rect 114848 398886 114876 494974
rect 116044 494902 116072 583918
rect 117240 564398 117268 702714
rect 119344 630692 119396 630698
rect 119344 630634 119396 630640
rect 117412 588600 117464 588606
rect 117412 588542 117464 588548
rect 117320 581188 117372 581194
rect 117320 581130 117372 581136
rect 117228 564392 117280 564398
rect 117228 564334 117280 564340
rect 116124 560992 116176 560998
rect 116124 560934 116176 560940
rect 116136 496262 116164 560934
rect 116216 544400 116268 544406
rect 116216 544342 116268 544348
rect 116124 496256 116176 496262
rect 116124 496198 116176 496204
rect 116136 495514 116164 496198
rect 116124 495508 116176 495514
rect 116124 495450 116176 495456
rect 116032 494896 116084 494902
rect 116032 494838 116084 494844
rect 115112 491292 115164 491298
rect 115112 491234 115164 491240
rect 115124 491201 115152 491234
rect 115110 491192 115166 491201
rect 115110 491127 115166 491136
rect 115848 477556 115900 477562
rect 115848 477498 115900 477504
rect 115860 477465 115888 477498
rect 116032 477488 116084 477494
rect 115846 477456 115902 477465
rect 116032 477430 116084 477436
rect 115846 477391 115902 477400
rect 115204 466540 115256 466546
rect 115204 466482 115256 466488
rect 115848 466540 115900 466546
rect 115848 466482 115900 466488
rect 115110 400208 115166 400217
rect 115110 400143 115166 400152
rect 115124 398954 115152 400143
rect 115112 398948 115164 398954
rect 115112 398890 115164 398896
rect 114836 398880 114888 398886
rect 114836 398822 114888 398828
rect 114928 390788 114980 390794
rect 114928 390730 114980 390736
rect 114190 390688 114246 390697
rect 114190 390623 114246 390632
rect 114204 387977 114232 390623
rect 114284 390516 114336 390522
rect 114284 390458 114336 390464
rect 114296 389366 114324 390458
rect 114284 389360 114336 389366
rect 114284 389302 114336 389308
rect 114190 387968 114246 387977
rect 114190 387903 114246 387912
rect 114204 385914 114232 387903
rect 113850 385886 114232 385914
rect 114296 385778 114324 389302
rect 114940 389201 114968 390730
rect 114926 389192 114982 389201
rect 114926 389127 114982 389136
rect 114940 385778 114968 389127
rect 100668 385688 100720 385694
rect 100668 385630 100720 385636
rect 106200 385370 106228 385750
rect 112720 385756 112772 385762
rect 114296 385750 114494 385778
rect 114940 385750 115138 385778
rect 112720 385698 112772 385704
rect 112810 385384 112866 385393
rect 106200 385354 106320 385370
rect 77484 385348 77892 385354
rect 77536 385342 77892 385348
rect 90272 385348 90324 385354
rect 77484 385290 77536 385296
rect 90272 385290 90324 385296
rect 100024 385348 100076 385354
rect 106200 385348 106332 385354
rect 106200 385342 106280 385348
rect 100024 385290 100076 385296
rect 112562 385342 112810 385370
rect 112810 385319 112866 385328
rect 106280 385290 106332 385296
rect 69768 373966 70164 373994
rect 69664 371884 69716 371890
rect 69664 371826 69716 371832
rect 69768 367810 69796 373966
rect 69756 367804 69808 367810
rect 69756 367746 69808 367752
rect 69400 364306 69704 364334
rect 69676 340082 69704 364306
rect 115216 359530 115244 466482
rect 115860 466342 115888 466482
rect 115848 466336 115900 466342
rect 115848 466278 115900 466284
rect 116044 398138 116072 477430
rect 116228 452606 116256 544342
rect 116676 529236 116728 529242
rect 116676 529178 116728 529184
rect 116584 496188 116636 496194
rect 116584 496130 116636 496136
rect 116216 452600 116268 452606
rect 116216 452542 116268 452548
rect 116032 398132 116084 398138
rect 116032 398074 116084 398080
rect 115296 389904 115348 389910
rect 115296 389846 115348 389852
rect 115308 365106 115336 389846
rect 115756 389156 115808 389162
rect 115756 389098 115808 389104
rect 115768 387682 115796 389098
rect 115846 388376 115902 388385
rect 115846 388311 115902 388320
rect 115860 387870 115888 388311
rect 115848 387864 115900 387870
rect 115848 387806 115900 387812
rect 115768 387654 115888 387682
rect 115860 385914 115888 387654
rect 115782 385886 115888 385914
rect 115940 385008 115992 385014
rect 115940 384950 115992 384956
rect 115952 384033 115980 384950
rect 115938 384024 115994 384033
rect 115938 383959 115994 383968
rect 115308 365078 115428 365106
rect 115294 359544 115350 359553
rect 115216 359502 115294 359530
rect 115294 359479 115350 359488
rect 115400 357434 115428 365078
rect 115308 357406 115428 357434
rect 115308 349217 115336 357406
rect 115294 349208 115350 349217
rect 115294 349143 115350 349152
rect 70306 345944 70362 345953
rect 70306 345879 70362 345888
rect 69676 340068 70058 340082
rect 69676 340054 70072 340068
rect 70044 338094 70072 340054
rect 70320 338910 70348 345879
rect 70398 341728 70454 341737
rect 70398 341663 70454 341672
rect 70412 339998 70440 341663
rect 115756 341624 115808 341630
rect 115756 341566 115808 341572
rect 115768 340762 115796 341566
rect 115216 340748 115796 340762
rect 115216 340734 115782 340748
rect 70490 340232 70546 340241
rect 70490 340167 70546 340176
rect 70400 339992 70452 339998
rect 70400 339934 70452 339940
rect 70308 338904 70360 338910
rect 70308 338846 70360 338852
rect 70504 338842 70532 340167
rect 70492 338836 70544 338842
rect 70492 338778 70544 338784
rect 70688 338162 70716 340068
rect 71044 339992 71096 339998
rect 71044 339934 71096 339940
rect 70676 338156 70728 338162
rect 70676 338098 70728 338104
rect 70032 338088 70084 338094
rect 70032 338030 70084 338036
rect 70688 337550 70716 338098
rect 70676 337544 70728 337550
rect 70676 337486 70728 337492
rect 69204 319456 69256 319462
rect 69204 319398 69256 319404
rect 69112 313948 69164 313954
rect 69112 313890 69164 313896
rect 69020 313336 69072 313342
rect 69020 313278 69072 313284
rect 66904 303612 66956 303618
rect 66904 303554 66956 303560
rect 66168 302456 66220 302462
rect 66168 302398 66220 302404
rect 66180 302161 66208 302398
rect 66166 302152 66222 302161
rect 66166 302087 66222 302096
rect 65984 290488 66036 290494
rect 65984 290430 66036 290436
rect 65616 288380 65668 288386
rect 65616 288322 65668 288328
rect 65524 287428 65576 287434
rect 65524 287370 65576 287376
rect 65536 262886 65564 287370
rect 66076 271992 66128 271998
rect 66076 271934 66128 271940
rect 65524 262880 65576 262886
rect 65524 262822 65576 262828
rect 65984 255400 66036 255406
rect 65984 255342 66036 255348
rect 65892 244248 65944 244254
rect 65892 244190 65944 244196
rect 65904 238882 65932 244190
rect 65892 238876 65944 238882
rect 65892 238818 65944 238824
rect 65996 234054 66024 255342
rect 65984 234048 66036 234054
rect 65984 233990 66036 233996
rect 66088 229906 66116 271934
rect 66916 270881 66944 303554
rect 68926 299568 68982 299577
rect 68926 299503 68982 299512
rect 67548 298308 67600 298314
rect 67548 298250 67600 298256
rect 67560 287065 67588 298250
rect 67640 296948 67692 296954
rect 67640 296890 67692 296896
rect 67652 290873 67680 296890
rect 67730 291136 67786 291145
rect 67730 291071 67786 291080
rect 67638 290864 67694 290873
rect 67638 290799 67694 290808
rect 67744 290494 67772 291071
rect 67732 290488 67784 290494
rect 67732 290430 67784 290436
rect 67638 289232 67694 289241
rect 67638 289167 67694 289176
rect 67652 288454 67680 289167
rect 67640 288448 67692 288454
rect 67640 288390 67692 288396
rect 67824 288380 67876 288386
rect 67824 288322 67876 288328
rect 67836 288153 67864 288322
rect 67822 288144 67878 288153
rect 67822 288079 67878 288088
rect 67822 287464 67878 287473
rect 67822 287399 67824 287408
rect 67876 287399 67878 287408
rect 67824 287370 67876 287376
rect 67546 287056 67602 287065
rect 67546 286991 67602 287000
rect 68940 286113 68968 299503
rect 68926 286104 68982 286113
rect 68926 286039 68982 286048
rect 68282 284472 68338 284481
rect 68282 284407 68338 284416
rect 67640 284300 67692 284306
rect 67640 284242 67692 284248
rect 67652 283393 67680 284242
rect 67638 283384 67694 283393
rect 67638 283319 67694 283328
rect 67730 280528 67786 280537
rect 67730 280463 67786 280472
rect 67638 280392 67694 280401
rect 67638 280327 67694 280336
rect 67652 280226 67680 280327
rect 67744 280294 67772 280463
rect 67732 280288 67784 280294
rect 67732 280230 67784 280236
rect 67640 280220 67692 280226
rect 67640 280162 67692 280168
rect 68008 280152 68060 280158
rect 68008 280094 68060 280100
rect 67640 280084 67692 280090
rect 67640 280026 67692 280032
rect 67652 279313 67680 280026
rect 68020 279721 68048 280094
rect 68006 279712 68062 279721
rect 68006 279647 68062 279656
rect 67638 279304 67694 279313
rect 67638 279239 67694 279248
rect 67730 277808 67786 277817
rect 67730 277743 67786 277752
rect 67638 277672 67694 277681
rect 67638 277607 67694 277616
rect 67652 277506 67680 277607
rect 67640 277500 67692 277506
rect 67640 277442 67692 277448
rect 67744 277438 67772 277743
rect 67732 277432 67784 277438
rect 67732 277374 67784 277380
rect 67730 276448 67786 276457
rect 67730 276383 67786 276392
rect 67638 276312 67694 276321
rect 67638 276247 67694 276256
rect 67652 276146 67680 276247
rect 67640 276140 67692 276146
rect 67640 276082 67692 276088
rect 67744 276078 67772 276383
rect 67732 276072 67784 276078
rect 67732 276014 67784 276020
rect 67730 275224 67786 275233
rect 67730 275159 67786 275168
rect 67638 274952 67694 274961
rect 67638 274887 67694 274896
rect 67652 274718 67680 274887
rect 67744 274786 67772 275159
rect 67732 274780 67784 274786
rect 67732 274722 67784 274728
rect 67640 274712 67692 274718
rect 67640 274654 67692 274660
rect 68008 274644 68060 274650
rect 68008 274586 68060 274592
rect 68020 274281 68048 274586
rect 68006 274272 68062 274281
rect 68006 274207 68062 274216
rect 67638 273592 67694 273601
rect 67638 273527 67694 273536
rect 67652 273290 67680 273527
rect 67640 273284 67692 273290
rect 67640 273226 67692 273232
rect 67638 272368 67694 272377
rect 67638 272303 67694 272312
rect 67652 271930 67680 272303
rect 68190 272232 68246 272241
rect 68190 272167 68246 272176
rect 68204 271998 68232 272167
rect 68192 271992 68244 271998
rect 68192 271934 68244 271940
rect 67640 271924 67692 271930
rect 67640 271866 67692 271872
rect 67638 271008 67694 271017
rect 67638 270943 67694 270952
rect 66902 270872 66958 270881
rect 66902 270807 66958 270816
rect 67652 270570 67680 270943
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 68296 269822 68324 284407
rect 68926 283792 68982 283801
rect 68926 283727 68982 283736
rect 68284 269816 68336 269822
rect 68284 269758 68336 269764
rect 67730 269648 67786 269657
rect 67730 269583 67786 269592
rect 67638 269512 67694 269521
rect 67638 269447 67694 269456
rect 67652 269142 67680 269447
rect 67744 269210 67772 269583
rect 67732 269204 67784 269210
rect 67732 269146 67784 269152
rect 67640 269136 67692 269142
rect 67640 269078 67692 269084
rect 67730 268288 67786 268297
rect 67730 268223 67786 268232
rect 67638 268152 67694 268161
rect 67638 268087 67694 268096
rect 67652 267782 67680 268087
rect 67744 267850 67772 268223
rect 67732 267844 67784 267850
rect 67732 267786 67784 267792
rect 67640 267776 67692 267782
rect 67640 267718 67692 267724
rect 67638 267064 67694 267073
rect 67638 266999 67640 267008
rect 67692 266999 67694 267008
rect 67640 266970 67692 266976
rect 67640 266416 67692 266422
rect 67638 266384 67640 266393
rect 67692 266384 67694 266393
rect 67638 266319 67694 266328
rect 67824 266348 67876 266354
rect 67824 266290 67876 266296
rect 67730 265568 67786 265577
rect 67730 265503 67786 265512
rect 67744 264994 67772 265503
rect 67836 265441 67864 266290
rect 67822 265432 67878 265441
rect 67822 265367 67878 265376
rect 67732 264988 67784 264994
rect 67732 264930 67784 264936
rect 67640 264920 67692 264926
rect 67638 264888 67640 264897
rect 67692 264888 67694 264897
rect 67638 264823 67694 264832
rect 67638 263664 67694 263673
rect 67638 263599 67640 263608
rect 67692 263599 67694 263608
rect 67640 263570 67692 263576
rect 67730 262848 67786 262857
rect 67730 262783 67786 262792
rect 67744 262342 67772 262783
rect 67732 262336 67784 262342
rect 67638 262304 67694 262313
rect 67732 262278 67784 262284
rect 67638 262239 67640 262248
rect 67692 262239 67694 262248
rect 67640 262210 67692 262216
rect 67730 261488 67786 261497
rect 67730 261423 67786 261432
rect 66168 260976 66220 260982
rect 67640 260976 67692 260982
rect 66168 260918 66220 260924
rect 67638 260944 67640 260953
rect 67692 260944 67694 260953
rect 66076 229900 66128 229906
rect 66076 229842 66128 229848
rect 66180 178770 66208 260918
rect 67744 260914 67772 261423
rect 67638 260879 67694 260888
rect 67732 260908 67784 260914
rect 67732 260850 67784 260856
rect 67640 260840 67692 260846
rect 67638 260808 67640 260817
rect 67692 260808 67694 260817
rect 67638 260743 67694 260752
rect 67638 259584 67694 259593
rect 67638 259519 67694 259528
rect 67652 259486 67680 259519
rect 67640 259480 67692 259486
rect 67640 259422 67692 259428
rect 67730 258768 67786 258777
rect 67730 258703 67786 258712
rect 67638 258224 67694 258233
rect 67744 258194 67772 258703
rect 67638 258159 67694 258168
rect 67732 258188 67784 258194
rect 67652 258126 67680 258159
rect 67732 258130 67784 258136
rect 67640 258120 67692 258126
rect 67640 258062 67692 258068
rect 67916 258052 67968 258058
rect 67916 257994 67968 258000
rect 67928 257281 67956 257994
rect 67914 257272 67970 257281
rect 67914 257207 67970 257216
rect 67638 256864 67694 256873
rect 67638 256799 67694 256808
rect 67652 256766 67680 256799
rect 67640 256760 67692 256766
rect 67640 256702 67692 256708
rect 67638 255912 67694 255921
rect 67638 255847 67694 255856
rect 67652 255406 67680 255847
rect 67640 255400 67692 255406
rect 67640 255342 67692 255348
rect 67730 255368 67786 255377
rect 67730 255303 67732 255312
rect 67784 255303 67786 255312
rect 67732 255274 67784 255280
rect 67640 255264 67692 255270
rect 67638 255232 67640 255241
rect 67692 255232 67694 255241
rect 67638 255167 67694 255176
rect 67638 254008 67694 254017
rect 67638 253943 67640 253952
rect 67692 253943 67694 253952
rect 67640 253914 67692 253920
rect 67638 253192 67694 253201
rect 67638 253127 67694 253136
rect 67652 252618 67680 253127
rect 67640 252612 67692 252618
rect 67640 252554 67692 252560
rect 67730 251832 67786 251841
rect 67730 251767 67786 251776
rect 67638 251424 67694 251433
rect 67638 251359 67694 251368
rect 67652 251326 67680 251359
rect 67640 251320 67692 251326
rect 67640 251262 67692 251268
rect 67744 251258 67772 251767
rect 67732 251252 67784 251258
rect 67732 251194 67784 251200
rect 68650 250472 68706 250481
rect 68650 250407 68706 250416
rect 67638 249928 67694 249937
rect 67638 249863 67694 249872
rect 67652 249830 67680 249863
rect 67640 249824 67692 249830
rect 67640 249766 67692 249772
rect 67730 249112 67786 249121
rect 67730 249047 67786 249056
rect 67638 248568 67694 248577
rect 67744 248538 67772 249047
rect 67638 248503 67694 248512
rect 67732 248532 67784 248538
rect 67652 248470 67680 248503
rect 67732 248474 67784 248480
rect 67640 248464 67692 248470
rect 67640 248406 67692 248412
rect 67730 247752 67786 247761
rect 67730 247687 67786 247696
rect 67638 247208 67694 247217
rect 67638 247143 67640 247152
rect 67692 247143 67694 247152
rect 67640 247114 67692 247120
rect 67744 247110 67772 247687
rect 67732 247104 67784 247110
rect 67732 247046 67784 247052
rect 67730 246392 67786 246401
rect 67730 246327 67786 246336
rect 67638 245848 67694 245857
rect 67638 245783 67694 245792
rect 67652 245750 67680 245783
rect 67640 245744 67692 245750
rect 67640 245686 67692 245692
rect 67744 245682 67772 246327
rect 67732 245676 67784 245682
rect 67732 245618 67784 245624
rect 67454 244352 67510 244361
rect 67454 244287 67510 244296
rect 67468 238202 67496 244287
rect 67546 243672 67602 243681
rect 67546 243607 67602 243616
rect 67456 238196 67508 238202
rect 67456 238138 67508 238144
rect 67560 185638 67588 243607
rect 67638 243128 67694 243137
rect 67638 243063 67694 243072
rect 67652 243030 67680 243063
rect 67640 243024 67692 243030
rect 67640 242966 67692 242972
rect 67638 241904 67694 241913
rect 67638 241839 67694 241848
rect 67652 241534 67680 241839
rect 67640 241528 67692 241534
rect 67640 241470 67692 241476
rect 68664 239465 68692 250407
rect 68650 239456 68706 239465
rect 68650 239391 68706 239400
rect 68940 232665 68968 283727
rect 69032 282169 69060 313278
rect 70308 311228 70360 311234
rect 70308 311170 70360 311176
rect 70320 300150 70348 311170
rect 70398 302288 70454 302297
rect 70398 302223 70454 302232
rect 70308 300144 70360 300150
rect 70308 300086 70360 300092
rect 69112 295996 69164 296002
rect 69112 295938 69164 295944
rect 69124 286793 69152 295938
rect 69848 295452 69900 295458
rect 69848 295394 69900 295400
rect 69860 288833 69888 295394
rect 70032 295248 70084 295254
rect 70032 295190 70084 295196
rect 70044 291924 70072 295190
rect 70412 291977 70440 302223
rect 71056 301481 71084 339934
rect 71332 337958 71360 340068
rect 71780 338088 71832 338094
rect 71780 338030 71832 338036
rect 71320 337952 71372 337958
rect 71320 337894 71372 337900
rect 71332 336938 71360 337894
rect 71320 336932 71372 336938
rect 71320 336874 71372 336880
rect 71792 334626 71820 338030
rect 71976 336598 72004 340068
rect 73264 339590 73292 340068
rect 73252 339584 73304 339590
rect 73252 339526 73304 339532
rect 73264 337618 73292 339526
rect 73908 339386 73936 340068
rect 73896 339380 73948 339386
rect 73896 339322 73948 339328
rect 73908 338065 73936 339322
rect 73894 338056 73950 338065
rect 73894 337991 73950 338000
rect 74446 338056 74502 338065
rect 74446 337991 74502 338000
rect 73252 337612 73304 337618
rect 73252 337554 73304 337560
rect 71964 336592 72016 336598
rect 71964 336534 72016 336540
rect 71780 334620 71832 334626
rect 71780 334562 71832 334568
rect 71976 333266 72004 336534
rect 71964 333260 72016 333266
rect 71964 333202 72016 333208
rect 72424 325712 72476 325718
rect 72424 325654 72476 325660
rect 71136 312588 71188 312594
rect 71136 312530 71188 312536
rect 71042 301472 71098 301481
rect 71042 301407 71098 301416
rect 71148 292369 71176 312530
rect 71780 302252 71832 302258
rect 71780 302194 71832 302200
rect 71320 294432 71372 294438
rect 71320 294374 71372 294380
rect 71134 292360 71190 292369
rect 71134 292295 71190 292304
rect 70412 291949 70702 291977
rect 71332 291963 71360 294374
rect 71792 291977 71820 302194
rect 72436 294438 72464 325654
rect 74460 315353 74488 337991
rect 74552 337890 74580 340068
rect 74540 337884 74592 337890
rect 74540 337826 74592 337832
rect 75184 337884 75236 337890
rect 75184 337826 75236 337832
rect 75196 319530 75224 337826
rect 75840 335238 75868 340068
rect 75918 339688 75974 339697
rect 75918 339623 75974 339632
rect 75828 335232 75880 335238
rect 75828 335174 75880 335180
rect 75840 334150 75868 335174
rect 75276 334144 75328 334150
rect 75276 334086 75328 334092
rect 75828 334144 75880 334150
rect 75828 334086 75880 334092
rect 75184 319524 75236 319530
rect 75184 319466 75236 319472
rect 75288 318073 75316 334086
rect 75274 318064 75330 318073
rect 75274 317999 75330 318008
rect 74446 315344 74502 315353
rect 73160 315308 73212 315314
rect 74446 315279 74502 315288
rect 73160 315250 73212 315256
rect 72424 294432 72476 294438
rect 72424 294374 72476 294380
rect 73172 294370 73200 315250
rect 75184 309256 75236 309262
rect 75184 309198 75236 309204
rect 75196 306374 75224 309198
rect 75932 308514 75960 339623
rect 76484 338026 76512 340068
rect 77128 339697 77156 340068
rect 77114 339688 77170 339697
rect 77114 339623 77170 339632
rect 76472 338020 76524 338026
rect 76472 337962 76524 337968
rect 76484 331974 76512 337962
rect 78416 337754 78444 340068
rect 79076 339810 79104 340068
rect 79076 339782 79456 339810
rect 76564 337748 76616 337754
rect 76564 337690 76616 337696
rect 78404 337748 78456 337754
rect 78404 337690 78456 337696
rect 76576 335170 76604 337690
rect 76656 336932 76708 336938
rect 76656 336874 76708 336880
rect 76564 335164 76616 335170
rect 76564 335106 76616 335112
rect 76472 331968 76524 331974
rect 76472 331910 76524 331916
rect 76576 309874 76604 335106
rect 76668 323610 76696 336874
rect 79428 336818 79456 339782
rect 79152 336790 79456 336818
rect 79152 336666 79180 336790
rect 79324 336728 79376 336734
rect 79324 336670 79376 336676
rect 79140 336660 79192 336666
rect 79140 336602 79192 336608
rect 79336 336462 79364 336670
rect 79324 336456 79376 336462
rect 79324 336398 79376 336404
rect 77300 330540 77352 330546
rect 77300 330482 77352 330488
rect 76656 323604 76708 323610
rect 76656 323546 76708 323552
rect 76564 309868 76616 309874
rect 76564 309810 76616 309816
rect 75920 308508 75972 308514
rect 75920 308450 75972 308456
rect 75104 306346 75224 306374
rect 73250 300928 73306 300937
rect 73250 300863 73306 300872
rect 73160 294364 73212 294370
rect 73160 294306 73212 294312
rect 72608 294296 72660 294302
rect 72608 294238 72660 294244
rect 71792 291949 71990 291977
rect 72620 291963 72648 294238
rect 73264 291963 73292 300863
rect 74448 298784 74500 298790
rect 74448 298726 74500 298732
rect 73620 294364 73672 294370
rect 73620 294306 73672 294312
rect 73632 291977 73660 294306
rect 74460 294302 74488 298726
rect 74540 295520 74592 295526
rect 74540 295462 74592 295468
rect 74448 294296 74500 294302
rect 74448 294238 74500 294244
rect 73632 291949 73922 291977
rect 74552 291963 74580 295462
rect 75104 295254 75132 306346
rect 75920 302320 75972 302326
rect 75920 302262 75972 302268
rect 75184 296812 75236 296818
rect 75184 296754 75236 296760
rect 75092 295248 75144 295254
rect 75092 295190 75144 295196
rect 75196 291963 75224 296754
rect 75826 294128 75882 294137
rect 75826 294063 75882 294072
rect 75840 291963 75868 294063
rect 75932 291977 75960 302262
rect 77312 294370 77340 330482
rect 79336 311370 79364 336398
rect 79428 316713 79456 336790
rect 79704 336734 79732 340068
rect 80946 339810 80974 340068
rect 80716 339782 80974 339810
rect 79692 336728 79744 336734
rect 79692 336670 79744 336676
rect 80716 333946 80744 339782
rect 81636 339522 81664 340068
rect 81624 339516 81676 339522
rect 81624 339458 81676 339464
rect 81636 337414 81664 339458
rect 81624 337408 81676 337414
rect 81624 337350 81676 337356
rect 80704 333940 80756 333946
rect 80704 333882 80756 333888
rect 80716 325038 80744 333882
rect 82280 332042 82308 340068
rect 83522 339810 83550 340068
rect 83476 339782 83550 339810
rect 83476 336666 83504 339782
rect 84212 337482 84240 340068
rect 84200 337476 84252 337482
rect 84200 337418 84252 337424
rect 83464 336660 83516 336666
rect 83464 336602 83516 336608
rect 82268 332036 82320 332042
rect 82268 331978 82320 331984
rect 80704 325032 80756 325038
rect 80704 324974 80756 324980
rect 83476 318102 83504 336602
rect 84856 336054 84884 340068
rect 86160 339810 86188 340068
rect 86160 339782 86264 339810
rect 86236 339454 86264 339782
rect 86224 339448 86276 339454
rect 86224 339390 86276 339396
rect 84844 336048 84896 336054
rect 84844 335990 84896 335996
rect 86236 322318 86264 339390
rect 86788 339318 86816 340068
rect 86776 339312 86828 339318
rect 86776 339254 86828 339260
rect 86788 338026 86816 339254
rect 87432 338094 87460 340068
rect 88736 339810 88764 340068
rect 88736 339782 89024 339810
rect 87420 338088 87472 338094
rect 87420 338030 87472 338036
rect 86776 338020 86828 338026
rect 86776 337962 86828 337968
rect 87604 338020 87656 338026
rect 87604 337962 87656 337968
rect 86224 322312 86276 322318
rect 86224 322254 86276 322260
rect 83464 318096 83516 318102
rect 83464 318038 83516 318044
rect 84292 316736 84344 316742
rect 79414 316704 79470 316713
rect 84292 316678 84344 316684
rect 79414 316639 79470 316648
rect 81440 311908 81492 311914
rect 81440 311850 81492 311856
rect 79324 311364 79376 311370
rect 79324 311306 79376 311312
rect 80060 309936 80112 309942
rect 80060 309878 80112 309884
rect 77392 304972 77444 304978
rect 77392 304914 77444 304920
rect 77300 294364 77352 294370
rect 77300 294306 77352 294312
rect 77116 293344 77168 293350
rect 77116 293286 77168 293292
rect 75932 291949 76498 291977
rect 77128 291963 77156 293286
rect 77404 291977 77432 304914
rect 79324 301028 79376 301034
rect 79324 300970 79376 300976
rect 78036 294364 78088 294370
rect 78036 294306 78088 294312
rect 77404 291949 77786 291977
rect 78048 291938 78076 294306
rect 79048 294092 79100 294098
rect 79048 294034 79100 294040
rect 79060 291963 79088 294034
rect 79336 291938 79364 300970
rect 80072 291977 80100 309878
rect 80980 294092 81032 294098
rect 80980 294034 81032 294040
rect 80072 291949 80362 291977
rect 80992 291963 81020 294034
rect 81452 291977 81480 311850
rect 81900 305108 81952 305114
rect 81900 305050 81952 305056
rect 81452 291949 81650 291977
rect 81912 291938 81940 305050
rect 83556 298444 83608 298450
rect 83556 298386 83608 298392
rect 82912 296880 82964 296886
rect 82912 296822 82964 296828
rect 82924 291963 82952 296822
rect 83568 291963 83596 298386
rect 84200 294704 84252 294710
rect 84200 294646 84252 294652
rect 84212 291963 84240 294646
rect 84304 294370 84332 316678
rect 84384 308440 84436 308446
rect 84384 308382 84436 308388
rect 84292 294364 84344 294370
rect 84292 294306 84344 294312
rect 84396 291938 84424 308382
rect 86960 306536 87012 306542
rect 86960 306478 87012 306484
rect 85580 306468 85632 306474
rect 85580 306410 85632 306416
rect 85212 294364 85264 294370
rect 85212 294306 85264 294312
rect 85224 291977 85252 294306
rect 85224 291949 85514 291977
rect 85592 291938 85620 306410
rect 86316 303748 86368 303754
rect 86316 303690 86368 303696
rect 86328 291977 86356 303690
rect 86328 291949 86802 291977
rect 86972 291938 87000 306478
rect 87616 300150 87644 337962
rect 88996 336530 89024 339782
rect 88984 336524 89036 336530
rect 88984 336466 89036 336472
rect 88996 322250 89024 336466
rect 89364 328438 89392 340068
rect 90008 339250 90036 340068
rect 89996 339244 90048 339250
rect 89996 339186 90048 339192
rect 90364 339244 90416 339250
rect 90364 339186 90416 339192
rect 89352 328432 89404 328438
rect 89352 328374 89404 328380
rect 88984 322244 89036 322250
rect 88984 322186 89036 322192
rect 89720 309188 89772 309194
rect 89720 309130 89772 309136
rect 88340 300960 88392 300966
rect 88340 300902 88392 300908
rect 87604 300144 87656 300150
rect 87604 300086 87656 300092
rect 88064 295588 88116 295594
rect 88064 295530 88116 295536
rect 88076 291963 88104 295530
rect 88352 294370 88380 300902
rect 88432 300892 88484 300898
rect 88432 300834 88484 300840
rect 88340 294364 88392 294370
rect 88340 294306 88392 294312
rect 88444 291977 88472 300834
rect 89076 294364 89128 294370
rect 89076 294306 89128 294312
rect 89088 291977 89116 294306
rect 89732 291977 89760 309130
rect 90376 305726 90404 339186
rect 91296 337754 91324 340068
rect 91284 337748 91336 337754
rect 91284 337690 91336 337696
rect 91008 337612 91060 337618
rect 91008 337554 91060 337560
rect 91020 333305 91048 337554
rect 91006 333296 91062 333305
rect 91006 333231 91062 333240
rect 91940 315994 91968 340068
rect 92584 333878 92612 340068
rect 92572 333872 92624 333878
rect 92572 333814 92624 333820
rect 92584 332654 92612 333814
rect 92572 332648 92624 332654
rect 92572 332590 92624 332596
rect 93124 332648 93176 332654
rect 93124 332590 93176 332596
rect 91928 315988 91980 315994
rect 91928 315930 91980 315936
rect 91100 311296 91152 311302
rect 91100 311238 91152 311244
rect 91112 309942 91140 311238
rect 91100 309936 91152 309942
rect 91100 309878 91152 309884
rect 90364 305720 90416 305726
rect 90364 305662 90416 305668
rect 93136 305658 93164 332590
rect 93228 329730 93256 340068
rect 93676 337748 93728 337754
rect 93676 337690 93728 337696
rect 93308 337544 93360 337550
rect 93308 337486 93360 337492
rect 93216 329724 93268 329730
rect 93216 329666 93268 329672
rect 93320 323678 93348 337486
rect 93688 335238 93716 337690
rect 93676 335232 93728 335238
rect 93676 335174 93728 335180
rect 93308 323672 93360 323678
rect 93308 323614 93360 323620
rect 93688 307086 93716 335174
rect 94516 334762 94544 340068
rect 95114 339810 95142 340068
rect 95068 339782 95142 339810
rect 94504 334756 94556 334762
rect 94504 334698 94556 334704
rect 95068 333946 95096 339782
rect 95804 337890 95832 340068
rect 96712 338088 96764 338094
rect 96712 338030 96764 338036
rect 95792 337884 95844 337890
rect 95792 337826 95844 337832
rect 95056 333940 95108 333946
rect 95056 333882 95108 333888
rect 93768 329112 93820 329118
rect 93768 329054 93820 329060
rect 93676 307080 93728 307086
rect 93676 307022 93728 307028
rect 93124 305652 93176 305658
rect 93124 305594 93176 305600
rect 90272 302524 90324 302530
rect 90272 302466 90324 302472
rect 90284 291977 90312 302466
rect 93216 298240 93268 298246
rect 93216 298182 93268 298188
rect 91928 297084 91980 297090
rect 91928 297026 91980 297032
rect 91282 294536 91338 294545
rect 91282 294471 91338 294480
rect 88444 291949 88734 291977
rect 89088 291949 89378 291977
rect 89732 291949 90022 291977
rect 90284 291949 90666 291977
rect 91296 291963 91324 294471
rect 91940 291963 91968 297026
rect 92572 295724 92624 295730
rect 92572 295666 92624 295672
rect 92584 291963 92612 295666
rect 93228 291963 93256 298182
rect 93780 295730 93808 329054
rect 95068 303822 95096 333882
rect 95148 332036 95200 332042
rect 95148 331978 95200 331984
rect 94504 303816 94556 303822
rect 94504 303758 94556 303764
rect 95056 303816 95108 303822
rect 95056 303758 95108 303764
rect 93952 302932 94004 302938
rect 93952 302874 94004 302880
rect 93768 295724 93820 295730
rect 93768 295666 93820 295672
rect 93964 294370 93992 302874
rect 94044 300076 94096 300082
rect 94044 300018 94096 300024
rect 93952 294364 94004 294370
rect 93952 294306 94004 294312
rect 93860 292732 93912 292738
rect 93860 292674 93912 292680
rect 93872 291963 93900 292674
rect 94056 291977 94084 300018
rect 94516 296002 94544 303758
rect 95160 300082 95188 331978
rect 96620 303816 96672 303822
rect 96620 303758 96672 303764
rect 95148 300076 95200 300082
rect 95148 300018 95200 300024
rect 95160 299674 95188 300018
rect 95148 299668 95200 299674
rect 95148 299610 95200 299616
rect 94504 295996 94556 296002
rect 94504 295938 94556 295944
rect 96632 294386 96660 303758
rect 96724 296041 96752 338030
rect 97092 337074 97120 340068
rect 97080 337068 97132 337074
rect 97080 337010 97132 337016
rect 97736 328370 97764 340068
rect 97908 338768 97960 338774
rect 97908 338710 97960 338716
rect 97920 338094 97948 338710
rect 97908 338088 97960 338094
rect 97908 338030 97960 338036
rect 98380 335306 98408 340068
rect 98644 338904 98696 338910
rect 98644 338846 98696 338852
rect 98368 335300 98420 335306
rect 98368 335242 98420 335248
rect 97724 328364 97776 328370
rect 97724 328306 97776 328312
rect 98656 297022 98684 338846
rect 99668 337482 99696 340068
rect 100312 337958 100340 340068
rect 100300 337952 100352 337958
rect 100300 337894 100352 337900
rect 99656 337476 99708 337482
rect 99656 337418 99708 337424
rect 100024 337068 100076 337074
rect 100024 337010 100076 337016
rect 100036 320142 100064 337010
rect 100956 329798 100984 340068
rect 102138 338192 102194 338201
rect 102138 338127 102194 338136
rect 102152 338094 102180 338127
rect 102140 338088 102192 338094
rect 102140 338030 102192 338036
rect 102048 337476 102100 337482
rect 102048 337418 102100 337424
rect 100944 329792 100996 329798
rect 100944 329734 100996 329740
rect 100024 320136 100076 320142
rect 100024 320078 100076 320084
rect 102060 307834 102088 337418
rect 102244 313274 102272 340068
rect 102232 313268 102284 313274
rect 102232 313210 102284 313216
rect 102888 311846 102916 340068
rect 103532 335306 103560 340068
rect 104820 336666 104848 340068
rect 104164 336660 104216 336666
rect 104164 336602 104216 336608
rect 104808 336660 104860 336666
rect 104808 336602 104860 336608
rect 103520 335300 103572 335306
rect 103520 335242 103572 335248
rect 102876 311840 102928 311846
rect 102876 311782 102928 311788
rect 104176 311234 104204 336602
rect 105464 321570 105492 340068
rect 106108 336734 106136 340068
rect 107396 339454 107424 340068
rect 107994 339810 108022 340068
rect 107948 339782 108022 339810
rect 107948 339590 107976 339782
rect 107936 339584 107988 339590
rect 107936 339526 107988 339532
rect 107384 339448 107436 339454
rect 107384 339390 107436 339396
rect 107568 339448 107620 339454
rect 107568 339390 107620 339396
rect 106096 336728 106148 336734
rect 106096 336670 106148 336676
rect 105452 321564 105504 321570
rect 105452 321506 105504 321512
rect 106108 318170 106136 336670
rect 106188 325100 106240 325106
rect 106188 325042 106240 325048
rect 106096 318164 106148 318170
rect 106096 318106 106148 318112
rect 104164 311228 104216 311234
rect 104164 311170 104216 311176
rect 102048 307828 102100 307834
rect 102048 307770 102100 307776
rect 103704 307828 103756 307834
rect 103704 307770 103756 307776
rect 103716 306374 103744 307770
rect 103716 306346 104296 306374
rect 102876 298172 102928 298178
rect 102876 298114 102928 298120
rect 101586 297392 101642 297401
rect 101586 297327 101642 297336
rect 98644 297016 98696 297022
rect 98644 296958 98696 296964
rect 96710 296032 96766 296041
rect 96710 295967 96766 295976
rect 94780 294364 94832 294370
rect 96632 294358 97212 294386
rect 94780 294306 94832 294312
rect 94056 291949 94530 291977
rect 94792 291938 94820 294306
rect 95790 294264 95846 294273
rect 95790 294199 95846 294208
rect 95804 291963 95832 294199
rect 96436 294024 96488 294030
rect 96436 293966 96488 293972
rect 96448 291963 96476 293966
rect 97080 293276 97132 293282
rect 97080 293218 97132 293224
rect 97092 292641 97120 293218
rect 97078 292632 97134 292641
rect 97078 292567 97134 292576
rect 97092 291963 97120 292567
rect 97184 291938 97212 294358
rect 98656 291977 98684 296958
rect 99656 295656 99708 295662
rect 99656 295598 99708 295604
rect 99012 294772 99064 294778
rect 99012 294714 99064 294720
rect 98394 291949 98684 291977
rect 99024 291963 99052 294714
rect 99668 291963 99696 295598
rect 100942 295488 100998 295497
rect 100942 295423 100998 295432
rect 100956 291963 100984 295423
rect 101600 291963 101628 297327
rect 102232 292596 102284 292602
rect 102232 292538 102284 292544
rect 102244 291963 102272 292538
rect 102888 291963 102916 298114
rect 103520 294228 103572 294234
rect 103520 294170 103572 294176
rect 103532 291963 103560 294170
rect 104268 291977 104296 306346
rect 105636 301572 105688 301578
rect 105636 301514 105688 301520
rect 104900 301436 104952 301442
rect 104900 301378 104952 301384
rect 104268 291949 104834 291977
rect 104912 291938 104940 301378
rect 105648 291977 105676 301514
rect 106200 301442 106228 325042
rect 106280 306400 106332 306406
rect 106332 306348 106872 306374
rect 106280 306346 106872 306348
rect 106280 306342 106332 306346
rect 106188 301436 106240 301442
rect 106188 301378 106240 301384
rect 106200 301102 106228 301378
rect 106188 301096 106240 301102
rect 106188 301038 106240 301044
rect 106740 295384 106792 295390
rect 106740 295326 106792 295332
rect 105648 291949 106122 291977
rect 106752 291963 106780 295326
rect 106844 291977 106872 306346
rect 107580 304366 107608 339390
rect 107948 335354 107976 339526
rect 107672 335326 107976 335354
rect 107672 324970 107700 335326
rect 108304 325712 108356 325718
rect 108684 325694 108712 340068
rect 109972 339425 110000 340068
rect 109958 339416 110014 339425
rect 109958 339351 110014 339360
rect 109972 338094 110000 339351
rect 109960 338088 110012 338094
rect 109960 338030 110012 338036
rect 110616 327078 110644 340068
rect 110604 327072 110656 327078
rect 110604 327014 110656 327020
rect 108356 325666 108712 325694
rect 108304 325654 108356 325660
rect 107660 324964 107712 324970
rect 107660 324906 107712 324912
rect 107660 309936 107712 309942
rect 107660 309878 107712 309884
rect 107672 306374 107700 309878
rect 108316 309126 108344 325654
rect 111260 325650 111288 340068
rect 112444 338904 112496 338910
rect 112444 338846 112496 338852
rect 111248 325644 111300 325650
rect 111248 325586 111300 325592
rect 112456 320890 112484 338846
rect 112548 338094 112576 340068
rect 113088 338972 113140 338978
rect 113088 338914 113140 338920
rect 112536 338088 112588 338094
rect 112536 338030 112588 338036
rect 112444 320884 112496 320890
rect 112444 320826 112496 320832
rect 108304 309120 108356 309126
rect 108304 309062 108356 309068
rect 107672 306346 108344 306374
rect 107568 304360 107620 304366
rect 107568 304302 107620 304308
rect 108026 293992 108082 294001
rect 108026 293927 108082 293936
rect 106844 291949 107410 291977
rect 108040 291963 108068 293927
rect 108316 291977 108344 306346
rect 110420 299600 110472 299606
rect 110420 299542 110472 299548
rect 109040 299532 109092 299538
rect 109040 299474 109092 299480
rect 109052 291977 109080 299474
rect 109960 294636 110012 294642
rect 109960 294578 110012 294584
rect 108316 291949 108698 291977
rect 109052 291949 109342 291977
rect 109972 291963 110000 294578
rect 110432 291977 110460 299542
rect 111246 295352 111302 295361
rect 111246 295287 111302 295296
rect 110432 291949 110630 291977
rect 111260 291963 111288 295287
rect 113100 293418 113128 338914
rect 113192 332110 113220 340068
rect 113836 339522 113864 340068
rect 113272 339516 113324 339522
rect 113272 339458 113324 339464
rect 113824 339516 113876 339522
rect 113824 339458 113876 339464
rect 113180 332104 113232 332110
rect 113180 332046 113232 332052
rect 113284 332042 113312 339458
rect 115124 338026 115152 340068
rect 115112 338020 115164 338026
rect 115112 337962 115164 337968
rect 113916 332580 113968 332586
rect 113916 332522 113968 332528
rect 113928 332110 113956 332522
rect 113916 332104 113968 332110
rect 113916 332046 113968 332052
rect 113272 332036 113324 332042
rect 113272 331978 113324 331984
rect 113824 318164 113876 318170
rect 113824 318106 113876 318112
rect 113178 296848 113234 296857
rect 113178 296783 113234 296792
rect 113192 294778 113220 296783
rect 113836 296750 113864 318106
rect 113928 316742 113956 332046
rect 115124 329118 115152 337962
rect 115112 329112 115164 329118
rect 115112 329054 115164 329060
rect 115216 316742 115244 340734
rect 115296 326392 115348 326398
rect 115296 326334 115348 326340
rect 113916 316736 113968 316742
rect 113916 316678 113968 316684
rect 115204 316736 115256 316742
rect 115204 316678 115256 316684
rect 114468 311160 114520 311166
rect 114468 311102 114520 311108
rect 114480 308446 114508 311102
rect 114468 308440 114520 308446
rect 114468 308382 114520 308388
rect 113916 299736 113968 299742
rect 113916 299678 113968 299684
rect 113456 296744 113508 296750
rect 113456 296686 113508 296692
rect 113824 296744 113876 296750
rect 113824 296686 113876 296692
rect 113180 294772 113232 294778
rect 113180 294714 113232 294720
rect 113088 293412 113140 293418
rect 113088 293354 113140 293360
rect 111890 292768 111946 292777
rect 111890 292703 111946 292712
rect 111904 291963 111932 292703
rect 112536 292664 112588 292670
rect 112536 292606 112588 292612
rect 112548 291963 112576 292606
rect 113468 291977 113496 296686
rect 113928 294710 113956 299678
rect 113916 294704 113968 294710
rect 113916 294646 113968 294652
rect 115112 294296 115164 294302
rect 115112 294238 115164 294244
rect 113824 294024 113876 294030
rect 113824 293966 113876 293972
rect 113206 291949 113496 291977
rect 113836 291963 113864 293966
rect 115124 291963 115152 294238
rect 115308 294166 115336 326334
rect 115952 325106 115980 383959
rect 116044 370433 116072 398074
rect 116596 396030 116624 496130
rect 116688 459610 116716 529178
rect 117332 488442 117360 581130
rect 117424 536790 117452 588542
rect 118792 585268 118844 585274
rect 118792 585210 118844 585216
rect 117964 567248 118016 567254
rect 117964 567190 118016 567196
rect 117412 536784 117464 536790
rect 117412 536726 117464 536732
rect 117424 535498 117452 536726
rect 117412 535492 117464 535498
rect 117412 535434 117464 535440
rect 117504 497684 117556 497690
rect 117504 497626 117556 497632
rect 117412 489184 117464 489190
rect 117410 489152 117412 489161
rect 117464 489152 117466 489161
rect 117410 489087 117466 489096
rect 117320 488436 117372 488442
rect 117320 488378 117372 488384
rect 117044 481704 117096 481710
rect 117044 481646 117096 481652
rect 117056 481545 117084 481646
rect 117042 481536 117098 481545
rect 117042 481471 117098 481480
rect 117320 479528 117372 479534
rect 117320 479470 117372 479476
rect 116676 459604 116728 459610
rect 116676 459546 116728 459552
rect 116688 459474 116716 459546
rect 116676 459468 116728 459474
rect 116676 459410 116728 459416
rect 116584 396024 116636 396030
rect 116584 395966 116636 395972
rect 116124 394120 116176 394126
rect 116124 394062 116176 394068
rect 116030 370424 116086 370433
rect 116030 370359 116086 370368
rect 116032 369912 116084 369918
rect 116032 369854 116084 369860
rect 115940 325100 115992 325106
rect 115940 325042 115992 325048
rect 115388 319524 115440 319530
rect 115388 319466 115440 319472
rect 115400 294302 115428 319466
rect 116044 315314 116072 369854
rect 116136 357105 116164 394062
rect 116214 391232 116270 391241
rect 116214 391167 116270 391176
rect 116228 371385 116256 391167
rect 117332 379545 117360 479470
rect 117516 440910 117544 497626
rect 117686 477456 117742 477465
rect 117686 477391 117742 477400
rect 117504 440904 117556 440910
rect 117504 440846 117556 440852
rect 117504 399560 117556 399566
rect 117504 399502 117556 399508
rect 117412 385756 117464 385762
rect 117412 385698 117464 385704
rect 117318 379536 117374 379545
rect 117318 379471 117374 379480
rect 116214 371376 116270 371385
rect 116214 371311 116270 371320
rect 116214 370696 116270 370705
rect 116214 370631 116270 370640
rect 116228 369918 116256 370631
rect 116216 369912 116268 369918
rect 116216 369854 116268 369860
rect 117320 369164 117372 369170
rect 117320 369106 117372 369112
rect 117332 368665 117360 369106
rect 117318 368656 117374 368665
rect 117424 368626 117452 385698
rect 117318 368591 117374 368600
rect 117412 368620 117464 368626
rect 117412 368562 117464 368568
rect 117412 368484 117464 368490
rect 117412 368426 117464 368432
rect 117320 368416 117372 368422
rect 117320 368358 117372 368364
rect 117332 367985 117360 368358
rect 117318 367976 117374 367985
rect 117318 367911 117374 367920
rect 117424 367305 117452 368426
rect 117410 367296 117466 367305
rect 117410 367231 117466 367240
rect 117320 367056 117372 367062
rect 117320 366998 117372 367004
rect 117332 365945 117360 366998
rect 117318 365936 117374 365945
rect 117318 365871 117374 365880
rect 117318 365256 117374 365265
rect 117318 365191 117374 365200
rect 117332 364886 117360 365191
rect 117320 364880 117372 364886
rect 117320 364822 117372 364828
rect 117320 362908 117372 362914
rect 117320 362850 117372 362856
rect 117332 362545 117360 362850
rect 117318 362536 117374 362545
rect 117318 362471 117374 362480
rect 117320 362228 117372 362234
rect 117320 362170 117372 362176
rect 117332 361865 117360 362170
rect 117318 361856 117374 361865
rect 117318 361791 117374 361800
rect 117318 361176 117374 361185
rect 117318 361111 117374 361120
rect 117332 360262 117360 361111
rect 117320 360256 117372 360262
rect 117320 360198 117372 360204
rect 116122 357096 116178 357105
rect 116122 357031 116178 357040
rect 117516 351665 117544 399502
rect 117596 394188 117648 394194
rect 117596 394130 117648 394136
rect 117608 355745 117636 394130
rect 117700 386345 117728 477391
rect 117976 476134 118004 567190
rect 118700 535492 118752 535498
rect 118700 535434 118752 535440
rect 117964 476128 118016 476134
rect 117964 476070 118016 476076
rect 117976 475930 118004 476070
rect 117964 475924 118016 475930
rect 117964 475866 118016 475872
rect 118712 437374 118740 535434
rect 118804 494834 118832 585210
rect 118884 576156 118936 576162
rect 118884 576098 118936 576104
rect 118792 494828 118844 494834
rect 118792 494770 118844 494776
rect 118896 491298 118924 576098
rect 119356 538150 119384 630634
rect 136652 592686 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700398 154160 703520
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 162124 700392 162176 700398
rect 162124 700334 162176 700340
rect 159364 683188 159416 683194
rect 159364 683130 159416 683136
rect 136640 592680 136692 592686
rect 136640 592622 136692 592628
rect 131304 586764 131356 586770
rect 131304 586706 131356 586712
rect 123024 586628 123076 586634
rect 123024 586570 123076 586576
rect 120080 585336 120132 585342
rect 120080 585278 120132 585284
rect 119436 555484 119488 555490
rect 119436 555426 119488 555432
rect 119344 538144 119396 538150
rect 119344 538086 119396 538092
rect 118884 491292 118936 491298
rect 118884 491234 118936 491240
rect 118792 489864 118844 489870
rect 118792 489806 118844 489812
rect 118804 488617 118832 489806
rect 118790 488608 118846 488617
rect 118790 488543 118846 488552
rect 118792 487552 118844 487558
rect 118792 487494 118844 487500
rect 118700 437368 118752 437374
rect 118700 437310 118752 437316
rect 118804 422278 118832 487494
rect 118884 472728 118936 472734
rect 118884 472670 118936 472676
rect 118896 471374 118924 472670
rect 118884 471368 118936 471374
rect 118884 471310 118936 471316
rect 119448 463690 119476 555426
rect 120092 493406 120120 585278
rect 121550 583808 121606 583817
rect 121550 583743 121606 583752
rect 121460 583024 121512 583030
rect 121460 582966 121512 582972
rect 120172 582548 120224 582554
rect 120172 582490 120224 582496
rect 120184 497622 120212 582490
rect 120172 497616 120224 497622
rect 120172 497558 120224 497564
rect 120264 497548 120316 497554
rect 120264 497490 120316 497496
rect 120080 493400 120132 493406
rect 120080 493342 120132 493348
rect 120080 492720 120132 492726
rect 120080 492662 120132 492668
rect 119988 466404 120040 466410
rect 119988 466346 120040 466352
rect 119436 463684 119488 463690
rect 119436 463626 119488 463632
rect 118792 422272 118844 422278
rect 118792 422214 118844 422220
rect 118804 420986 118832 422214
rect 118792 420980 118844 420986
rect 118792 420922 118844 420928
rect 119344 420980 119396 420986
rect 119344 420922 119396 420928
rect 119356 389366 119384 420922
rect 118792 389360 118844 389366
rect 118792 389302 118844 389308
rect 119344 389360 119396 389366
rect 119344 389302 119396 389308
rect 118700 387116 118752 387122
rect 118700 387058 118752 387064
rect 117686 386336 117742 386345
rect 117686 386271 117742 386280
rect 118514 384976 118570 384985
rect 118514 384911 118570 384920
rect 118528 383722 118556 384911
rect 118516 383716 118568 383722
rect 118516 383658 118568 383664
rect 118608 383648 118660 383654
rect 118606 383616 118608 383625
rect 118660 383616 118662 383625
rect 118606 383551 118662 383560
rect 118606 381576 118662 381585
rect 118606 381511 118608 381520
rect 118660 381511 118662 381520
rect 118608 381482 118660 381488
rect 118606 380896 118662 380905
rect 118606 380831 118608 380840
rect 118660 380831 118662 380840
rect 118608 380802 118660 380808
rect 118332 380180 118384 380186
rect 118332 380122 118384 380128
rect 118344 379545 118372 380122
rect 118330 379536 118386 379545
rect 118330 379471 118386 379480
rect 118608 378888 118660 378894
rect 118606 378856 118608 378865
rect 118660 378856 118662 378865
rect 118606 378791 118662 378800
rect 118608 378208 118660 378214
rect 118606 378176 118608 378185
rect 118660 378176 118662 378185
rect 118606 378111 118662 378120
rect 118422 376816 118478 376825
rect 118422 376751 118424 376760
rect 118476 376751 118478 376760
rect 118424 376722 118476 376728
rect 118608 376712 118660 376718
rect 118608 376654 118660 376660
rect 117780 376304 117832 376310
rect 117780 376246 117832 376252
rect 117792 376145 117820 376246
rect 117778 376136 117834 376145
rect 117778 376071 117834 376080
rect 118620 375465 118648 376654
rect 118606 375456 118662 375465
rect 118606 375391 118662 375400
rect 118608 375352 118660 375358
rect 118608 375294 118660 375300
rect 118620 374105 118648 375294
rect 118606 374096 118662 374105
rect 118606 374031 118662 374040
rect 118608 373992 118660 373998
rect 118608 373934 118660 373940
rect 118620 373425 118648 373934
rect 118606 373416 118662 373425
rect 118606 373351 118662 373360
rect 117870 370696 117926 370705
rect 117870 370631 117926 370640
rect 117884 370530 117912 370631
rect 117872 370524 117924 370530
rect 117872 370466 117924 370472
rect 118054 370016 118110 370025
rect 118054 369951 118110 369960
rect 118068 369918 118096 369951
rect 118056 369912 118108 369918
rect 118056 369854 118108 369860
rect 117688 368620 117740 368626
rect 117688 368562 117740 368568
rect 117700 363662 117728 368562
rect 117688 363656 117740 363662
rect 117688 363598 117740 363604
rect 117700 363225 117728 363598
rect 117686 363216 117742 363225
rect 117686 363151 117742 363160
rect 117870 359136 117926 359145
rect 117870 359071 117926 359080
rect 117884 358834 117912 359071
rect 117872 358828 117924 358834
rect 117872 358770 117924 358776
rect 118606 358456 118662 358465
rect 118606 358391 118662 358400
rect 118620 358086 118648 358391
rect 118608 358080 118660 358086
rect 118608 358022 118660 358028
rect 118146 357096 118202 357105
rect 118146 357031 118202 357040
rect 118160 356114 118188 357031
rect 118606 356416 118662 356425
rect 118606 356351 118662 356360
rect 118620 356182 118648 356351
rect 118608 356176 118660 356182
rect 118608 356118 118660 356124
rect 118148 356108 118200 356114
rect 118148 356050 118200 356056
rect 117594 355736 117650 355745
rect 117594 355671 117650 355680
rect 118606 355736 118662 355745
rect 118606 355671 118662 355680
rect 118620 355366 118648 355671
rect 118608 355360 118660 355366
rect 118608 355302 118660 355308
rect 118516 354680 118568 354686
rect 118516 354622 118568 354628
rect 118528 353705 118556 354622
rect 118606 354376 118662 354385
rect 118606 354311 118662 354320
rect 118620 354074 118648 354311
rect 118608 354068 118660 354074
rect 118608 354010 118660 354016
rect 118514 353696 118570 353705
rect 118514 353631 118570 353640
rect 118606 353016 118662 353025
rect 118606 352951 118662 352960
rect 118620 352578 118648 352951
rect 118608 352572 118660 352578
rect 118608 352514 118660 352520
rect 118056 351892 118108 351898
rect 118056 351834 118108 351840
rect 117502 351656 117558 351665
rect 117502 351591 117558 351600
rect 118068 350985 118096 351834
rect 118606 351656 118662 351665
rect 118606 351591 118662 351600
rect 118620 351286 118648 351591
rect 118608 351280 118660 351286
rect 118608 351222 118660 351228
rect 118054 350976 118110 350985
rect 118054 350911 118110 350920
rect 118606 350296 118662 350305
rect 118606 350231 118662 350240
rect 118620 349858 118648 350231
rect 118608 349852 118660 349858
rect 118608 349794 118660 349800
rect 118608 349104 118660 349110
rect 118608 349046 118660 349052
rect 117870 348936 117926 348945
rect 117870 348871 117926 348880
rect 117884 347818 117912 348871
rect 118620 348265 118648 349046
rect 118606 348256 118662 348265
rect 118606 348191 118662 348200
rect 117872 347812 117924 347818
rect 117872 347754 117924 347760
rect 117412 347744 117464 347750
rect 117412 347686 117464 347692
rect 117424 347585 117452 347686
rect 117410 347576 117466 347585
rect 117410 347511 117466 347520
rect 118608 346384 118660 346390
rect 118608 346326 118660 346332
rect 118514 346216 118570 346225
rect 118514 346151 118570 346160
rect 118528 345710 118556 346151
rect 118516 345704 118568 345710
rect 118516 345646 118568 345652
rect 118620 345545 118648 346326
rect 118606 345536 118662 345545
rect 118606 345471 118662 345480
rect 118608 345024 118660 345030
rect 118608 344966 118660 344972
rect 118620 344865 118648 344966
rect 118606 344856 118662 344865
rect 118606 344791 118662 344800
rect 117780 343596 117832 343602
rect 117780 343538 117832 343544
rect 117792 342825 117820 343538
rect 118606 343496 118662 343505
rect 118606 343431 118662 343440
rect 118620 342922 118648 343431
rect 118608 342916 118660 342922
rect 118608 342858 118660 342864
rect 117778 342816 117834 342825
rect 117778 342751 117834 342760
rect 118608 342236 118660 342242
rect 118608 342178 118660 342184
rect 118620 342145 118648 342178
rect 118606 342136 118662 342145
rect 118606 342071 118662 342080
rect 117502 340776 117558 340785
rect 117502 340711 117558 340720
rect 117516 340270 117544 340711
rect 117504 340264 117556 340270
rect 117504 340206 117556 340212
rect 118424 340196 118476 340202
rect 118424 340138 118476 340144
rect 118436 340105 118464 340138
rect 117318 340096 117374 340105
rect 117318 340031 117374 340040
rect 118422 340096 118478 340105
rect 118422 340031 118478 340040
rect 116584 331968 116636 331974
rect 116584 331910 116636 331916
rect 116032 315308 116084 315314
rect 116032 315250 116084 315256
rect 115940 302388 115992 302394
rect 115940 302330 115992 302336
rect 115388 294296 115440 294302
rect 115388 294238 115440 294244
rect 115296 294160 115348 294166
rect 115296 294102 115348 294108
rect 114558 291952 114614 291961
rect 78048 291910 78418 291938
rect 79336 291910 79706 291938
rect 81912 291910 82282 291938
rect 84396 291910 84858 291938
rect 85592 291910 86146 291938
rect 86972 291910 87434 291938
rect 94792 291910 95162 291938
rect 97184 291910 97738 291938
rect 103980 291916 104032 291922
rect 104912 291910 105466 291938
rect 114494 291910 114558 291938
rect 115308 291938 115336 294102
rect 115952 291977 115980 302330
rect 116596 293350 116624 331910
rect 117332 327729 117360 340031
rect 118712 335238 118740 387058
rect 118804 338978 118832 389302
rect 119356 389162 119384 389302
rect 119344 389156 119396 389162
rect 119344 389098 119396 389104
rect 119344 388068 119396 388074
rect 119344 388010 119396 388016
rect 119356 378826 119384 388010
rect 119344 378820 119396 378826
rect 119344 378762 119396 378768
rect 119068 365696 119120 365702
rect 119068 365638 119120 365644
rect 119080 364857 119108 365638
rect 119896 365084 119948 365090
rect 119896 365026 119948 365032
rect 119908 364886 119936 365026
rect 119896 364880 119948 364886
rect 119066 364848 119122 364857
rect 119896 364822 119948 364828
rect 119066 364783 119122 364792
rect 118884 360324 118936 360330
rect 118884 360266 118936 360272
rect 118896 359825 118924 360266
rect 118882 359816 118938 359825
rect 118882 359751 118938 359760
rect 119344 354000 119396 354006
rect 119344 353942 119396 353948
rect 118792 338972 118844 338978
rect 118792 338914 118844 338920
rect 119356 338065 119384 353942
rect 119342 338056 119398 338065
rect 119342 337991 119398 338000
rect 118700 335232 118752 335238
rect 118700 335174 118752 335180
rect 117964 331900 118016 331906
rect 117964 331842 118016 331848
rect 117318 327720 117374 327729
rect 117318 327655 117374 327664
rect 117976 311778 118004 331842
rect 117964 311772 118016 311778
rect 117964 311714 118016 311720
rect 116676 309800 116728 309806
rect 116676 309742 116728 309748
rect 116688 302394 116716 309742
rect 118882 307728 118938 307737
rect 118882 307663 118938 307672
rect 118896 306406 118924 307663
rect 118884 306400 118936 306406
rect 118884 306342 118936 306348
rect 116676 302388 116728 302394
rect 116676 302330 116728 302336
rect 117688 298376 117740 298382
rect 117688 298318 117740 298324
rect 117228 294228 117280 294234
rect 117228 294170 117280 294176
rect 117136 294092 117188 294098
rect 117136 294034 117188 294040
rect 116584 293344 116636 293350
rect 116584 293286 116636 293292
rect 117148 291990 117176 294034
rect 117240 293282 117268 294170
rect 117228 293276 117280 293282
rect 117228 293218 117280 293224
rect 117136 291984 117188 291990
rect 115952 291949 116426 291977
rect 115308 291910 115770 291938
rect 117700 291963 117728 298318
rect 119908 295633 119936 364822
rect 120000 360330 120028 466346
rect 120092 388550 120120 492662
rect 120172 476128 120224 476134
rect 120172 476070 120224 476076
rect 120080 388544 120132 388550
rect 120080 388486 120132 388492
rect 120080 385212 120132 385218
rect 120080 385154 120132 385160
rect 119988 360324 120040 360330
rect 119988 360266 120040 360272
rect 119894 295624 119950 295633
rect 119894 295559 119950 295568
rect 119620 294704 119672 294710
rect 119620 294646 119672 294652
rect 118330 292904 118386 292913
rect 118330 292839 118386 292848
rect 118344 292534 118372 292839
rect 118332 292528 118384 292534
rect 118332 292470 118384 292476
rect 118344 291963 118372 292470
rect 117136 291926 117188 291932
rect 119632 291924 119660 294646
rect 119804 292528 119856 292534
rect 119804 292470 119856 292476
rect 117228 291916 117280 291922
rect 114558 291887 114614 291896
rect 104032 291864 104178 291870
rect 103980 291858 104178 291864
rect 103992 291842 104178 291858
rect 117070 291864 117228 291870
rect 119344 291916 119396 291922
rect 117070 291858 117280 291864
rect 119002 291864 119344 291870
rect 119002 291858 119396 291864
rect 117070 291842 117268 291858
rect 119002 291842 119384 291858
rect 69846 288824 69902 288833
rect 69846 288759 69902 288768
rect 119816 287054 119844 292470
rect 119988 291916 120040 291922
rect 119988 291858 120040 291864
rect 119896 291848 119948 291854
rect 119896 291790 119948 291796
rect 119908 291242 119936 291790
rect 120000 291310 120028 291858
rect 119988 291304 120040 291310
rect 119988 291246 120040 291252
rect 119896 291236 119948 291242
rect 119896 291178 119948 291184
rect 119816 287026 120028 287054
rect 69110 286784 69166 286793
rect 69110 286719 69166 286728
rect 69018 282160 69074 282169
rect 69018 282095 69074 282104
rect 69018 274272 69074 274281
rect 69018 274207 69074 274216
rect 68926 232656 68982 232665
rect 68926 232591 68982 232600
rect 69032 196654 69060 274207
rect 120000 268394 120028 287026
rect 119988 268388 120040 268394
rect 119988 268330 120040 268336
rect 69110 252648 69166 252657
rect 69110 252583 69166 252592
rect 69020 196648 69072 196654
rect 69020 196590 69072 196596
rect 67548 185632 67600 185638
rect 67548 185574 67600 185580
rect 69124 178838 69152 252583
rect 120092 247625 120120 385154
rect 120184 369170 120212 476070
rect 120276 439550 120304 497490
rect 120356 494964 120408 494970
rect 120356 494906 120408 494912
rect 120264 439544 120316 439550
rect 120264 439486 120316 439492
rect 120368 438734 120396 494906
rect 121472 489870 121500 582966
rect 121564 538966 121592 583743
rect 122840 582480 122892 582486
rect 122840 582422 122892 582428
rect 122748 575544 122800 575550
rect 122748 575486 122800 575492
rect 122104 574048 122156 574054
rect 122104 573990 122156 573996
rect 122116 573374 122144 573990
rect 122104 573368 122156 573374
rect 122104 573310 122156 573316
rect 122116 572801 122144 573310
rect 122102 572792 122158 572801
rect 122102 572727 122158 572736
rect 121552 538960 121604 538966
rect 121552 538902 121604 538908
rect 121644 537600 121696 537606
rect 121644 537542 121696 537548
rect 121552 495508 121604 495514
rect 121552 495450 121604 495456
rect 121460 489864 121512 489870
rect 121460 489806 121512 489812
rect 121472 489190 121500 489806
rect 121460 489184 121512 489190
rect 121460 489126 121512 489132
rect 121460 484424 121512 484430
rect 121460 484366 121512 484372
rect 120356 438728 120408 438734
rect 120356 438670 120408 438676
rect 120908 438728 120960 438734
rect 120908 438670 120960 438676
rect 120920 438258 120948 438670
rect 120908 438252 120960 438258
rect 120908 438194 120960 438200
rect 120724 396908 120776 396914
rect 120724 396850 120776 396856
rect 120264 396024 120316 396030
rect 120264 395966 120316 395972
rect 120276 387802 120304 395966
rect 120264 387796 120316 387802
rect 120264 387738 120316 387744
rect 120276 387025 120304 387738
rect 120262 387016 120318 387025
rect 120262 386951 120318 386960
rect 120264 385688 120316 385694
rect 120264 385630 120316 385636
rect 120276 376310 120304 385630
rect 120264 376304 120316 376310
rect 120264 376246 120316 376252
rect 120172 369164 120224 369170
rect 120172 369106 120224 369112
rect 120170 338056 120226 338065
rect 120170 337991 120226 338000
rect 120184 337890 120212 337991
rect 120172 337884 120224 337890
rect 120172 337826 120224 337832
rect 120184 336802 120212 337826
rect 120172 336796 120224 336802
rect 120172 336738 120224 336744
rect 120736 329866 120764 396850
rect 121472 380866 121500 484366
rect 121564 392630 121592 495450
rect 121656 438802 121684 537542
rect 122760 485761 122788 575486
rect 122852 494766 122880 582422
rect 122932 581052 122984 581058
rect 122932 580994 122984 581000
rect 122944 497486 122972 580994
rect 123036 532030 123064 586570
rect 128452 586560 128504 586566
rect 128452 586502 128504 586508
rect 125692 583840 125744 583846
rect 125692 583782 125744 583788
rect 124312 564392 124364 564398
rect 124312 564334 124364 564340
rect 124220 559020 124272 559026
rect 124220 558962 124272 558968
rect 123484 538280 123536 538286
rect 123484 538222 123536 538228
rect 123024 532024 123076 532030
rect 123024 531966 123076 531972
rect 122932 497480 122984 497486
rect 122932 497422 122984 497428
rect 122840 494760 122892 494766
rect 122840 494702 122892 494708
rect 122840 493400 122892 493406
rect 122840 493342 122892 493348
rect 122746 485752 122802 485761
rect 122746 485687 122802 485696
rect 121736 466268 121788 466274
rect 121736 466210 121788 466216
rect 121644 438796 121696 438802
rect 121644 438738 121696 438744
rect 121656 438326 121684 438738
rect 121644 438320 121696 438326
rect 121644 438262 121696 438268
rect 121748 393314 121776 466210
rect 121656 393286 121776 393314
rect 121552 392624 121604 392630
rect 121552 392566 121604 392572
rect 121552 392148 121604 392154
rect 121552 392090 121604 392096
rect 121460 380860 121512 380866
rect 121460 380802 121512 380808
rect 121368 362228 121420 362234
rect 121368 362170 121420 362176
rect 120172 329860 120224 329866
rect 120172 329802 120224 329808
rect 120724 329860 120776 329866
rect 120724 329802 120776 329808
rect 120184 329730 120212 329802
rect 120172 329724 120224 329730
rect 120172 329666 120224 329672
rect 120172 311364 120224 311370
rect 120172 311306 120224 311312
rect 120184 256465 120212 311306
rect 120170 256456 120226 256465
rect 120170 256391 120226 256400
rect 120170 251016 120226 251025
rect 120170 250951 120226 250960
rect 120078 247616 120134 247625
rect 120078 247551 120134 247560
rect 69202 245032 69258 245041
rect 69202 244967 69258 244976
rect 69216 237386 69244 244967
rect 119896 240168 119948 240174
rect 69952 240094 70058 240122
rect 119646 240116 119896 240122
rect 119646 240110 119948 240116
rect 119646 240094 119936 240110
rect 69952 238134 69980 240094
rect 70688 238754 70716 240037
rect 71320 239850 71348 240037
rect 70412 238726 70716 238754
rect 71240 239822 71348 239850
rect 69940 238128 69992 238134
rect 69940 238070 69992 238076
rect 69204 237380 69256 237386
rect 69204 237322 69256 237328
rect 70412 200802 70440 238726
rect 71240 227118 71268 239822
rect 71976 238754 72004 240037
rect 72424 239556 72476 239562
rect 72424 239498 72476 239504
rect 71792 238726 72004 238754
rect 71228 227112 71280 227118
rect 71228 227054 71280 227060
rect 71792 213382 71820 238726
rect 71780 213376 71832 213382
rect 71780 213318 71832 213324
rect 70400 200796 70452 200802
rect 70400 200738 70452 200744
rect 72436 186998 72464 239498
rect 72620 238649 72648 240037
rect 73252 239850 73280 240037
rect 73172 239822 73280 239850
rect 72606 238640 72662 238649
rect 72606 238575 72662 238584
rect 73172 187134 73200 239822
rect 73908 238066 73936 240037
rect 73896 238060 73948 238066
rect 73896 238002 73948 238008
rect 74552 209166 74580 240037
rect 75196 238754 75224 240037
rect 75828 239850 75856 240037
rect 74644 238726 75224 238754
rect 75748 239822 75856 239850
rect 75920 239828 75972 239834
rect 74644 220114 74672 238726
rect 75748 224942 75776 239822
rect 75920 239770 75972 239776
rect 75736 224936 75788 224942
rect 75736 224878 75788 224884
rect 74632 220108 74684 220114
rect 74632 220050 74684 220056
rect 75932 210458 75960 239770
rect 76484 238882 76512 240037
rect 77116 239834 77144 240037
rect 77104 239828 77156 239834
rect 77104 239770 77156 239776
rect 76012 238876 76064 238882
rect 76012 238818 76064 238824
rect 76472 238876 76524 238882
rect 76472 238818 76524 238824
rect 76024 211886 76052 238818
rect 77772 232626 77800 240037
rect 78416 238754 78444 240037
rect 79060 238754 79088 240037
rect 79692 239850 79720 240037
rect 77864 238726 78444 238754
rect 78692 238726 79088 238754
rect 79612 239822 79720 239850
rect 80060 239828 80112 239834
rect 77760 232620 77812 232626
rect 77760 232562 77812 232568
rect 77864 219434 77892 238726
rect 77944 238128 77996 238134
rect 77944 238070 77996 238076
rect 77312 219406 77892 219434
rect 76012 211880 76064 211886
rect 76012 211822 76064 211828
rect 75920 210452 75972 210458
rect 75920 210394 75972 210400
rect 74540 209160 74592 209166
rect 74540 209102 74592 209108
rect 77312 199578 77340 219406
rect 77956 216034 77984 238070
rect 77944 216028 77996 216034
rect 77944 215970 77996 215976
rect 77300 199572 77352 199578
rect 77300 199514 77352 199520
rect 78692 189922 78720 238726
rect 79612 219434 79640 239822
rect 80060 239770 80112 239776
rect 80072 225622 80100 239770
rect 80348 238754 80376 240037
rect 80980 239834 81008 240037
rect 80968 239828 81020 239834
rect 80968 239770 81020 239776
rect 80164 238726 80376 238754
rect 80164 229809 80192 238726
rect 81636 237250 81664 240037
rect 82280 238754 82308 240037
rect 82912 239850 82940 240037
rect 83556 239850 83584 240037
rect 82004 238726 82308 238754
rect 82832 239822 82940 239850
rect 83476 239822 83584 239850
rect 81624 237244 81676 237250
rect 81624 237186 81676 237192
rect 81636 236026 81664 237186
rect 81624 236020 81676 236026
rect 81624 235962 81676 235968
rect 80150 229800 80206 229809
rect 80150 229735 80206 229744
rect 80060 225616 80112 225622
rect 80060 225558 80112 225564
rect 82004 219434 82032 238726
rect 82084 236020 82136 236026
rect 82084 235962 82136 235968
rect 78784 219406 79640 219434
rect 81544 219406 82032 219434
rect 78784 214742 78812 219406
rect 81544 216646 81572 219406
rect 81532 216640 81584 216646
rect 81532 216582 81584 216588
rect 78772 214736 78824 214742
rect 78772 214678 78824 214684
rect 78680 189916 78732 189922
rect 78680 189858 78732 189864
rect 73160 187128 73212 187134
rect 73160 187070 73212 187076
rect 72424 186992 72476 186998
rect 72424 186934 72476 186940
rect 82096 180130 82124 235962
rect 82832 229022 82860 239822
rect 83476 229090 83504 239822
rect 84212 229974 84240 240037
rect 84856 238754 84884 240037
rect 84396 238726 84884 238754
rect 84200 229968 84252 229974
rect 84200 229910 84252 229916
rect 84396 229786 84424 238726
rect 85500 237454 85528 240037
rect 85488 237448 85540 237454
rect 85488 237390 85540 237396
rect 86144 237182 86172 240037
rect 86788 238678 86816 240037
rect 87432 238754 87460 240037
rect 88064 239850 88092 240037
rect 86972 238726 87460 238754
rect 87984 239822 88092 239850
rect 86776 238672 86828 238678
rect 86776 238614 86828 238620
rect 86788 237522 86816 238614
rect 86224 237516 86276 237522
rect 86224 237458 86276 237464
rect 86776 237516 86828 237522
rect 86776 237458 86828 237464
rect 86132 237176 86184 237182
rect 86132 237118 86184 237124
rect 86144 233918 86172 237118
rect 86132 233912 86184 233918
rect 86132 233854 86184 233860
rect 84476 229968 84528 229974
rect 84476 229910 84528 229916
rect 84212 229758 84424 229786
rect 83464 229084 83516 229090
rect 83464 229026 83516 229032
rect 82820 229016 82872 229022
rect 82820 228958 82872 228964
rect 83476 221474 83504 229026
rect 83464 221468 83516 221474
rect 83464 221410 83516 221416
rect 82084 180124 82136 180130
rect 82084 180066 82136 180072
rect 84212 178906 84240 229758
rect 84488 229650 84516 229910
rect 84304 229622 84516 229650
rect 84304 220153 84332 229622
rect 84290 220144 84346 220153
rect 84290 220079 84346 220088
rect 86236 206310 86264 237458
rect 86316 237448 86368 237454
rect 86316 237390 86368 237396
rect 86328 206378 86356 237390
rect 86316 206372 86368 206378
rect 86316 206314 86368 206320
rect 86224 206304 86276 206310
rect 86224 206246 86276 206252
rect 86972 184414 87000 238726
rect 87984 219434 88012 239822
rect 88720 238754 88748 240037
rect 87064 219406 88012 219434
rect 88352 238726 88748 238754
rect 89364 238754 89392 240037
rect 89364 238726 89668 238754
rect 87064 207806 87092 219406
rect 87052 207800 87104 207806
rect 87052 207742 87104 207748
rect 88352 187202 88380 238726
rect 89640 235958 89668 238726
rect 90008 237454 90036 240037
rect 90652 238754 90680 240037
rect 91296 238754 91324 240037
rect 90100 238726 90680 238754
rect 91112 238726 91324 238754
rect 89996 237448 90048 237454
rect 89996 237390 90048 237396
rect 89628 235952 89680 235958
rect 89628 235894 89680 235900
rect 89640 195294 89668 235894
rect 90100 224330 90128 238726
rect 90362 237960 90418 237969
rect 90362 237895 90418 237904
rect 90088 224324 90140 224330
rect 90088 224266 90140 224272
rect 90376 203658 90404 237895
rect 91112 227730 91140 238726
rect 91940 238678 91968 240037
rect 92480 239828 92532 239834
rect 92480 239770 92532 239776
rect 91928 238672 91980 238678
rect 91928 238614 91980 238620
rect 91744 237448 91796 237454
rect 91744 237390 91796 237396
rect 91100 227724 91152 227730
rect 91100 227666 91152 227672
rect 91756 203726 91784 237390
rect 91744 203720 91796 203726
rect 91744 203662 91796 203668
rect 90364 203652 90416 203658
rect 90364 203594 90416 203600
rect 92492 196722 92520 239770
rect 92584 198150 92612 240037
rect 93216 239834 93244 240037
rect 93204 239828 93256 239834
rect 93204 239770 93256 239776
rect 92664 239420 92716 239426
rect 92664 239362 92716 239368
rect 92676 238610 92704 239362
rect 92664 238604 92716 238610
rect 92664 238546 92716 238552
rect 93872 233866 93900 240037
rect 94516 238754 94544 240037
rect 95148 239850 95176 240037
rect 94056 238726 94544 238754
rect 95068 239822 95176 239850
rect 95240 239828 95292 239834
rect 93872 233838 93992 233866
rect 93860 233776 93912 233782
rect 93860 233718 93912 233724
rect 92572 198144 92624 198150
rect 92572 198086 92624 198092
rect 92480 196716 92532 196722
rect 92480 196658 92532 196664
rect 89628 195288 89680 195294
rect 89628 195230 89680 195236
rect 93872 193866 93900 233718
rect 93964 213246 93992 233838
rect 94056 233782 94084 238726
rect 94044 233776 94096 233782
rect 94044 233718 94096 233724
rect 95068 231198 95096 239822
rect 95240 239770 95292 239776
rect 95056 231192 95108 231198
rect 95056 231134 95108 231140
rect 93952 213240 94004 213246
rect 93952 213182 94004 213188
rect 93860 193860 93912 193866
rect 93860 193802 93912 193808
rect 88340 187196 88392 187202
rect 88340 187138 88392 187144
rect 86960 184408 87012 184414
rect 86960 184350 87012 184356
rect 95252 184278 95280 239770
rect 95804 238754 95832 240037
rect 96436 239834 96464 240037
rect 96424 239828 96476 239834
rect 96424 239770 96476 239776
rect 96620 239828 96672 239834
rect 96620 239770 96672 239776
rect 95344 238726 95832 238754
rect 95344 231742 95372 238726
rect 95332 231736 95384 231742
rect 95332 231678 95384 231684
rect 95240 184272 95292 184278
rect 95240 184214 95292 184220
rect 96632 182850 96660 239770
rect 97092 238754 97120 240037
rect 97724 239834 97752 240037
rect 97712 239828 97764 239834
rect 97712 239770 97764 239776
rect 96724 238726 97120 238754
rect 98380 238746 98408 240037
rect 99012 239850 99040 240037
rect 98564 239822 99040 239850
rect 98368 238740 98420 238746
rect 96724 184346 96752 238726
rect 98368 238682 98420 238688
rect 98564 219434 98592 239822
rect 98644 239488 98696 239494
rect 98644 239430 98696 239436
rect 98104 219406 98592 219434
rect 98104 205630 98132 219406
rect 98092 205624 98144 205630
rect 98092 205566 98144 205572
rect 98656 202230 98684 239430
rect 99668 238754 99696 240037
rect 100300 239850 100328 240037
rect 100944 239850 100972 240037
rect 99392 238726 99696 238754
rect 100220 239822 100328 239850
rect 100760 239828 100812 239834
rect 98644 202224 98696 202230
rect 98644 202166 98696 202172
rect 99392 188426 99420 238726
rect 100220 219434 100248 239822
rect 100760 239770 100812 239776
rect 100864 239822 100972 239850
rect 101588 239834 101616 240037
rect 101576 239828 101628 239834
rect 99484 219406 100248 219434
rect 99484 202298 99512 219406
rect 100772 203794 100800 239770
rect 100864 209234 100892 239822
rect 101576 239770 101628 239776
rect 102244 238134 102272 240037
rect 102876 239850 102904 240037
rect 102796 239822 102904 239850
rect 102232 238128 102284 238134
rect 102232 238070 102284 238076
rect 102796 219434 102824 239822
rect 103532 238610 103560 240037
rect 104176 239442 104204 240037
rect 104808 239850 104836 240037
rect 103992 239414 104204 239442
rect 104728 239822 104836 239850
rect 104900 239828 104952 239834
rect 103992 238754 104020 239414
rect 104728 238754 104756 239822
rect 104900 239770 104952 239776
rect 103624 238726 104020 238754
rect 104084 238726 104756 238754
rect 103520 238604 103572 238610
rect 103520 238546 103572 238552
rect 103532 237454 103560 238546
rect 103520 237448 103572 237454
rect 103520 237390 103572 237396
rect 103624 221610 103652 238726
rect 103612 221604 103664 221610
rect 103612 221546 103664 221552
rect 104084 219434 104112 238726
rect 104164 237448 104216 237454
rect 104164 237390 104216 237396
rect 104176 221474 104204 237390
rect 104164 221468 104216 221474
rect 104164 221410 104216 221416
rect 102152 219406 102824 219434
rect 103716 219406 104112 219434
rect 100852 209228 100904 209234
rect 100852 209170 100904 209176
rect 100760 203788 100812 203794
rect 100760 203730 100812 203736
rect 99472 202292 99524 202298
rect 99472 202234 99524 202240
rect 102152 193934 102180 219406
rect 103716 195430 103744 219406
rect 103704 195424 103756 195430
rect 103704 195366 103756 195372
rect 102140 193928 102192 193934
rect 102140 193870 102192 193876
rect 100668 190596 100720 190602
rect 100668 190538 100720 190544
rect 99380 188420 99432 188426
rect 99380 188362 99432 188368
rect 96712 184340 96764 184346
rect 96712 184282 96764 184288
rect 96620 182844 96672 182850
rect 96620 182786 96672 182792
rect 97080 180872 97132 180878
rect 97080 180814 97132 180820
rect 84200 178900 84252 178906
rect 84200 178842 84252 178848
rect 69112 178832 69164 178838
rect 69112 178774 69164 178780
rect 66168 178764 66220 178770
rect 66168 178706 66220 178712
rect 97092 177721 97120 180814
rect 97078 177712 97134 177721
rect 97078 177647 97134 177656
rect 100680 176769 100708 190538
rect 102048 189100 102100 189106
rect 102048 189042 102100 189048
rect 100760 178696 100812 178702
rect 100760 178638 100812 178644
rect 100772 177342 100800 178638
rect 102060 177721 102088 189042
rect 104912 187066 104940 239770
rect 105464 238270 105492 240037
rect 106096 239834 106124 240037
rect 106084 239828 106136 239834
rect 106084 239770 106136 239776
rect 106752 238754 106780 240037
rect 107384 239850 107412 240037
rect 106292 238726 106780 238754
rect 107304 239822 107412 239850
rect 105452 238264 105504 238270
rect 105452 238206 105504 238212
rect 106292 208350 106320 238726
rect 107304 231810 107332 239822
rect 108040 238754 108068 240037
rect 108672 239850 108700 240037
rect 109960 239850 109988 240037
rect 107672 238726 108068 238754
rect 108592 239822 108700 239850
rect 109880 239822 109988 239850
rect 107292 231804 107344 231810
rect 107292 231746 107344 231752
rect 107304 219434 107332 231746
rect 106936 219406 107332 219434
rect 106280 208344 106332 208350
rect 106280 208286 106332 208292
rect 106936 197985 106964 219406
rect 106922 197976 106978 197985
rect 106922 197911 106978 197920
rect 106188 190528 106240 190534
rect 106188 190470 106240 190476
rect 104900 187060 104952 187066
rect 104900 187002 104952 187008
rect 106200 177721 106228 190470
rect 107672 184210 107700 238726
rect 108592 229838 108620 239822
rect 109880 238754 109908 239822
rect 109696 238726 109908 238754
rect 109696 234598 109724 238726
rect 110616 237250 110644 240037
rect 111260 238754 111288 240037
rect 111892 239850 111920 240037
rect 110984 238726 111288 238754
rect 111812 239822 111920 239850
rect 110604 237244 110656 237250
rect 110604 237186 110656 237192
rect 110616 236026 110644 237186
rect 110604 236020 110656 236026
rect 110604 235962 110656 235968
rect 109684 234592 109736 234598
rect 109684 234534 109736 234540
rect 108580 229832 108632 229838
rect 108580 229774 108632 229780
rect 109696 223650 109724 234534
rect 109684 223644 109736 223650
rect 109684 223586 109736 223592
rect 107660 184204 107712 184210
rect 107660 184146 107712 184152
rect 109696 180198 109724 223586
rect 110984 219434 111012 238726
rect 111064 236020 111116 236026
rect 111064 235962 111116 235968
rect 110432 219406 111012 219434
rect 110432 182986 110460 219406
rect 110420 182980 110472 182986
rect 110420 182922 110472 182928
rect 110696 182232 110748 182238
rect 110696 182174 110748 182180
rect 109684 180192 109736 180198
rect 109684 180134 109736 180140
rect 108120 179444 108172 179450
rect 108120 179386 108172 179392
rect 102046 177712 102102 177721
rect 102046 177647 102102 177656
rect 106186 177712 106242 177721
rect 106186 177647 106242 177656
rect 100760 177336 100812 177342
rect 100760 177278 100812 177284
rect 108132 177041 108160 179386
rect 109960 177948 110012 177954
rect 109960 177890 110012 177896
rect 108118 177032 108174 177041
rect 108118 176967 108174 176976
rect 107016 176928 107068 176934
rect 107016 176870 107068 176876
rect 103336 176860 103388 176866
rect 103336 176802 103388 176808
rect 103348 176769 103376 176802
rect 107028 176769 107056 176870
rect 109972 176769 110000 177890
rect 110708 177721 110736 182174
rect 110694 177712 110750 177721
rect 110694 177647 110750 177656
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 103334 176760 103390 176769
rect 103334 176695 103390 176704
rect 107014 176760 107070 176769
rect 107014 176695 107070 176704
rect 109958 176760 110014 176769
rect 109958 176695 110014 176704
rect 104624 176112 104676 176118
rect 104624 176054 104676 176060
rect 104636 175545 104664 176054
rect 111076 175982 111104 235962
rect 111812 196858 111840 239822
rect 112548 238814 112576 240037
rect 113192 239442 113220 240037
rect 113192 239414 113312 239442
rect 113180 239352 113232 239358
rect 113180 239294 113232 239300
rect 112536 238808 112588 238814
rect 112536 238750 112588 238756
rect 112548 233986 112576 238750
rect 112536 233980 112588 233986
rect 112536 233922 112588 233928
rect 113192 215286 113220 239294
rect 113284 235278 113312 239414
rect 113836 238649 113864 240037
rect 114480 239358 114508 240037
rect 114560 239828 114612 239834
rect 114560 239770 114612 239776
rect 114468 239352 114520 239358
rect 114468 239294 114520 239300
rect 113822 238640 113878 238649
rect 113822 238575 113878 238584
rect 113272 235272 113324 235278
rect 113272 235214 113324 235220
rect 113180 215280 113232 215286
rect 113180 215222 113232 215228
rect 114572 210594 114600 239770
rect 115124 238754 115152 240037
rect 115756 239834 115784 240037
rect 115744 239828 115796 239834
rect 115744 239770 115796 239776
rect 116412 238754 116440 240037
rect 114664 238726 115152 238754
rect 115952 238726 116440 238754
rect 114664 226273 114692 238726
rect 114650 226264 114706 226273
rect 114650 226199 114706 226208
rect 114560 210588 114612 210594
rect 114560 210530 114612 210536
rect 115952 199646 115980 238726
rect 117056 238513 117084 240037
rect 117320 239828 117372 239834
rect 117320 239770 117372 239776
rect 117042 238504 117098 238513
rect 117042 238439 117098 238448
rect 116584 237448 116636 237454
rect 116584 237390 116636 237396
rect 116596 237318 116624 237390
rect 116584 237312 116636 237318
rect 116584 237254 116636 237260
rect 115940 199640 115992 199646
rect 115940 199582 115992 199588
rect 111800 196852 111852 196858
rect 111800 196794 111852 196800
rect 116596 189786 116624 237254
rect 117332 200870 117360 239770
rect 117700 237454 117728 240037
rect 118344 239834 118372 240037
rect 118332 239828 118384 239834
rect 118332 239770 118384 239776
rect 118988 238754 119016 240037
rect 118988 238726 119384 238754
rect 117688 237448 117740 237454
rect 117688 237390 117740 237396
rect 119356 235929 119384 238726
rect 119342 235920 119398 235929
rect 119342 235855 119398 235864
rect 117320 200864 117372 200870
rect 117320 200806 117372 200812
rect 119356 191146 119384 235855
rect 120184 205018 120212 250951
rect 121380 241505 121408 362170
rect 121460 323740 121512 323746
rect 121460 323682 121512 323688
rect 121472 248402 121500 323682
rect 121564 311302 121592 392090
rect 121656 391950 121684 393286
rect 121644 391944 121696 391950
rect 121644 391886 121696 391892
rect 121656 358086 121684 391886
rect 122012 388544 122064 388550
rect 122012 388486 122064 388492
rect 122024 383654 122052 388486
rect 122852 387705 122880 493342
rect 123024 492040 123076 492046
rect 123024 491982 123076 491988
rect 122932 483676 122984 483682
rect 122932 483618 122984 483624
rect 122944 483313 122972 483618
rect 122930 483304 122986 483313
rect 122930 483239 122986 483248
rect 122932 438932 122984 438938
rect 122932 438874 122984 438880
rect 122102 387696 122158 387705
rect 122102 387631 122158 387640
rect 122838 387696 122894 387705
rect 122838 387631 122894 387640
rect 122116 386617 122144 387631
rect 122102 386608 122158 386617
rect 122102 386543 122104 386552
rect 122156 386543 122158 386552
rect 122104 386514 122156 386520
rect 122116 386483 122144 386514
rect 122024 383626 122144 383654
rect 122116 365022 122144 383626
rect 122196 380860 122248 380866
rect 122196 380802 122248 380808
rect 122208 380225 122236 380802
rect 122194 380216 122250 380225
rect 122194 380151 122250 380160
rect 122840 378888 122892 378894
rect 122840 378830 122892 378836
rect 122196 378208 122248 378214
rect 122196 378150 122248 378156
rect 122104 365016 122156 365022
rect 122104 364958 122156 364964
rect 121644 358080 121696 358086
rect 121644 358022 121696 358028
rect 122104 345704 122156 345710
rect 122104 345646 122156 345652
rect 121644 319456 121696 319462
rect 121644 319398 121696 319404
rect 121552 311296 121604 311302
rect 121552 311238 121604 311244
rect 121550 291816 121606 291825
rect 121550 291751 121552 291760
rect 121604 291751 121606 291760
rect 121552 291722 121604 291728
rect 121550 291136 121606 291145
rect 121550 291071 121606 291080
rect 121564 289882 121592 291071
rect 121552 289876 121604 289882
rect 121552 289818 121604 289824
rect 121552 288380 121604 288386
rect 121552 288322 121604 288328
rect 121564 287745 121592 288322
rect 121550 287736 121606 287745
rect 121550 287671 121606 287680
rect 121550 287056 121606 287065
rect 121656 287054 121684 319398
rect 121734 289096 121790 289105
rect 121734 289031 121790 289040
rect 121748 288454 121776 289031
rect 121736 288448 121788 288454
rect 121736 288390 121788 288396
rect 121826 288416 121882 288425
rect 121826 288351 121882 288360
rect 121840 287094 121868 288351
rect 121828 287088 121880 287094
rect 121656 287026 121776 287054
rect 121828 287030 121880 287036
rect 121550 286991 121552 287000
rect 121604 286991 121606 287000
rect 121552 286962 121604 286968
rect 121550 286376 121606 286385
rect 121550 286311 121552 286320
rect 121604 286311 121606 286320
rect 121552 286282 121604 286288
rect 121550 285016 121606 285025
rect 121550 284951 121606 284960
rect 121564 284442 121592 284951
rect 121552 284436 121604 284442
rect 121552 284378 121604 284384
rect 121644 284368 121696 284374
rect 121642 284336 121644 284345
rect 121696 284336 121698 284345
rect 121642 284271 121698 284280
rect 121550 283656 121606 283665
rect 121550 283591 121552 283600
rect 121604 283591 121606 283600
rect 121552 283562 121604 283568
rect 121550 282976 121606 282985
rect 121550 282911 121552 282920
rect 121604 282911 121606 282920
rect 121552 282882 121604 282888
rect 121642 282296 121698 282305
rect 121642 282231 121698 282240
rect 121656 281654 121684 282231
rect 121644 281648 121696 281654
rect 121550 281616 121606 281625
rect 121644 281590 121696 281596
rect 121550 281551 121552 281560
rect 121604 281551 121606 281560
rect 121552 281522 121604 281528
rect 121642 280936 121698 280945
rect 121642 280871 121698 280880
rect 121552 280288 121604 280294
rect 121550 280256 121552 280265
rect 121604 280256 121606 280265
rect 121656 280226 121684 280871
rect 121550 280191 121606 280200
rect 121644 280220 121696 280226
rect 121644 280162 121696 280168
rect 121642 279576 121698 279585
rect 121642 279511 121698 279520
rect 121550 278896 121606 278905
rect 121550 278831 121552 278840
rect 121604 278831 121606 278840
rect 121552 278802 121604 278808
rect 121656 278798 121684 279511
rect 121644 278792 121696 278798
rect 121644 278734 121696 278740
rect 121550 277536 121606 277545
rect 121550 277471 121606 277480
rect 121564 277438 121592 277471
rect 121552 277432 121604 277438
rect 121552 277374 121604 277380
rect 121748 276865 121776 287026
rect 121734 276856 121790 276865
rect 121734 276791 121790 276800
rect 121550 276176 121606 276185
rect 121550 276111 121606 276120
rect 121564 276078 121592 276111
rect 121552 276072 121604 276078
rect 121552 276014 121604 276020
rect 121644 276004 121696 276010
rect 121644 275946 121696 275952
rect 121656 275505 121684 275946
rect 121642 275496 121698 275505
rect 121642 275431 121698 275440
rect 121748 275398 121776 276791
rect 121736 275392 121788 275398
rect 121736 275334 121788 275340
rect 121550 274816 121606 274825
rect 121550 274751 121606 274760
rect 121564 274718 121592 274751
rect 121552 274712 121604 274718
rect 121552 274654 121604 274660
rect 121552 274576 121604 274582
rect 121552 274518 121604 274524
rect 121564 274145 121592 274518
rect 121550 274136 121606 274145
rect 121550 274071 121606 274080
rect 121550 273456 121606 273465
rect 121550 273391 121606 273400
rect 121564 273290 121592 273391
rect 121552 273284 121604 273290
rect 121552 273226 121604 273232
rect 121552 273148 121604 273154
rect 121552 273090 121604 273096
rect 121564 272785 121592 273090
rect 121550 272776 121606 272785
rect 121550 272711 121606 272720
rect 121550 272096 121606 272105
rect 121550 272031 121606 272040
rect 121564 271930 121592 272031
rect 121552 271924 121604 271930
rect 121552 271866 121604 271872
rect 121550 271416 121606 271425
rect 121550 271351 121606 271360
rect 121564 270570 121592 271351
rect 121552 270564 121604 270570
rect 121552 270506 121604 270512
rect 121642 270056 121698 270065
rect 121642 269991 121698 270000
rect 121550 269376 121606 269385
rect 121550 269311 121606 269320
rect 121564 269210 121592 269311
rect 121552 269204 121604 269210
rect 121552 269146 121604 269152
rect 121656 269142 121684 269991
rect 121644 269136 121696 269142
rect 121644 269078 121696 269084
rect 121642 268696 121698 268705
rect 121642 268631 121698 268640
rect 121550 268016 121606 268025
rect 121550 267951 121606 267960
rect 121564 267782 121592 267951
rect 121656 267850 121684 268631
rect 121644 267844 121696 267850
rect 121644 267786 121696 267792
rect 121552 267776 121604 267782
rect 121552 267718 121604 267724
rect 121642 267336 121698 267345
rect 121642 267271 121698 267280
rect 121550 266656 121606 266665
rect 121550 266591 121606 266600
rect 121564 266490 121592 266591
rect 121552 266484 121604 266490
rect 121552 266426 121604 266432
rect 121656 266422 121684 267271
rect 121644 266416 121696 266422
rect 121644 266358 121696 266364
rect 121642 265976 121698 265985
rect 121642 265911 121698 265920
rect 121550 265296 121606 265305
rect 121550 265231 121606 265240
rect 121564 264994 121592 265231
rect 121552 264988 121604 264994
rect 121552 264930 121604 264936
rect 121656 264246 121684 265911
rect 121734 264616 121790 264625
rect 121734 264551 121790 264560
rect 121644 264240 121696 264246
rect 121644 264182 121696 264188
rect 121550 263936 121606 263945
rect 121550 263871 121606 263880
rect 121564 263702 121592 263871
rect 121552 263696 121604 263702
rect 121552 263638 121604 263644
rect 121552 263560 121604 263566
rect 121552 263502 121604 263508
rect 121564 263265 121592 263502
rect 121748 263498 121776 264551
rect 121736 263492 121788 263498
rect 121736 263434 121788 263440
rect 121550 263256 121606 263265
rect 121550 263191 121606 263200
rect 121550 262576 121606 262585
rect 121550 262511 121606 262520
rect 121564 262274 121592 262511
rect 121552 262268 121604 262274
rect 121552 262210 121604 262216
rect 121644 262200 121696 262206
rect 121644 262142 121696 262148
rect 121656 261225 121684 262142
rect 121734 261896 121790 261905
rect 121734 261831 121790 261840
rect 121642 261216 121698 261225
rect 121642 261151 121698 261160
rect 121552 260840 121604 260846
rect 121552 260782 121604 260788
rect 121564 260545 121592 260782
rect 121550 260536 121606 260545
rect 121550 260471 121606 260480
rect 121748 260234 121776 261831
rect 121736 260228 121788 260234
rect 121736 260170 121788 260176
rect 121550 259856 121606 259865
rect 121550 259791 121606 259800
rect 121564 259486 121592 259791
rect 121552 259480 121604 259486
rect 121552 259422 121604 259428
rect 121644 259412 121696 259418
rect 121644 259354 121696 259360
rect 121550 259176 121606 259185
rect 121550 259111 121606 259120
rect 121564 258126 121592 259111
rect 121656 258505 121684 259354
rect 121642 258496 121698 258505
rect 121642 258431 121698 258440
rect 121552 258120 121604 258126
rect 121552 258062 121604 258068
rect 121642 257816 121698 257825
rect 121642 257751 121698 257760
rect 121550 257136 121606 257145
rect 121550 257071 121606 257080
rect 121564 256698 121592 257071
rect 121656 256766 121684 257751
rect 121644 256760 121696 256766
rect 121644 256702 121696 256708
rect 121552 256692 121604 256698
rect 121552 256634 121604 256640
rect 121642 256456 121698 256465
rect 121642 256391 121698 256400
rect 121550 254416 121606 254425
rect 121550 254351 121606 254360
rect 121564 253978 121592 254351
rect 121552 253972 121604 253978
rect 121552 253914 121604 253920
rect 121550 253736 121606 253745
rect 121550 253671 121606 253680
rect 121564 252686 121592 253671
rect 121656 253230 121684 256391
rect 121644 253224 121696 253230
rect 121644 253166 121696 253172
rect 121642 253056 121698 253065
rect 121642 252991 121698 253000
rect 121552 252680 121604 252686
rect 121552 252622 121604 252628
rect 121656 252618 121684 252991
rect 121644 252612 121696 252618
rect 121644 252554 121696 252560
rect 121552 252544 121604 252550
rect 121552 252486 121604 252492
rect 121564 252385 121592 252486
rect 121550 252376 121606 252385
rect 121550 252311 121606 252320
rect 121550 251696 121606 251705
rect 121550 251631 121606 251640
rect 121564 251258 121592 251631
rect 121552 251252 121604 251258
rect 121552 251194 121604 251200
rect 122116 251025 122144 345646
rect 122208 338910 122236 378150
rect 122196 338904 122248 338910
rect 122196 338846 122248 338852
rect 122562 314256 122618 314265
rect 122562 314191 122618 314200
rect 122576 313342 122604 314191
rect 122564 313336 122616 313342
rect 122564 313278 122616 313284
rect 122852 302938 122880 378830
rect 122944 336666 122972 438874
rect 123036 395350 123064 491982
rect 123496 439006 123524 538222
rect 124232 466342 124260 558962
rect 124324 471986 124352 564334
rect 124402 554024 124458 554033
rect 124402 553959 124458 553968
rect 124312 471980 124364 471986
rect 124312 471922 124364 471928
rect 124220 466336 124272 466342
rect 124220 466278 124272 466284
rect 124220 463752 124272 463758
rect 124220 463694 124272 463700
rect 123484 439000 123536 439006
rect 123760 439000 123812 439006
rect 123484 438942 123536 438948
rect 123758 438968 123760 438977
rect 123812 438968 123814 438977
rect 123758 438903 123814 438912
rect 123116 400988 123168 400994
rect 123116 400930 123168 400936
rect 123024 395344 123076 395350
rect 123024 395286 123076 395292
rect 123022 378992 123078 379001
rect 123022 378927 123078 378936
rect 123036 378894 123064 378927
rect 123024 378888 123076 378894
rect 123024 378830 123076 378836
rect 122932 336660 122984 336666
rect 122932 336602 122984 336608
rect 123128 328438 123156 400930
rect 123484 390720 123536 390726
rect 123484 390662 123536 390668
rect 123116 328432 123168 328438
rect 123116 328374 123168 328380
rect 122840 302932 122892 302938
rect 122840 302874 122892 302880
rect 123496 291786 123524 390662
rect 124232 354074 124260 463694
rect 124416 462330 124444 553959
rect 125600 550656 125652 550662
rect 125600 550598 125652 550604
rect 124954 541648 125010 541657
rect 124954 541583 125010 541592
rect 124404 462324 124456 462330
rect 124404 462266 124456 462272
rect 124864 452600 124916 452606
rect 124864 452542 124916 452548
rect 124312 399492 124364 399498
rect 124312 399434 124364 399440
rect 124220 354068 124272 354074
rect 124220 354010 124272 354016
rect 124232 353326 124260 354010
rect 124220 353320 124272 353326
rect 124220 353262 124272 353268
rect 124220 352572 124272 352578
rect 124220 352514 124272 352520
rect 124128 328432 124180 328438
rect 124128 328374 124180 328380
rect 124140 327826 124168 328374
rect 124128 327820 124180 327826
rect 124128 327762 124180 327768
rect 123668 305788 123720 305794
rect 123668 305730 123720 305736
rect 123576 294296 123628 294302
rect 123576 294238 123628 294244
rect 123484 291780 123536 291786
rect 123484 291722 123536 291728
rect 123484 289808 123536 289814
rect 123484 289750 123536 289756
rect 122378 289504 122434 289513
rect 122378 289439 122434 289448
rect 122392 288522 122420 289439
rect 123496 289134 123524 289750
rect 123484 289128 123536 289134
rect 123484 289070 123536 289076
rect 122380 288516 122432 288522
rect 122380 288458 122432 288464
rect 122748 286408 122800 286414
rect 122748 286350 122800 286356
rect 122760 285705 122788 286350
rect 122746 285696 122802 285705
rect 122746 285631 122802 285640
rect 122760 280838 122788 285631
rect 122748 280832 122800 280838
rect 122748 280774 122800 280780
rect 122286 255096 122342 255105
rect 122286 255031 122342 255040
rect 122102 251016 122158 251025
rect 122102 250951 122158 250960
rect 121550 250336 121606 250345
rect 121550 250271 121606 250280
rect 121564 249830 121592 250271
rect 122116 249898 122144 250951
rect 122104 249892 122156 249898
rect 122104 249834 122156 249840
rect 121552 249824 121604 249830
rect 121552 249766 121604 249772
rect 121550 248976 121606 248985
rect 121550 248911 121606 248920
rect 121564 248470 121592 248911
rect 121552 248464 121604 248470
rect 121552 248406 121604 248412
rect 121460 248396 121512 248402
rect 121460 248338 121512 248344
rect 121736 248396 121788 248402
rect 121736 248338 121788 248344
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121472 247178 121500 248231
rect 121642 247616 121698 247625
rect 121642 247551 121698 247560
rect 121460 247172 121512 247178
rect 121460 247114 121512 247120
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 121458 246256 121514 246265
rect 121458 246191 121514 246200
rect 121472 245682 121500 246191
rect 121564 245750 121592 246871
rect 121656 246362 121684 247551
rect 121644 246356 121696 246362
rect 121644 246298 121696 246304
rect 121552 245744 121604 245750
rect 121552 245686 121604 245692
rect 121460 245676 121512 245682
rect 121460 245618 121512 245624
rect 121642 245576 121698 245585
rect 121642 245511 121698 245520
rect 121550 244896 121606 244905
rect 121550 244831 121606 244840
rect 121458 244216 121514 244225
rect 121458 244151 121514 244160
rect 121472 243030 121500 244151
rect 121460 243024 121512 243030
rect 121460 242966 121512 242972
rect 121460 242888 121512 242894
rect 121458 242856 121460 242865
rect 121512 242856 121514 242865
rect 121564 242826 121592 244831
rect 121458 242791 121514 242800
rect 121552 242820 121604 242826
rect 121552 242762 121604 242768
rect 121366 241496 121422 241505
rect 121366 241431 121422 241440
rect 121458 240816 121514 240825
rect 121656 240786 121684 245511
rect 121748 243574 121776 248338
rect 122300 244934 122328 255031
rect 122288 244928 122340 244934
rect 122288 244870 122340 244876
rect 121736 243568 121788 243574
rect 121734 243536 121736 243545
rect 121788 243536 121790 243545
rect 121734 243471 121790 243480
rect 121458 240751 121514 240760
rect 121644 240780 121696 240786
rect 121472 240242 121500 240751
rect 121644 240722 121696 240728
rect 121460 240236 121512 240242
rect 121460 240178 121512 240184
rect 121458 240136 121514 240145
rect 121458 240071 121514 240080
rect 121472 238814 121500 240071
rect 121460 238808 121512 238814
rect 121460 238750 121512 238756
rect 123496 238678 123524 289070
rect 123588 265674 123616 294238
rect 123680 289814 123708 305730
rect 123760 294160 123812 294166
rect 123760 294102 123812 294108
rect 123668 289808 123720 289814
rect 123668 289750 123720 289756
rect 123772 278050 123800 294102
rect 123760 278044 123812 278050
rect 123760 277986 123812 277992
rect 123576 265668 123628 265674
rect 123576 265610 123628 265616
rect 124034 248296 124090 248305
rect 124034 248231 124090 248240
rect 124048 247110 124076 248231
rect 124036 247104 124088 247110
rect 124036 247046 124088 247052
rect 124232 239834 124260 352514
rect 124324 333946 124352 399434
rect 124404 387184 124456 387190
rect 124404 387126 124456 387132
rect 124416 338774 124444 387126
rect 124876 342242 124904 452542
rect 124968 444961 124996 541583
rect 125612 458182 125640 550598
rect 125704 492114 125732 583782
rect 127072 581120 127124 581126
rect 127072 581062 127124 581068
rect 125784 565956 125836 565962
rect 125784 565898 125836 565904
rect 125692 492108 125744 492114
rect 125692 492050 125744 492056
rect 125796 475998 125824 565898
rect 126980 497616 127032 497622
rect 126980 497558 127032 497564
rect 125876 494828 125928 494834
rect 125876 494770 125928 494776
rect 125784 475992 125836 475998
rect 125784 475934 125836 475940
rect 125600 458176 125652 458182
rect 125600 458118 125652 458124
rect 125598 453384 125654 453393
rect 125598 453319 125600 453328
rect 125652 453319 125654 453328
rect 125600 453290 125652 453296
rect 124954 444952 125010 444961
rect 124954 444887 125010 444896
rect 125784 438320 125836 438326
rect 125784 438262 125836 438268
rect 125692 396772 125744 396778
rect 125692 396714 125744 396720
rect 125600 353320 125652 353326
rect 125600 353262 125652 353268
rect 124864 342236 124916 342242
rect 124864 342178 124916 342184
rect 124864 341556 124916 341562
rect 124864 341498 124916 341504
rect 124404 338768 124456 338774
rect 124404 338710 124456 338716
rect 124312 333940 124364 333946
rect 124312 333882 124364 333888
rect 124402 316024 124458 316033
rect 124402 315959 124404 315968
rect 124456 315959 124458 315968
rect 124404 315930 124456 315936
rect 124312 310548 124364 310554
rect 124312 310490 124364 310496
rect 124324 274582 124352 310490
rect 124876 304298 124904 341498
rect 125508 311772 125560 311778
rect 125508 311714 125560 311720
rect 125520 310554 125548 311714
rect 125508 310548 125560 310554
rect 125508 310490 125560 310496
rect 124864 304292 124916 304298
rect 124864 304234 124916 304240
rect 124404 301504 124456 301510
rect 124404 301446 124456 301452
rect 124416 286822 124444 301446
rect 124864 291780 124916 291786
rect 124864 291722 124916 291728
rect 124404 286816 124456 286822
rect 124404 286758 124456 286764
rect 124416 286346 124444 286758
rect 124404 286340 124456 286346
rect 124404 286282 124456 286288
rect 124312 274576 124364 274582
rect 124312 274518 124364 274524
rect 124876 257378 124904 291722
rect 124956 283620 125008 283626
rect 124956 283562 125008 283568
rect 124968 273222 124996 283562
rect 124956 273216 125008 273222
rect 124956 273158 125008 273164
rect 124864 257372 124916 257378
rect 124864 257314 124916 257320
rect 124312 249892 124364 249898
rect 124312 249834 124364 249840
rect 124324 246430 124352 249834
rect 124312 246424 124364 246430
rect 124312 246366 124364 246372
rect 124220 239828 124272 239834
rect 124220 239770 124272 239776
rect 123484 238672 123536 238678
rect 123484 238614 123536 238620
rect 125612 235958 125640 353262
rect 125704 337482 125732 396714
rect 125796 337958 125824 438262
rect 125888 390726 125916 494770
rect 125968 462324 126020 462330
rect 125968 462266 126020 462272
rect 125876 390720 125928 390726
rect 125876 390662 125928 390668
rect 125980 352578 126008 462266
rect 126992 393990 127020 497558
rect 127084 491230 127112 581062
rect 127624 556232 127676 556238
rect 127624 556174 127676 556180
rect 127164 493468 127216 493474
rect 127164 493410 127216 493416
rect 127072 491224 127124 491230
rect 127072 491166 127124 491172
rect 127072 440360 127124 440366
rect 127072 440302 127124 440308
rect 126980 393984 127032 393990
rect 126980 393926 127032 393932
rect 126980 390652 127032 390658
rect 126980 390594 127032 390600
rect 125968 352572 126020 352578
rect 125968 352514 126020 352520
rect 126152 342916 126204 342922
rect 126152 342858 126204 342864
rect 126164 342417 126192 342858
rect 126150 342408 126206 342417
rect 126150 342343 126152 342352
rect 126204 342343 126206 342352
rect 126152 342314 126204 342320
rect 125784 337952 125836 337958
rect 125784 337894 125836 337900
rect 126888 337952 126940 337958
rect 126888 337894 126940 337900
rect 126900 337550 126928 337894
rect 126888 337544 126940 337550
rect 126888 337486 126940 337492
rect 125692 337476 125744 337482
rect 125692 337418 125744 337424
rect 125784 329860 125836 329866
rect 125784 329802 125836 329808
rect 125692 295724 125744 295730
rect 125692 295666 125744 295672
rect 125600 235952 125652 235958
rect 125600 235894 125652 235900
rect 120172 205012 120224 205018
rect 120172 204954 120224 204960
rect 125704 202162 125732 295666
rect 125796 286414 125824 329802
rect 126244 293412 126296 293418
rect 126244 293354 126296 293360
rect 125784 286408 125836 286414
rect 125784 286350 125836 286356
rect 126256 258738 126284 293354
rect 126244 258732 126296 258738
rect 126244 258674 126296 258680
rect 126992 231742 127020 390594
rect 127084 336734 127112 440302
rect 127176 395418 127204 493410
rect 127636 465118 127664 556174
rect 128360 534744 128412 534750
rect 128360 534686 128412 534692
rect 127624 465112 127676 465118
rect 127624 465054 127676 465060
rect 128372 437442 128400 534686
rect 128464 498846 128492 586502
rect 131120 585200 131172 585206
rect 131120 585142 131172 585148
rect 129832 584112 129884 584118
rect 129832 584054 129884 584060
rect 128636 572756 128688 572762
rect 128636 572698 128688 572704
rect 128544 537668 128596 537674
rect 128544 537610 128596 537616
rect 128452 498840 128504 498846
rect 128450 498808 128452 498817
rect 128504 498808 128506 498817
rect 128450 498743 128506 498752
rect 128452 487892 128504 487898
rect 128452 487834 128504 487840
rect 128360 437436 128412 437442
rect 128360 437378 128412 437384
rect 127256 403640 127308 403646
rect 127256 403582 127308 403588
rect 127164 395412 127216 395418
rect 127164 395354 127216 395360
rect 127072 336728 127124 336734
rect 127072 336670 127124 336676
rect 127268 313274 127296 403582
rect 128360 389292 128412 389298
rect 128360 389234 128412 389240
rect 127256 313268 127308 313274
rect 127256 313210 127308 313216
rect 127268 312497 127296 313210
rect 127254 312488 127310 312497
rect 127254 312423 127310 312432
rect 127624 304360 127676 304366
rect 127624 304302 127676 304308
rect 127636 242962 127664 304302
rect 127624 242956 127676 242962
rect 127624 242898 127676 242904
rect 127636 238513 127664 242898
rect 127622 238504 127678 238513
rect 127622 238439 127678 238448
rect 126980 231736 127032 231742
rect 126980 231678 127032 231684
rect 127440 231736 127492 231742
rect 127440 231678 127492 231684
rect 127452 231130 127480 231678
rect 127440 231124 127492 231130
rect 127440 231066 127492 231072
rect 128372 229022 128400 389234
rect 128464 385014 128492 487834
rect 128556 445058 128584 537610
rect 128648 481642 128676 572698
rect 129844 493338 129872 584054
rect 130016 561740 130068 561746
rect 130016 561682 130068 561688
rect 129924 538892 129976 538898
rect 129924 538834 129976 538840
rect 129832 493332 129884 493338
rect 129832 493274 129884 493280
rect 128636 481636 128688 481642
rect 128636 481578 128688 481584
rect 128648 480962 128676 481578
rect 128636 480956 128688 480962
rect 128636 480898 128688 480904
rect 129740 471980 129792 471986
rect 129740 471922 129792 471928
rect 128544 445052 128596 445058
rect 128544 444994 128596 445000
rect 128636 403708 128688 403714
rect 128636 403650 128688 403656
rect 128544 389360 128596 389366
rect 128544 389302 128596 389308
rect 128452 385008 128504 385014
rect 128452 384950 128504 384956
rect 128452 342372 128504 342378
rect 128452 342314 128504 342320
rect 128464 238649 128492 342314
rect 128556 298790 128584 389302
rect 128648 341630 128676 403650
rect 129752 365702 129780 471922
rect 129936 438938 129964 538834
rect 130028 470558 130056 561682
rect 131132 496126 131160 585142
rect 131212 499588 131264 499594
rect 131212 499530 131264 499536
rect 131120 496120 131172 496126
rect 131120 496062 131172 496068
rect 130108 494760 130160 494766
rect 130108 494702 130160 494708
rect 130016 470552 130068 470558
rect 130016 470494 130068 470500
rect 130028 469946 130056 470494
rect 130016 469940 130068 469946
rect 130016 469882 130068 469888
rect 129924 438932 129976 438938
rect 129924 438874 129976 438880
rect 129924 438252 129976 438258
rect 129924 438194 129976 438200
rect 129830 388376 129886 388385
rect 129830 388311 129886 388320
rect 129740 365696 129792 365702
rect 129740 365638 129792 365644
rect 128636 341624 128688 341630
rect 128636 341566 128688 341572
rect 129740 334008 129792 334014
rect 129740 333950 129792 333956
rect 128636 316804 128688 316810
rect 128636 316746 128688 316752
rect 128544 298784 128596 298790
rect 128544 298726 128596 298732
rect 128544 286816 128596 286822
rect 128544 286758 128596 286764
rect 128556 282198 128584 286758
rect 128544 282192 128596 282198
rect 128544 282134 128596 282140
rect 128648 263498 128676 316746
rect 129752 287054 129780 333950
rect 129844 312594 129872 388311
rect 129936 335306 129964 438194
rect 130016 402280 130068 402286
rect 130016 402222 130068 402228
rect 129924 335300 129976 335306
rect 129924 335242 129976 335248
rect 129936 334014 129964 335242
rect 129924 334008 129976 334014
rect 129924 333950 129976 333956
rect 130028 328370 130056 402222
rect 130120 389842 130148 494702
rect 131224 396846 131252 499530
rect 131316 491978 131344 586706
rect 133144 578332 133196 578338
rect 133144 578274 133196 578280
rect 132592 546508 132644 546514
rect 132592 546450 132644 546456
rect 131396 497480 131448 497486
rect 131396 497422 131448 497428
rect 131304 491972 131356 491978
rect 131304 491914 131356 491920
rect 131304 400920 131356 400926
rect 131304 400862 131356 400868
rect 131212 396840 131264 396846
rect 131212 396782 131264 396788
rect 131212 391332 131264 391338
rect 131212 391274 131264 391280
rect 130384 389904 130436 389910
rect 130384 389846 130436 389852
rect 130108 389836 130160 389842
rect 130108 389778 130160 389784
rect 130396 388385 130424 389846
rect 130382 388376 130438 388385
rect 130382 388311 130438 388320
rect 131120 369164 131172 369170
rect 131120 369106 131172 369112
rect 130016 328364 130068 328370
rect 130016 328306 130068 328312
rect 130384 328364 130436 328370
rect 130384 328306 130436 328312
rect 130396 327758 130424 328306
rect 130384 327752 130436 327758
rect 130384 327694 130436 327700
rect 129832 312588 129884 312594
rect 129832 312530 129884 312536
rect 130384 299736 130436 299742
rect 130384 299678 130436 299684
rect 129752 287026 129872 287054
rect 129844 273154 129872 287026
rect 129832 273148 129884 273154
rect 129832 273090 129884 273096
rect 129844 272610 129872 273090
rect 129832 272604 129884 272610
rect 129832 272546 129884 272552
rect 129648 268456 129700 268462
rect 129648 268398 129700 268404
rect 129660 267850 129688 268398
rect 129648 267844 129700 267850
rect 129648 267786 129700 267792
rect 128636 263492 128688 263498
rect 128636 263434 128688 263440
rect 128912 263492 128964 263498
rect 128912 263434 128964 263440
rect 128924 262954 128952 263434
rect 128912 262948 128964 262954
rect 128912 262890 128964 262896
rect 129660 250510 129688 267786
rect 129648 250504 129700 250510
rect 129648 250446 129700 250452
rect 128450 238640 128506 238649
rect 128450 238575 128506 238584
rect 128360 229016 128412 229022
rect 128360 228958 128412 228964
rect 128372 228410 128400 228958
rect 128360 228404 128412 228410
rect 128360 228346 128412 228352
rect 125692 202156 125744 202162
rect 125692 202098 125744 202104
rect 119344 191140 119396 191146
rect 119344 191082 119396 191088
rect 116584 189780 116636 189786
rect 116584 189722 116636 189728
rect 130396 188494 130424 299678
rect 131132 297401 131160 369106
rect 131224 339590 131252 391274
rect 131212 339584 131264 339590
rect 131212 339526 131264 339532
rect 131316 320142 131344 400862
rect 131408 392698 131436 497422
rect 132500 494896 132552 494902
rect 132500 494838 132552 494844
rect 131764 475992 131816 475998
rect 131764 475934 131816 475940
rect 131396 392692 131448 392698
rect 131396 392634 131448 392640
rect 131776 368558 131804 475934
rect 132512 386510 132540 494838
rect 132604 455462 132632 546450
rect 132684 537532 132736 537538
rect 132684 537474 132736 537480
rect 132592 455456 132644 455462
rect 132592 455398 132644 455404
rect 132500 386504 132552 386510
rect 132500 386446 132552 386452
rect 131396 368552 131448 368558
rect 131396 368494 131448 368500
rect 131764 368552 131816 368558
rect 131764 368494 131816 368500
rect 131408 368422 131436 368494
rect 131396 368416 131448 368422
rect 131396 368358 131448 368364
rect 131396 356720 131448 356726
rect 131396 356662 131448 356668
rect 131408 356182 131436 356662
rect 131396 356176 131448 356182
rect 131396 356118 131448 356124
rect 131764 356176 131816 356182
rect 131764 356118 131816 356124
rect 131304 320136 131356 320142
rect 131304 320078 131356 320084
rect 131672 320136 131724 320142
rect 131672 320078 131724 320084
rect 131684 319433 131712 320078
rect 131670 319424 131726 319433
rect 131670 319359 131726 319368
rect 131118 297392 131174 297401
rect 131118 297327 131174 297336
rect 131120 293344 131172 293350
rect 131120 293286 131172 293292
rect 131132 276010 131160 293286
rect 131120 276004 131172 276010
rect 131120 275946 131172 275952
rect 131132 275330 131160 275946
rect 131120 275324 131172 275330
rect 131120 275266 131172 275272
rect 131776 227730 131804 356118
rect 132512 237250 132540 386446
rect 132604 346390 132632 455398
rect 132696 440366 132724 537474
rect 133156 487830 133184 578274
rect 135260 578264 135312 578270
rect 135260 578206 135312 578212
rect 133880 564460 133932 564466
rect 133880 564402 133932 564408
rect 133144 487824 133196 487830
rect 133144 487766 133196 487772
rect 133892 472666 133920 564402
rect 134248 545148 134300 545154
rect 134248 545090 134300 545096
rect 134156 542428 134208 542434
rect 134156 542370 134208 542376
rect 133880 472660 133932 472666
rect 133880 472602 133932 472608
rect 133892 470594 133920 472602
rect 133892 470566 134104 470594
rect 133972 459604 134024 459610
rect 133972 459546 134024 459552
rect 132868 441652 132920 441658
rect 132868 441594 132920 441600
rect 132684 440360 132736 440366
rect 132684 440302 132736 440308
rect 132776 401056 132828 401062
rect 132776 400998 132828 401004
rect 132592 346384 132644 346390
rect 132592 346326 132644 346332
rect 132788 335354 132816 400998
rect 132880 339454 132908 441594
rect 133880 440292 133932 440298
rect 133880 440234 133932 440240
rect 133788 346384 133840 346390
rect 133788 346326 133840 346332
rect 133800 345710 133828 346326
rect 133788 345704 133840 345710
rect 133788 345646 133840 345652
rect 132868 339448 132920 339454
rect 132868 339390 132920 339396
rect 132696 335326 132816 335354
rect 132696 325650 132724 335326
rect 132684 325644 132736 325650
rect 132684 325586 132736 325592
rect 133788 325644 133840 325650
rect 133788 325586 133840 325592
rect 133800 324970 133828 325586
rect 133788 324964 133840 324970
rect 133788 324906 133840 324912
rect 133892 321570 133920 440234
rect 133984 349858 134012 459546
rect 134076 367062 134104 470566
rect 134168 451926 134196 542370
rect 134260 454714 134288 545090
rect 135272 487150 135300 578206
rect 137284 574116 137336 574122
rect 137284 574058 137336 574064
rect 136824 559564 136876 559570
rect 136824 559506 136876 559512
rect 136836 558958 136864 559506
rect 136824 558952 136876 558958
rect 136824 558894 136876 558900
rect 135444 549364 135496 549370
rect 135444 549306 135496 549312
rect 135260 487144 135312 487150
rect 135260 487086 135312 487092
rect 135352 486464 135404 486470
rect 135352 486406 135404 486412
rect 134248 454708 134300 454714
rect 134248 454650 134300 454656
rect 134156 451920 134208 451926
rect 134156 451862 134208 451868
rect 135260 438184 135312 438190
rect 135260 438126 135312 438132
rect 134522 385656 134578 385665
rect 134522 385591 134578 385600
rect 134064 367056 134116 367062
rect 134064 366998 134116 367004
rect 134064 360324 134116 360330
rect 134064 360266 134116 360272
rect 133972 349852 134024 349858
rect 133972 349794 134024 349800
rect 133984 341562 134012 349794
rect 133972 341556 134024 341562
rect 133972 341498 134024 341504
rect 133880 321564 133932 321570
rect 133880 321506 133932 321512
rect 133144 297084 133196 297090
rect 133144 297026 133196 297032
rect 132500 237244 132552 237250
rect 132500 237186 132552 237192
rect 131212 227724 131264 227730
rect 131212 227666 131264 227672
rect 131764 227724 131816 227730
rect 131764 227666 131816 227672
rect 131224 227050 131252 227666
rect 131212 227044 131264 227050
rect 131212 226986 131264 226992
rect 133156 199714 133184 297026
rect 133878 296984 133934 296993
rect 133878 296919 133934 296928
rect 133144 199708 133196 199714
rect 133144 199650 133196 199656
rect 130384 188488 130436 188494
rect 130384 188430 130436 188436
rect 133144 186380 133196 186386
rect 133144 186322 133196 186328
rect 124128 185020 124180 185026
rect 124128 184962 124180 184968
rect 121368 183592 121420 183598
rect 121368 183534 121420 183540
rect 118516 181008 118568 181014
rect 118516 180950 118568 180956
rect 114376 180940 114428 180946
rect 114376 180882 114428 180888
rect 114008 179580 114060 179586
rect 114008 179522 114060 179528
rect 114020 177041 114048 179522
rect 114388 177721 114416 180882
rect 115848 179512 115900 179518
rect 115848 179454 115900 179460
rect 114374 177712 114430 177721
rect 114374 177647 114430 177656
rect 115860 177041 115888 179454
rect 118528 177721 118556 180950
rect 119528 178016 119580 178022
rect 119528 177958 119580 177964
rect 118514 177712 118570 177721
rect 118514 177647 118570 177656
rect 114006 177032 114062 177041
rect 114006 176967 114062 176976
rect 115846 177032 115902 177041
rect 115846 176967 115902 176976
rect 119540 176769 119568 177958
rect 121380 177721 121408 183534
rect 121458 179480 121514 179489
rect 121458 179415 121514 179424
rect 121472 177954 121500 179415
rect 122104 178084 122156 178090
rect 122104 178026 122156 178032
rect 121460 177948 121512 177954
rect 121460 177890 121512 177896
rect 121366 177712 121422 177721
rect 121366 177647 121422 177656
rect 122116 176769 122144 178026
rect 124140 177177 124168 184962
rect 126888 184952 126940 184958
rect 126888 184894 126940 184900
rect 126900 177721 126928 184894
rect 130752 182300 130804 182306
rect 130752 182242 130804 182248
rect 127900 177948 127952 177954
rect 127900 177890 127952 177896
rect 126886 177712 126942 177721
rect 126886 177647 126942 177656
rect 124126 177168 124182 177177
rect 124126 177103 124182 177112
rect 124496 176996 124548 177002
rect 124496 176938 124548 176944
rect 124508 176769 124536 176938
rect 127912 176769 127940 177890
rect 130764 177721 130792 182242
rect 132408 181076 132460 181082
rect 132408 181018 132460 181024
rect 132420 177721 132448 181018
rect 133156 177954 133184 186322
rect 133892 178702 133920 296919
rect 134076 287026 134104 360266
rect 134536 309942 134564 385591
rect 134616 334688 134668 334694
rect 134616 334630 134668 334636
rect 134524 309936 134576 309942
rect 134524 309878 134576 309884
rect 134064 287020 134116 287026
rect 134064 286962 134116 286968
rect 134076 286346 134104 286962
rect 134064 286340 134116 286346
rect 134064 286282 134116 286288
rect 134628 260914 134656 334630
rect 135272 329798 135300 438126
rect 135364 381546 135392 486406
rect 135456 458862 135484 549306
rect 136732 487824 136784 487830
rect 136732 487766 136784 487772
rect 136548 487144 136600 487150
rect 136548 487086 136600 487092
rect 136560 486538 136588 487086
rect 136548 486532 136600 486538
rect 136548 486474 136600 486480
rect 136640 478916 136692 478922
rect 136640 478858 136692 478864
rect 135444 458856 135496 458862
rect 135444 458798 135496 458804
rect 135456 458250 135484 458798
rect 135444 458244 135496 458250
rect 135444 458186 135496 458192
rect 135444 394052 135496 394058
rect 135444 393994 135496 394000
rect 135352 381540 135404 381546
rect 135352 381482 135404 381488
rect 135260 329792 135312 329798
rect 135260 329734 135312 329740
rect 135168 321564 135220 321570
rect 135168 321506 135220 321512
rect 135180 320890 135208 321506
rect 135168 320884 135220 320890
rect 135168 320826 135220 320832
rect 135168 309936 135220 309942
rect 135168 309878 135220 309884
rect 135180 309806 135208 309878
rect 135168 309800 135220 309806
rect 135168 309742 135220 309748
rect 135364 292534 135392 381482
rect 135456 311846 135484 393994
rect 136652 373994 136680 478858
rect 136744 383654 136772 487766
rect 136836 466410 136864 558894
rect 137296 483070 137324 574058
rect 159376 574054 159404 683130
rect 162136 585818 162164 700334
rect 170324 697610 170352 703520
rect 202800 703390 202828 703520
rect 201500 703384 201552 703390
rect 201500 703326 201552 703332
rect 202788 703384 202840 703390
rect 202788 703326 202840 703332
rect 170312 697604 170364 697610
rect 170312 697546 170364 697552
rect 162124 585812 162176 585818
rect 162124 585754 162176 585760
rect 159364 574048 159416 574054
rect 159364 573990 159416 573996
rect 140780 571396 140832 571402
rect 140780 571338 140832 571344
rect 138112 560380 138164 560386
rect 138112 560322 138164 560328
rect 138020 552084 138072 552090
rect 138020 552026 138072 552032
rect 137284 483064 137336 483070
rect 137284 483006 137336 483012
rect 136824 466404 136876 466410
rect 136824 466346 136876 466352
rect 138032 459542 138060 552026
rect 138124 469878 138152 560322
rect 139492 560312 139544 560318
rect 139492 560254 139544 560260
rect 139400 493332 139452 493338
rect 139400 493274 139452 493280
rect 138112 469872 138164 469878
rect 138112 469814 138164 469820
rect 138112 465112 138164 465118
rect 138112 465054 138164 465060
rect 138020 459536 138072 459542
rect 138020 459478 138072 459484
rect 136824 398268 136876 398274
rect 136824 398210 136876 398216
rect 136732 383648 136784 383654
rect 136732 383590 136784 383596
rect 136744 382974 136772 383590
rect 136732 382968 136784 382974
rect 136732 382910 136784 382916
rect 136652 373966 136772 373994
rect 136744 370530 136772 373966
rect 136732 370524 136784 370530
rect 136732 370466 136784 370472
rect 136640 367056 136692 367062
rect 136640 366998 136692 367004
rect 136548 329792 136600 329798
rect 136548 329734 136600 329740
rect 136560 329118 136588 329734
rect 136548 329112 136600 329118
rect 136548 329054 136600 329060
rect 135444 311840 135496 311846
rect 135444 311782 135496 311788
rect 136548 311840 136600 311846
rect 136548 311782 136600 311788
rect 136560 311234 136588 311782
rect 136548 311228 136600 311234
rect 136548 311170 136600 311176
rect 135904 302524 135956 302530
rect 135904 302466 135956 302472
rect 135352 292528 135404 292534
rect 135352 292470 135404 292476
rect 134616 260908 134668 260914
rect 134616 260850 134668 260856
rect 134892 260908 134944 260914
rect 134892 260850 134944 260856
rect 134904 259418 134932 260850
rect 134892 259412 134944 259418
rect 134892 259354 134944 259360
rect 135916 245002 135944 302466
rect 135904 244996 135956 245002
rect 135904 244938 135956 244944
rect 136652 226273 136680 366998
rect 136744 366382 136772 370466
rect 136732 366376 136784 366382
rect 136732 366318 136784 366324
rect 136836 327078 136864 398210
rect 138020 392080 138072 392086
rect 138020 392022 138072 392028
rect 137284 390584 137336 390590
rect 136914 390552 136970 390561
rect 137284 390526 137336 390532
rect 136914 390487 136970 390496
rect 136928 389230 136956 390487
rect 136916 389224 136968 389230
rect 136916 389166 136968 389172
rect 136824 327072 136876 327078
rect 136824 327014 136876 327020
rect 137100 327072 137152 327078
rect 137100 327014 137152 327020
rect 137112 326505 137140 327014
rect 137098 326496 137154 326505
rect 137098 326431 137154 326440
rect 137296 263634 137324 390526
rect 137284 263628 137336 263634
rect 137284 263570 137336 263576
rect 137296 262206 137324 263570
rect 137284 262200 137336 262206
rect 137284 262142 137336 262148
rect 136638 226264 136694 226273
rect 136638 226199 136694 226208
rect 136652 225729 136680 226199
rect 136638 225720 136694 225729
rect 136638 225655 136694 225664
rect 138032 208350 138060 392022
rect 138124 356726 138152 465054
rect 138204 445800 138256 445806
rect 138204 445742 138256 445748
rect 138112 356720 138164 356726
rect 138112 356662 138164 356668
rect 138216 345014 138244 445742
rect 139412 389910 139440 493274
rect 139504 471306 139532 560254
rect 139584 549296 139636 549302
rect 139584 549238 139636 549244
rect 139492 471300 139544 471306
rect 139492 471242 139544 471248
rect 139504 470626 139532 471242
rect 139492 470620 139544 470626
rect 139492 470562 139544 470568
rect 139492 458244 139544 458250
rect 139492 458186 139544 458192
rect 139400 389904 139452 389910
rect 139400 389846 139452 389852
rect 139504 349110 139532 458186
rect 139596 456754 139624 549238
rect 140792 480214 140820 571338
rect 142160 569968 142212 569974
rect 142160 569910 142212 569916
rect 141516 554056 141568 554062
rect 141516 553998 141568 554004
rect 141528 553450 141556 553998
rect 140964 553444 141016 553450
rect 140964 553386 141016 553392
rect 141516 553444 141568 553450
rect 141516 553386 141568 553392
rect 140872 543788 140924 543794
rect 140872 543730 140924 543736
rect 140780 480208 140832 480214
rect 140780 480150 140832 480156
rect 140792 479534 140820 480150
rect 140780 479528 140832 479534
rect 140780 479470 140832 479476
rect 139584 456748 139636 456754
rect 139584 456690 139636 456696
rect 140320 456748 140372 456754
rect 140320 456690 140372 456696
rect 140332 456074 140360 456690
rect 140320 456068 140372 456074
rect 140320 456010 140372 456016
rect 140780 449948 140832 449954
rect 140780 449890 140832 449896
rect 139584 392692 139636 392698
rect 139584 392634 139636 392640
rect 139492 349104 139544 349110
rect 139492 349046 139544 349052
rect 138124 344986 138244 345014
rect 138124 338094 138152 344986
rect 138112 338088 138164 338094
rect 138112 338030 138164 338036
rect 138124 337482 138152 338030
rect 138112 337476 138164 337482
rect 138112 337418 138164 337424
rect 139596 268462 139624 392634
rect 139768 349104 139820 349110
rect 139768 349046 139820 349052
rect 139780 348430 139808 349046
rect 139768 348424 139820 348430
rect 139768 348366 139820 348372
rect 140792 338026 140820 449890
rect 140884 431866 140912 543730
rect 140976 462398 141004 553386
rect 141056 496120 141108 496126
rect 141056 496062 141108 496068
rect 140964 462392 141016 462398
rect 140964 462334 141016 462340
rect 140872 431860 140924 431866
rect 140872 431802 140924 431808
rect 140884 431254 140912 431802
rect 140872 431248 140924 431254
rect 140872 431190 140924 431196
rect 140872 398200 140924 398206
rect 140872 398142 140924 398148
rect 140884 345030 140912 398142
rect 140976 354686 141004 462334
rect 141068 388482 141096 496062
rect 142172 476066 142200 569910
rect 142252 565888 142304 565894
rect 142252 565830 142304 565836
rect 142160 476060 142212 476066
rect 142160 476002 142212 476008
rect 142264 474706 142292 565830
rect 201512 559570 201540 703326
rect 218992 700398 219020 703520
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 235184 700330 235212 703520
rect 267660 703322 267688 703520
rect 267648 703316 267700 703322
rect 267648 703258 267700 703264
rect 283852 700330 283880 703520
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 238024 700324 238076 700330
rect 238024 700266 238076 700272
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 238036 596834 238064 700266
rect 238024 596828 238076 596834
rect 238024 596770 238076 596776
rect 204904 564460 204956 564466
rect 204904 564402 204956 564408
rect 201500 559564 201552 559570
rect 201500 559506 201552 559512
rect 142436 539640 142488 539646
rect 142436 539582 142488 539588
rect 142252 474700 142304 474706
rect 142252 474642 142304 474648
rect 142344 470620 142396 470626
rect 142344 470562 142396 470568
rect 142252 469872 142304 469878
rect 142252 469814 142304 469820
rect 142160 445052 142212 445058
rect 142160 444994 142212 445000
rect 141056 388476 141108 388482
rect 141056 388418 141108 388424
rect 141792 361548 141844 361554
rect 141792 361490 141844 361496
rect 141804 360262 141832 361490
rect 141424 360256 141476 360262
rect 141424 360198 141476 360204
rect 141792 360256 141844 360262
rect 141792 360198 141844 360204
rect 140964 354680 141016 354686
rect 140964 354622 141016 354628
rect 140976 353326 141004 354622
rect 140964 353320 141016 353326
rect 140964 353262 141016 353268
rect 140872 345024 140924 345030
rect 140872 344966 140924 344972
rect 140884 344350 140912 344966
rect 140872 344344 140924 344350
rect 140872 344286 140924 344292
rect 140872 342304 140924 342310
rect 140872 342246 140924 342252
rect 140780 338020 140832 338026
rect 140780 337962 140832 337968
rect 140780 337544 140832 337550
rect 140780 337486 140832 337492
rect 139584 268456 139636 268462
rect 139584 268398 139636 268404
rect 140792 263566 140820 337486
rect 140780 263560 140832 263566
rect 140780 263502 140832 263508
rect 140792 262886 140820 263502
rect 140780 262880 140832 262886
rect 140780 262822 140832 262828
rect 140884 248414 140912 342246
rect 141436 311166 141464 360198
rect 141424 311160 141476 311166
rect 141424 311102 141476 311108
rect 142172 309126 142200 444994
rect 142264 361554 142292 469814
rect 142356 362234 142384 470562
rect 142448 449206 142476 539582
rect 204916 538218 204944 564402
rect 299492 541657 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703254 332548 703520
rect 332508 703248 332560 703254
rect 332508 703190 332560 703196
rect 348804 703186 348832 703520
rect 348792 703180 348844 703186
rect 348792 703122 348844 703128
rect 364996 703050 365024 703520
rect 397472 703118 397500 703520
rect 397460 703112 397512 703118
rect 397460 703054 397512 703060
rect 364984 703044 365036 703050
rect 364984 702986 365036 702992
rect 364996 701758 365024 702986
rect 413664 702982 413692 703520
rect 413652 702976 413704 702982
rect 413652 702918 413704 702924
rect 429856 702846 429884 703520
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 429200 702840 429252 702846
rect 429200 702782 429252 702788
rect 429844 702840 429896 702846
rect 429844 702782 429896 702788
rect 364984 701752 365036 701758
rect 364984 701694 365036 701700
rect 425704 616140 425756 616146
rect 425704 616082 425756 616088
rect 299478 541648 299534 541657
rect 299478 541583 299534 541592
rect 425716 539578 425744 616082
rect 425060 539572 425112 539578
rect 425060 539514 425112 539520
rect 425704 539572 425756 539578
rect 425704 539514 425756 539520
rect 425072 538286 425100 539514
rect 425060 538280 425112 538286
rect 425060 538222 425112 538228
rect 204904 538212 204956 538218
rect 204904 538154 204956 538160
rect 420920 534744 420972 534750
rect 420920 534686 420972 534692
rect 143540 491972 143592 491978
rect 143540 491914 143592 491920
rect 142436 449200 142488 449206
rect 142436 449142 142488 449148
rect 142436 389836 142488 389842
rect 142436 389778 142488 389784
rect 142344 362228 142396 362234
rect 142344 362170 142396 362176
rect 142252 361548 142304 361554
rect 142252 361490 142304 361496
rect 142252 353320 142304 353326
rect 142252 353262 142304 353268
rect 142160 309120 142212 309126
rect 142160 309062 142212 309068
rect 140792 248386 140912 248414
rect 140792 242826 140820 248386
rect 140780 242820 140832 242826
rect 140780 242762 140832 242768
rect 140792 242214 140820 242762
rect 140780 242208 140832 242214
rect 140780 242150 140832 242156
rect 142264 224942 142292 353262
rect 142448 288386 142476 389778
rect 143552 385665 143580 491914
rect 150532 486532 150584 486538
rect 150532 486474 150584 486480
rect 147956 483064 148008 483070
rect 147956 483006 148008 483012
rect 146300 480956 146352 480962
rect 146300 480898 146352 480904
rect 145012 479528 145064 479534
rect 145012 479470 145064 479476
rect 143724 454708 143776 454714
rect 143724 454650 143776 454656
rect 143538 385656 143594 385665
rect 143538 385591 143594 385600
rect 143632 376780 143684 376786
rect 143632 376722 143684 376728
rect 143540 358080 143592 358086
rect 143540 358022 143592 358028
rect 143448 309120 143500 309126
rect 143448 309062 143500 309068
rect 143460 308446 143488 309062
rect 143448 308440 143500 308446
rect 143448 308382 143500 308388
rect 142804 292732 142856 292738
rect 142804 292674 142856 292680
rect 142436 288380 142488 288386
rect 142436 288322 142488 288328
rect 142252 224936 142304 224942
rect 142252 224878 142304 224884
rect 138020 208344 138072 208350
rect 138020 208286 138072 208292
rect 138032 207670 138060 208286
rect 138020 207664 138072 207670
rect 138020 207606 138072 207612
rect 135904 187740 135956 187746
rect 135904 187682 135956 187688
rect 133880 178696 133932 178702
rect 133880 178638 133932 178644
rect 135916 178022 135944 187682
rect 142816 183054 142844 292674
rect 143448 288380 143500 288386
rect 143448 288322 143500 288328
rect 143460 287706 143488 288322
rect 143448 287700 143500 287706
rect 143448 287642 143500 287648
rect 143448 224936 143500 224942
rect 143448 224878 143500 224884
rect 143460 224262 143488 224878
rect 143448 224256 143500 224262
rect 143448 224198 143500 224204
rect 143552 205630 143580 358022
rect 143644 267734 143672 376722
rect 143736 343602 143764 454650
rect 143816 449200 143868 449206
rect 143816 449142 143868 449148
rect 143724 343596 143776 343602
rect 143724 343538 143776 343544
rect 143828 339522 143856 449142
rect 144918 448624 144974 448633
rect 144918 448559 144974 448568
rect 144828 343596 144880 343602
rect 144828 343538 144880 343544
rect 144840 342922 144868 343538
rect 144828 342916 144880 342922
rect 144828 342858 144880 342864
rect 143816 339516 143868 339522
rect 143816 339458 143868 339464
rect 144932 332586 144960 448559
rect 145024 375358 145052 479470
rect 145104 382968 145156 382974
rect 145104 382910 145156 382916
rect 145012 375352 145064 375358
rect 145012 375294 145064 375300
rect 144920 332580 144972 332586
rect 144920 332522 144972 332528
rect 145116 301510 145144 382910
rect 146312 376718 146340 480898
rect 146392 471368 146444 471374
rect 146392 471310 146444 471316
rect 146404 470626 146432 471310
rect 146392 470620 146444 470626
rect 146392 470562 146444 470568
rect 146300 376712 146352 376718
rect 146300 376654 146352 376660
rect 146208 375352 146260 375358
rect 146208 375294 146260 375300
rect 146220 374649 146248 375294
rect 146206 374640 146262 374649
rect 146206 374575 146262 374584
rect 146300 368552 146352 368558
rect 146300 368494 146352 368500
rect 146208 332580 146260 332586
rect 146208 332522 146260 332528
rect 146220 331906 146248 332522
rect 146208 331900 146260 331906
rect 146208 331842 146260 331848
rect 145104 301504 145156 301510
rect 145104 301446 145156 301452
rect 144184 295656 144236 295662
rect 144184 295598 144236 295604
rect 144196 283529 144224 295598
rect 144182 283520 144238 283529
rect 144182 283455 144238 283464
rect 143644 267706 143764 267734
rect 143736 252550 143764 267706
rect 146312 260846 146340 368494
rect 146404 365090 146432 470562
rect 147864 460964 147916 460970
rect 147864 460906 147916 460912
rect 147772 451920 147824 451926
rect 147772 451862 147824 451868
rect 146944 396092 146996 396098
rect 146944 396034 146996 396040
rect 146392 365084 146444 365090
rect 146392 365026 146444 365032
rect 146956 303958 146984 396034
rect 147680 393372 147732 393378
rect 147680 393314 147732 393320
rect 146944 303952 146996 303958
rect 146944 303894 146996 303900
rect 146956 294710 146984 303894
rect 147036 298444 147088 298450
rect 147036 298386 147088 298392
rect 146944 294704 146996 294710
rect 146944 294646 146996 294652
rect 146300 260840 146352 260846
rect 146300 260782 146352 260788
rect 146760 260840 146812 260846
rect 146760 260782 146812 260788
rect 146772 260166 146800 260782
rect 146760 260160 146812 260166
rect 146760 260102 146812 260108
rect 143724 252544 143776 252550
rect 143724 252486 143776 252492
rect 144828 252544 144880 252550
rect 144828 252486 144880 252492
rect 144840 251870 144868 252486
rect 144828 251864 144880 251870
rect 144828 251806 144880 251812
rect 143540 205624 143592 205630
rect 143540 205566 143592 205572
rect 144828 205624 144880 205630
rect 144828 205566 144880 205572
rect 144840 205018 144868 205566
rect 144828 205012 144880 205018
rect 144828 204954 144880 204960
rect 147048 193905 147076 298386
rect 147692 242894 147720 393314
rect 147784 340202 147812 451862
rect 147876 351898 147904 460906
rect 147968 378146 147996 483006
rect 149152 456068 149204 456074
rect 149152 456010 149204 456016
rect 147956 378140 148008 378146
rect 147956 378082 148008 378088
rect 147968 377466 147996 378082
rect 147956 377460 148008 377466
rect 147956 377402 148008 377408
rect 149060 376712 149112 376718
rect 149060 376654 149112 376660
rect 147864 351892 147916 351898
rect 147864 351834 147916 351840
rect 147876 351218 147904 351834
rect 147864 351212 147916 351218
rect 147864 351154 147916 351160
rect 147772 340196 147824 340202
rect 147772 340138 147824 340144
rect 147772 322312 147824 322318
rect 147772 322254 147824 322260
rect 147680 242888 147732 242894
rect 147680 242830 147732 242836
rect 147784 215286 147812 322254
rect 149072 229090 149100 376654
rect 149164 347750 149192 456010
rect 150440 393440 150492 393446
rect 150440 393382 150492 393388
rect 149152 347744 149204 347750
rect 149152 347686 149204 347692
rect 149704 347744 149756 347750
rect 149704 347686 149756 347692
rect 149716 347138 149744 347686
rect 149704 347132 149756 347138
rect 149704 347074 149756 347080
rect 150452 273222 150480 393382
rect 150544 368393 150572 486474
rect 151820 476808 151872 476814
rect 151820 476750 151872 476756
rect 150624 474700 150676 474706
rect 150624 474642 150676 474648
rect 150636 368490 150664 474642
rect 150716 431248 150768 431254
rect 150716 431190 150768 431196
rect 150624 368484 150676 368490
rect 150624 368426 150676 368432
rect 150530 368384 150586 368393
rect 150530 368319 150586 368328
rect 150728 340270 150756 431190
rect 151832 373998 151860 476750
rect 152004 469940 152056 469946
rect 152004 469882 152056 469888
rect 151912 456816 151964 456822
rect 151912 456758 151964 456764
rect 151820 373992 151872 373998
rect 151820 373934 151872 373940
rect 151832 373289 151860 373934
rect 151818 373280 151874 373289
rect 151818 373215 151874 373224
rect 151820 369912 151872 369918
rect 151820 369854 151872 369860
rect 151176 368484 151228 368490
rect 151176 368426 151228 368432
rect 150990 368384 151046 368393
rect 150990 368319 151046 368328
rect 151004 367713 151032 368319
rect 151188 367742 151216 368426
rect 151176 367736 151228 367742
rect 150990 367704 151046 367713
rect 151176 367678 151228 367684
rect 150990 367639 151046 367648
rect 150716 340264 150768 340270
rect 150716 340206 150768 340212
rect 150728 335354 150756 340206
rect 150544 335326 150756 335354
rect 150440 273216 150492 273222
rect 150440 273158 150492 273164
rect 150452 272542 150480 273158
rect 150440 272536 150492 272542
rect 150440 272478 150492 272484
rect 150544 237386 150572 335326
rect 150532 237380 150584 237386
rect 150532 237322 150584 237328
rect 150544 236706 150572 237322
rect 150532 236700 150584 236706
rect 150532 236642 150584 236648
rect 149060 229084 149112 229090
rect 149060 229026 149112 229032
rect 149072 228614 149100 229026
rect 149060 228608 149112 228614
rect 149060 228550 149112 228556
rect 151084 224392 151136 224398
rect 151084 224334 151136 224340
rect 147772 215280 147824 215286
rect 147772 215222 147824 215228
rect 147784 214674 147812 215222
rect 147772 214668 147824 214674
rect 147772 214610 147824 214616
rect 147034 193896 147090 193905
rect 147034 193831 147090 193840
rect 151096 185774 151124 224334
rect 151832 216646 151860 369854
rect 151924 345778 151952 456758
rect 152016 362914 152044 469882
rect 289084 403028 289136 403034
rect 289084 402970 289136 402976
rect 160744 398880 160796 398886
rect 160744 398822 160796 398828
rect 154580 394800 154632 394806
rect 154580 394742 154632 394748
rect 152096 367736 152148 367742
rect 152096 367678 152148 367684
rect 152004 362908 152056 362914
rect 152004 362850 152056 362856
rect 151912 345772 151964 345778
rect 151912 345714 151964 345720
rect 152108 294642 152136 367678
rect 153108 362908 153160 362914
rect 153108 362850 153160 362856
rect 153120 362234 153148 362850
rect 153108 362228 153160 362234
rect 153108 362170 153160 362176
rect 152096 294636 152148 294642
rect 152096 294578 152148 294584
rect 152462 291952 152518 291961
rect 152462 291887 152518 291896
rect 151820 216640 151872 216646
rect 151820 216582 151872 216588
rect 151084 185768 151136 185774
rect 151084 185710 151136 185716
rect 152476 184482 152504 291887
rect 154592 256698 154620 394742
rect 158720 351280 158772 351286
rect 158720 351222 158772 351228
rect 158732 347070 158760 351222
rect 158720 347064 158772 347070
rect 158720 347006 158772 347012
rect 159364 311296 159416 311302
rect 159364 311238 159416 311244
rect 155224 295588 155276 295594
rect 155224 295530 155276 295536
rect 154580 256692 154632 256698
rect 154580 256634 154632 256640
rect 154592 256086 154620 256634
rect 154580 256080 154632 256086
rect 154580 256022 154632 256028
rect 153108 216640 153160 216646
rect 153108 216582 153160 216588
rect 153120 215966 153148 216582
rect 153108 215960 153160 215966
rect 153108 215902 153160 215908
rect 155236 189990 155264 295530
rect 159376 256018 159404 311238
rect 159364 256012 159416 256018
rect 159364 255954 159416 255960
rect 159364 245744 159416 245750
rect 159364 245686 159416 245692
rect 155224 189984 155276 189990
rect 155224 189926 155276 189932
rect 152464 184476 152516 184482
rect 152464 184418 152516 184424
rect 142804 183048 142856 183054
rect 142804 182990 142856 182996
rect 159376 180266 159404 245686
rect 160756 181762 160784 398822
rect 188344 397588 188396 397594
rect 188344 397530 188396 397536
rect 178684 396772 178736 396778
rect 178684 396714 178736 396720
rect 170404 395344 170456 395350
rect 170404 395286 170456 395292
rect 162124 333328 162176 333334
rect 162124 333270 162176 333276
rect 160836 297016 160888 297022
rect 160836 296958 160888 296964
rect 160848 271182 160876 296958
rect 160836 271176 160888 271182
rect 160836 271118 160888 271124
rect 160744 181756 160796 181762
rect 160744 181698 160796 181704
rect 159364 180260 159416 180266
rect 159364 180202 159416 180208
rect 135904 178016 135956 178022
rect 135904 177958 135956 177964
rect 133144 177948 133196 177954
rect 133144 177890 133196 177896
rect 130750 177712 130806 177721
rect 130750 177647 130806 177656
rect 132406 177712 132462 177721
rect 132406 177647 132462 177656
rect 162136 177313 162164 333270
rect 169024 302456 169076 302462
rect 169024 302398 169076 302404
rect 166264 299668 166316 299674
rect 166264 299610 166316 299616
rect 164884 271924 164936 271930
rect 164884 271866 164936 271872
rect 162122 177304 162178 177313
rect 162122 177239 162178 177248
rect 134432 177064 134484 177070
rect 134432 177006 134484 177012
rect 134444 176769 134472 177006
rect 136088 176792 136140 176798
rect 119526 176760 119582 176769
rect 119526 176695 119582 176704
rect 122102 176760 122158 176769
rect 122102 176695 122158 176704
rect 124494 176760 124550 176769
rect 124494 176695 124550 176704
rect 127898 176760 127954 176769
rect 127898 176695 127954 176704
rect 133142 176760 133198 176769
rect 133142 176695 133144 176704
rect 133196 176695 133198 176704
rect 134430 176760 134486 176769
rect 134430 176695 134486 176704
rect 136086 176760 136088 176769
rect 136140 176760 136142 176769
rect 136086 176695 136142 176704
rect 133144 176666 133196 176672
rect 128176 176316 128228 176322
rect 128176 176258 128228 176264
rect 111064 175976 111116 175982
rect 111064 175918 111116 175924
rect 116952 175976 117004 175982
rect 116952 175918 117004 175924
rect 116964 175545 116992 175918
rect 128188 175545 128216 176258
rect 158904 176248 158956 176254
rect 158904 176190 158956 176196
rect 148232 176180 148284 176186
rect 148232 176122 148284 176128
rect 129464 176044 129516 176050
rect 129464 175986 129516 175992
rect 129476 175545 129504 175986
rect 148244 175545 148272 176122
rect 158916 175545 158944 176190
rect 104622 175536 104678 175545
rect 104622 175471 104678 175480
rect 116950 175536 117006 175545
rect 116950 175471 117006 175480
rect 128174 175536 128230 175545
rect 128174 175471 128230 175480
rect 129462 175536 129518 175545
rect 129462 175471 129518 175480
rect 148230 175536 148286 175545
rect 148230 175471 148286 175480
rect 158902 175536 158958 175545
rect 158902 175471 158958 175480
rect 164896 174049 164924 271866
rect 166276 181490 166304 299610
rect 169036 249082 169064 302398
rect 169024 249076 169076 249082
rect 169024 249018 169076 249024
rect 167828 185020 167880 185026
rect 167828 184962 167880 184968
rect 166356 183592 166408 183598
rect 166356 183534 166408 183540
rect 166264 181484 166316 181490
rect 166264 181426 166316 181432
rect 164976 181076 165028 181082
rect 164976 181018 165028 181024
rect 164882 174040 164938 174049
rect 164882 173975 164938 173984
rect 164988 173874 165016 181018
rect 166264 179580 166316 179586
rect 166264 179522 166316 179528
rect 165528 177064 165580 177070
rect 165528 177006 165580 177012
rect 165252 176928 165304 176934
rect 165252 176870 165304 176876
rect 165264 174554 165292 176870
rect 165540 175234 165568 177006
rect 165528 175228 165580 175234
rect 165528 175170 165580 175176
rect 165252 174548 165304 174554
rect 165252 174490 165304 174496
rect 165618 174040 165674 174049
rect 165618 173975 165674 173984
rect 164976 173868 165028 173874
rect 164976 173810 165028 173816
rect 66074 129296 66130 129305
rect 66074 129231 66130 129240
rect 65522 128072 65578 128081
rect 65522 128007 65578 128016
rect 65536 127022 65564 128007
rect 65524 127016 65576 127022
rect 65524 126958 65576 126964
rect 65982 102368 66038 102377
rect 65982 102303 66038 102312
rect 65996 85542 66024 102303
rect 66088 94761 66116 129231
rect 67362 126304 67418 126313
rect 67362 126239 67418 126248
rect 66166 125216 66222 125225
rect 66166 125151 66222 125160
rect 66074 94752 66130 94761
rect 66074 94687 66130 94696
rect 65984 85536 66036 85542
rect 65984 85478 66036 85484
rect 66180 84153 66208 125151
rect 67376 94897 67404 126239
rect 67546 123584 67602 123593
rect 67546 123519 67602 123528
rect 67454 122632 67510 122641
rect 67454 122567 67510 122576
rect 67362 94888 67418 94897
rect 67362 94823 67418 94832
rect 67468 91089 67496 122567
rect 67454 91080 67510 91089
rect 67454 91015 67510 91024
rect 67560 89729 67588 123519
rect 67638 120864 67694 120873
rect 67638 120799 67694 120808
rect 67546 89720 67602 89729
rect 67652 89690 67680 120799
rect 67730 100736 67786 100745
rect 67730 100671 67786 100680
rect 67546 89655 67602 89664
rect 67640 89684 67692 89690
rect 67640 89626 67692 89632
rect 67744 88330 67772 100671
rect 165632 95674 165660 173975
rect 166276 164218 166304 179522
rect 166368 168298 166396 183534
rect 166540 182300 166592 182306
rect 166540 182242 166592 182248
rect 166448 178084 166500 178090
rect 166448 178026 166500 178032
rect 166460 168366 166488 178026
rect 166552 173806 166580 182242
rect 167736 180940 167788 180946
rect 167736 180882 167788 180888
rect 167000 176316 167052 176322
rect 167000 176258 167052 176264
rect 166540 173800 166592 173806
rect 166540 173742 166592 173748
rect 167012 172514 167040 176258
rect 167000 172508 167052 172514
rect 167000 172450 167052 172456
rect 167642 171592 167698 171601
rect 167642 171527 167698 171536
rect 166448 168360 166500 168366
rect 166448 168302 166500 168308
rect 166356 168292 166408 168298
rect 166356 168234 166408 168240
rect 166264 164212 166316 164218
rect 166264 164154 166316 164160
rect 167656 151094 167684 171527
rect 167748 165510 167776 180882
rect 167840 169726 167868 184962
rect 169024 182232 169076 182238
rect 169024 182174 169076 182180
rect 167920 179512 167972 179518
rect 167920 179454 167972 179460
rect 167828 169720 167880 169726
rect 167828 169662 167880 169668
rect 167932 165578 167960 179454
rect 167920 165572 167972 165578
rect 167920 165514 167972 165520
rect 167736 165504 167788 165510
rect 167736 165446 167788 165452
rect 169036 162858 169064 182174
rect 169208 179444 169260 179450
rect 169208 179386 169260 179392
rect 169116 176860 169168 176866
rect 169116 176802 169168 176808
rect 169024 162852 169076 162858
rect 169024 162794 169076 162800
rect 169128 158710 169156 176802
rect 169220 161430 169248 179386
rect 169300 176112 169352 176118
rect 169300 176054 169352 176060
rect 169208 161424 169260 161430
rect 169208 161366 169260 161372
rect 169312 160070 169340 176054
rect 169300 160064 169352 160070
rect 169300 160006 169352 160012
rect 169116 158704 169168 158710
rect 169116 158646 169168 158652
rect 167644 151088 167696 151094
rect 167644 151030 167696 151036
rect 169024 143608 169076 143614
rect 169024 143550 169076 143556
rect 167644 142860 167696 142866
rect 167644 142802 167696 142808
rect 166264 136672 166316 136678
rect 166264 136614 166316 136620
rect 164884 95668 164936 95674
rect 164884 95610 164936 95616
rect 165620 95668 165672 95674
rect 165620 95610 165672 95616
rect 126518 94208 126574 94217
rect 126518 94143 126574 94152
rect 152094 94208 152150 94217
rect 152094 94143 152096 94152
rect 126532 94110 126560 94143
rect 152148 94143 152150 94152
rect 152096 94114 152148 94120
rect 126520 94104 126572 94110
rect 112350 94072 112406 94081
rect 126520 94046 126572 94052
rect 126702 94072 126758 94081
rect 112350 94007 112406 94016
rect 126702 94007 126704 94016
rect 112364 93974 112392 94007
rect 126756 94007 126758 94016
rect 126704 93978 126756 93984
rect 112352 93968 112404 93974
rect 96158 93936 96214 93945
rect 112352 93910 112404 93916
rect 96158 93871 96160 93880
rect 96212 93871 96214 93880
rect 96160 93842 96212 93848
rect 100942 93528 100998 93537
rect 100942 93463 100998 93472
rect 109222 93528 109278 93537
rect 109222 93463 109278 93472
rect 116766 93528 116822 93537
rect 116766 93463 116822 93472
rect 121734 93528 121790 93537
rect 121734 93463 121790 93472
rect 133142 93528 133198 93537
rect 133142 93463 133144 93472
rect 100956 93158 100984 93463
rect 103334 93256 103390 93265
rect 109236 93226 109264 93463
rect 116780 93294 116808 93463
rect 121748 93362 121776 93463
rect 133196 93463 133198 93472
rect 151726 93528 151782 93537
rect 151726 93463 151782 93472
rect 133144 93434 133196 93440
rect 151740 93430 151768 93463
rect 151728 93424 151780 93430
rect 151728 93366 151780 93372
rect 121736 93356 121788 93362
rect 121736 93298 121788 93304
rect 116768 93288 116820 93294
rect 110142 93256 110198 93265
rect 103334 93191 103390 93200
rect 109224 93220 109276 93226
rect 100944 93152 100996 93158
rect 100944 93094 100996 93100
rect 88984 92472 89036 92478
rect 74814 92440 74870 92449
rect 74814 92375 74870 92384
rect 85854 92440 85910 92449
rect 85854 92375 85910 92384
rect 88062 92440 88118 92449
rect 88062 92375 88118 92384
rect 88982 92440 88984 92449
rect 89036 92440 89038 92449
rect 88982 92375 89038 92384
rect 97538 92440 97594 92449
rect 97538 92375 97594 92384
rect 98826 92440 98882 92449
rect 98826 92375 98882 92384
rect 74828 91186 74856 92375
rect 85486 91216 85542 91225
rect 74816 91180 74868 91186
rect 85486 91151 85542 91160
rect 74816 91122 74868 91128
rect 67732 88324 67784 88330
rect 67732 88266 67784 88272
rect 66166 84144 66222 84153
rect 66166 84079 66222 84088
rect 85500 77246 85528 91151
rect 85868 91118 85896 92375
rect 86774 91216 86830 91225
rect 86774 91151 86830 91160
rect 85856 91112 85908 91118
rect 85856 91054 85908 91060
rect 86788 86834 86816 91151
rect 88076 91050 88104 92375
rect 90730 91760 90786 91769
rect 90730 91695 90786 91704
rect 88984 91180 89036 91186
rect 88984 91122 89036 91128
rect 88064 91044 88116 91050
rect 88064 90986 88116 90992
rect 88996 86970 89024 91122
rect 90744 89554 90772 91695
rect 95054 91352 95110 91361
rect 95054 91287 95110 91296
rect 92386 91216 92442 91225
rect 92386 91151 92442 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 90732 89548 90784 89554
rect 90732 89490 90784 89496
rect 88984 86964 89036 86970
rect 88984 86906 89036 86912
rect 86776 86828 86828 86834
rect 86776 86770 86828 86776
rect 92400 79966 92428 91151
rect 93780 81190 93808 91151
rect 95068 82686 95096 91287
rect 95146 91216 95202 91225
rect 97552 91186 97580 92375
rect 97814 91216 97870 91225
rect 95146 91151 95202 91160
rect 97540 91180 97592 91186
rect 95056 82680 95108 82686
rect 95056 82622 95108 82628
rect 93768 81184 93820 81190
rect 93768 81126 93820 81132
rect 92388 79960 92440 79966
rect 92388 79902 92440 79908
rect 95160 78606 95188 91151
rect 97814 91151 97870 91160
rect 97540 91122 97592 91128
rect 97828 81258 97856 91151
rect 98840 90982 98868 92375
rect 103242 92304 103298 92313
rect 103242 92239 103298 92248
rect 99194 91352 99250 91361
rect 99194 91287 99250 91296
rect 100574 91352 100630 91361
rect 100574 91287 100630 91296
rect 101862 91352 101918 91361
rect 101862 91287 101918 91296
rect 98828 90976 98880 90982
rect 98828 90918 98880 90924
rect 99208 82793 99236 91287
rect 99286 91216 99342 91225
rect 99286 91151 99342 91160
rect 99194 82784 99250 82793
rect 99194 82719 99250 82728
rect 97816 81252 97868 81258
rect 97816 81194 97868 81200
rect 99300 80073 99328 91151
rect 100588 86766 100616 91287
rect 100666 91216 100722 91225
rect 100666 91151 100722 91160
rect 100576 86760 100628 86766
rect 100576 86702 100628 86708
rect 100680 84114 100708 91151
rect 101876 85474 101904 91287
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 101864 85468 101916 85474
rect 101864 85410 101916 85416
rect 100668 84108 100720 84114
rect 100668 84050 100720 84056
rect 99286 80064 99342 80073
rect 99286 79999 99342 80008
rect 95148 78600 95200 78606
rect 95148 78542 95200 78548
rect 102060 78538 102088 91151
rect 103256 90846 103284 92239
rect 103348 92206 103376 93191
rect 116768 93230 116820 93236
rect 110142 93191 110198 93200
rect 109224 93162 109276 93168
rect 103336 92200 103388 92206
rect 103336 92142 103388 92148
rect 106094 91352 106150 91361
rect 106094 91287 106150 91296
rect 107566 91352 107622 91361
rect 107566 91287 107622 91296
rect 104254 91216 104310 91225
rect 104254 91151 104310 91160
rect 104806 91216 104862 91225
rect 104806 91151 104862 91160
rect 103244 90840 103296 90846
rect 103244 90782 103296 90788
rect 104268 88194 104296 91151
rect 104256 88188 104308 88194
rect 104256 88130 104308 88136
rect 104820 82618 104848 91151
rect 106108 84046 106136 91287
rect 106186 91216 106242 91225
rect 106186 91151 106242 91160
rect 107474 91216 107530 91225
rect 107474 91151 107530 91160
rect 106096 84040 106148 84046
rect 106096 83982 106148 83988
rect 104808 82612 104860 82618
rect 104808 82554 104860 82560
rect 106200 81433 106228 91151
rect 107488 84182 107516 91151
rect 107476 84176 107528 84182
rect 107476 84118 107528 84124
rect 107580 82822 107608 91287
rect 107934 91216 107990 91225
rect 107934 91151 107990 91160
rect 108946 91216 109002 91225
rect 108946 91151 109002 91160
rect 107948 86698 107976 91151
rect 107936 86692 107988 86698
rect 107936 86634 107988 86640
rect 107568 82816 107620 82822
rect 107568 82758 107620 82764
rect 106186 81424 106242 81433
rect 106186 81359 106242 81368
rect 108960 79937 108988 91151
rect 110156 89622 110184 93191
rect 114466 92440 114522 92449
rect 114466 92375 114522 92384
rect 114926 92440 114982 92449
rect 114926 92375 114982 92384
rect 115478 92440 115534 92449
rect 115478 92375 115534 92384
rect 118054 92440 118110 92449
rect 118054 92375 118056 92384
rect 114480 92274 114508 92375
rect 114468 92268 114520 92274
rect 114468 92210 114520 92216
rect 110326 91216 110382 91225
rect 110326 91151 110382 91160
rect 110694 91216 110750 91225
rect 110694 91151 110750 91160
rect 111706 91216 111762 91225
rect 111706 91151 111762 91160
rect 113086 91216 113142 91225
rect 113086 91151 113142 91160
rect 113362 91216 113418 91225
rect 113362 91151 113418 91160
rect 114374 91216 114430 91225
rect 114374 91151 114430 91160
rect 110144 89616 110196 89622
rect 110144 89558 110196 89564
rect 108946 79928 109002 79937
rect 108946 79863 109002 79872
rect 102048 78532 102100 78538
rect 102048 78474 102100 78480
rect 85488 77240 85540 77246
rect 85488 77182 85540 77188
rect 110340 77178 110368 91151
rect 110708 88233 110736 91151
rect 110694 88224 110750 88233
rect 110694 88159 110750 88168
rect 111720 81394 111748 91151
rect 111708 81388 111760 81394
rect 111708 81330 111760 81336
rect 113100 79830 113128 91151
rect 113376 85406 113404 91151
rect 113364 85400 113416 85406
rect 113364 85342 113416 85348
rect 114388 85338 114416 91151
rect 114940 90914 114968 92375
rect 115492 92342 115520 92375
rect 118108 92375 118110 92384
rect 132406 92440 132462 92449
rect 132406 92375 132462 92384
rect 151542 92440 151598 92449
rect 151542 92375 151598 92384
rect 118056 92346 118108 92352
rect 115480 92336 115532 92342
rect 115480 92278 115532 92284
rect 122838 92168 122894 92177
rect 132420 92138 132448 92375
rect 122838 92103 122894 92112
rect 132408 92132 132460 92138
rect 119802 91624 119858 91633
rect 119802 91559 119858 91568
rect 115754 91216 115810 91225
rect 117134 91216 117190 91225
rect 115754 91151 115810 91160
rect 116124 91180 116176 91186
rect 114928 90908 114980 90914
rect 114928 90850 114980 90856
rect 114376 85332 114428 85338
rect 114376 85274 114428 85280
rect 113088 79824 113140 79830
rect 113088 79766 113140 79772
rect 115768 78674 115796 91151
rect 117134 91151 117190 91160
rect 118606 91216 118662 91225
rect 118606 91151 118662 91160
rect 116124 91122 116176 91128
rect 116136 88262 116164 91122
rect 116124 88256 116176 88262
rect 116124 88198 116176 88204
rect 117148 86630 117176 91151
rect 117136 86624 117188 86630
rect 117136 86566 117188 86572
rect 118620 83978 118648 91151
rect 119816 89418 119844 91559
rect 120722 91352 120778 91361
rect 120722 91287 120778 91296
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 119804 89412 119856 89418
rect 119804 89354 119856 89360
rect 118608 83972 118660 83978
rect 118608 83914 118660 83920
rect 120000 82754 120028 91151
rect 120736 88126 120764 91287
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 120724 88120 120776 88126
rect 120724 88062 120776 88068
rect 119988 82748 120040 82754
rect 119988 82690 120040 82696
rect 115756 78668 115808 78674
rect 115756 78610 115808 78616
rect 121380 78470 121408 91151
rect 122104 91112 122156 91118
rect 122104 91054 122156 91060
rect 121368 78464 121420 78470
rect 121368 78406 121420 78412
rect 110328 77172 110380 77178
rect 110328 77114 110380 77120
rect 122116 75886 122144 91054
rect 122852 89486 122880 92103
rect 132408 92074 132460 92080
rect 136454 91624 136510 91633
rect 136454 91559 136510 91568
rect 124034 91352 124090 91361
rect 124034 91287 124090 91296
rect 125414 91352 125470 91361
rect 125414 91287 125470 91296
rect 122840 89480 122892 89486
rect 122840 89422 122892 89428
rect 124048 85270 124076 91287
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 124036 85264 124088 85270
rect 124036 85206 124088 85212
rect 124140 83910 124168 91151
rect 124128 83904 124180 83910
rect 124128 83846 124180 83852
rect 125428 81326 125456 91287
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 126518 91216 126574 91225
rect 126518 91151 126574 91160
rect 129462 91216 129518 91225
rect 129462 91151 129518 91160
rect 130750 91216 130806 91225
rect 130750 91151 130806 91160
rect 135166 91216 135222 91225
rect 135166 91151 135222 91160
rect 125416 81320 125468 81326
rect 125416 81262 125468 81268
rect 125520 79898 125548 91151
rect 126532 86902 126560 91151
rect 129476 88058 129504 91151
rect 129464 88052 129516 88058
rect 129464 87994 129516 88000
rect 126520 86896 126572 86902
rect 126520 86838 126572 86844
rect 130764 85513 130792 91151
rect 130750 85504 130806 85513
rect 130750 85439 130806 85448
rect 135180 82550 135208 91151
rect 136468 89350 136496 91559
rect 151556 90778 151584 92375
rect 151634 92168 151690 92177
rect 151634 92103 151690 92112
rect 151544 90772 151596 90778
rect 151544 90714 151596 90720
rect 151648 90710 151676 92103
rect 151636 90704 151688 90710
rect 151636 90646 151688 90652
rect 136456 89344 136508 89350
rect 136456 89286 136508 89292
rect 135168 82544 135220 82550
rect 135168 82486 135220 82492
rect 125508 79892 125560 79898
rect 125508 79834 125560 79840
rect 122104 75880 122156 75886
rect 122104 75822 122156 75828
rect 93860 75268 93912 75274
rect 93860 75210 93912 75216
rect 69020 75200 69072 75206
rect 69020 75142 69072 75148
rect 67638 64152 67694 64161
rect 67638 64087 67694 64096
rect 64880 60104 64932 60110
rect 64880 60046 64932 60052
rect 64788 29640 64840 29646
rect 64788 29582 64840 29588
rect 64604 20664 64656 20670
rect 64604 20606 64656 20612
rect 64892 16574 64920 60046
rect 60752 16546 60872 16574
rect 62132 16546 63264 16574
rect 64892 16546 65104 16574
rect 60844 480 60872 16546
rect 62028 9036 62080 9042
rect 62028 8978 62080 8984
rect 62040 480 62068 8978
rect 63236 480 63264 16546
rect 64328 2100 64380 2106
rect 64328 2042 64380 2048
rect 64340 480 64368 2042
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65076 354 65104 16546
rect 66720 14544 66772 14550
rect 66720 14486 66772 14492
rect 66732 480 66760 14486
rect 65494 354 65606 480
rect 65076 326 65606 354
rect 65494 -960 65606 326
rect 66690 -960 66802 480
rect 67652 354 67680 64087
rect 69032 3534 69060 75142
rect 89720 71052 89772 71058
rect 89720 70994 89772 71000
rect 86960 69692 87012 69698
rect 86960 69634 87012 69640
rect 75920 68400 75972 68406
rect 75920 68342 75972 68348
rect 73160 65544 73212 65550
rect 73160 65486 73212 65492
rect 70400 62824 70452 62830
rect 70400 62766 70452 62772
rect 69112 58676 69164 58682
rect 69112 58618 69164 58624
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 69124 480 69152 58618
rect 70412 16574 70440 62766
rect 71780 57316 71832 57322
rect 71780 57258 71832 57264
rect 71792 16574 71820 57258
rect 73172 16574 73200 65486
rect 74540 61464 74592 61470
rect 74540 61406 74592 61412
rect 74552 16574 74580 61406
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69940 3528 69992 3534
rect 69940 3470 69992 3476
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69952 354 69980 3470
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69952 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 68342
rect 85580 58812 85632 58818
rect 85580 58754 85632 58760
rect 82820 54664 82872 54670
rect 82820 54606 82872 54612
rect 80060 32496 80112 32502
rect 80060 32438 80112 32444
rect 80072 16574 80100 32438
rect 81440 28280 81492 28286
rect 81440 28222 81492 28228
rect 81452 16574 81480 28222
rect 82832 16574 82860 54606
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 77392 11824 77444 11830
rect 77392 11766 77444 11772
rect 77404 480 77432 11766
rect 79692 6248 79744 6254
rect 79692 6190 79744 6196
rect 78588 3596 78640 3602
rect 78588 3538 78640 3544
rect 78600 480 78628 3538
rect 79704 480 79732 6190
rect 80900 480 80928 16546
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 84200 14612 84252 14618
rect 84200 14554 84252 14560
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 14554
rect 85592 6914 85620 58754
rect 85672 50448 85724 50454
rect 85672 50390 85724 50396
rect 85684 16574 85712 50390
rect 86972 16574 87000 69634
rect 88984 68332 89036 68338
rect 88984 68274 89036 68280
rect 85684 16546 86448 16574
rect 86972 16546 87552 16574
rect 85592 6886 85712 6914
rect 85684 480 85712 6886
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 16546
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 16546
rect 88996 3602 89024 68274
rect 89732 16574 89760 70994
rect 92480 43512 92532 43518
rect 92480 43454 92532 43460
rect 91100 38004 91152 38010
rect 91100 37946 91152 37952
rect 91112 16574 91140 37946
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 88984 3596 89036 3602
rect 88984 3538 89036 3544
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 89180 480 89208 3470
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 43454
rect 93872 3602 93900 75210
rect 104900 73908 104952 73914
rect 104900 73850 104952 73856
rect 102140 73840 102192 73846
rect 102140 73782 102192 73788
rect 93952 56024 94004 56030
rect 93952 55966 94004 55972
rect 93860 3596 93912 3602
rect 93860 3538 93912 3544
rect 93964 480 93992 55966
rect 99380 49088 99432 49094
rect 99380 49030 99432 49036
rect 95240 45008 95292 45014
rect 95240 44950 95292 44956
rect 95252 16574 95280 44950
rect 99392 16574 99420 49030
rect 100760 18760 100812 18766
rect 100760 18702 100812 18708
rect 95252 16546 95832 16574
rect 99392 16546 99880 16574
rect 94780 3596 94832 3602
rect 94780 3538 94832 3544
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3538
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97448 13184 97500 13190
rect 97448 13126 97500 13132
rect 97460 480 97488 13126
rect 98184 11756 98236 11762
rect 98184 11698 98236 11704
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 11698
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 18702
rect 102152 16574 102180 73782
rect 103520 17332 103572 17338
rect 103520 17274 103572 17280
rect 103532 16574 103560 17274
rect 104912 16574 104940 73850
rect 115940 71120 115992 71126
rect 115940 71062 115992 71068
rect 106280 65612 106332 65618
rect 106280 65554 106332 65560
rect 106292 16574 106320 65554
rect 111800 60172 111852 60178
rect 111800 60114 111852 60120
rect 110420 54732 110472 54738
rect 110420 54674 110472 54680
rect 110432 16574 110460 54674
rect 111812 16574 111840 60114
rect 114560 51740 114612 51746
rect 114560 51682 114612 51688
rect 113180 50516 113232 50522
rect 113180 50458 113232 50464
rect 113192 16574 113220 50458
rect 114572 16574 114600 51682
rect 115952 16574 115980 71062
rect 122840 68468 122892 68474
rect 122840 68410 122892 68416
rect 117320 53236 117372 53242
rect 117320 53178 117372 53184
rect 102152 16546 102272 16574
rect 103532 16546 104112 16574
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 110432 16546 110552 16574
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 102244 480 102272 16546
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103348 480 103376 3538
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 16546
rect 105740 480 105768 16546
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108120 15972 108172 15978
rect 108120 15914 108172 15920
rect 108132 480 108160 15914
rect 109316 7676 109368 7682
rect 109316 7618 109368 7624
rect 109328 480 109356 7618
rect 110524 480 110552 16546
rect 111616 2168 111668 2174
rect 111616 2110 111668 2116
rect 111628 480 111656 2110
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 53178
rect 120080 51808 120132 51814
rect 120080 51750 120132 51756
rect 118700 47660 118752 47666
rect 118700 47602 118752 47608
rect 118712 6914 118740 47602
rect 118792 24268 118844 24274
rect 118792 24210 118844 24216
rect 118804 16574 118832 24210
rect 120092 16574 120120 51750
rect 121460 44940 121512 44946
rect 121460 44882 121512 44888
rect 121472 16574 121500 44882
rect 122852 16574 122880 68410
rect 132500 53168 132552 53174
rect 132500 53110 132552 53116
rect 132512 16574 132540 53110
rect 135260 35284 135312 35290
rect 135260 35226 135312 35232
rect 118804 16546 119936 16574
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 132512 16546 133000 16574
rect 118712 6886 118832 6914
rect 118804 480 118832 6886
rect 119908 480 119936 16546
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124680 10328 124732 10334
rect 124680 10270 124732 10276
rect 124692 480 124720 10270
rect 125876 3664 125928 3670
rect 125876 3606 125928 3612
rect 125888 480 125916 3606
rect 129372 2236 129424 2242
rect 129372 2178 129424 2184
rect 129384 480 129412 2178
rect 132972 480 133000 16546
rect 135272 3398 135300 35226
rect 164424 14476 164476 14482
rect 164424 14418 164476 14424
rect 135260 3392 135312 3398
rect 135260 3334 135312 3340
rect 136456 3392 136508 3398
rect 136456 3334 136508 3340
rect 136468 480 136496 3334
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 14418
rect 164896 3670 164924 95610
rect 166276 93294 166304 136614
rect 166356 111852 166408 111858
rect 166356 111794 166408 111800
rect 166264 93288 166316 93294
rect 166264 93230 166316 93236
rect 166368 86766 166396 111794
rect 167656 108769 167684 142802
rect 167828 122868 167880 122874
rect 167828 122810 167880 122816
rect 167736 114572 167788 114578
rect 167736 114514 167788 114520
rect 167642 108760 167698 108769
rect 167642 108695 167698 108704
rect 167644 106344 167696 106350
rect 167644 106286 167696 106292
rect 166448 98048 166500 98054
rect 166448 97990 166500 97996
rect 166460 86834 166488 97990
rect 166908 95940 166960 95946
rect 166908 95882 166960 95888
rect 166920 92478 166948 95882
rect 166908 92472 166960 92478
rect 166908 92414 166960 92420
rect 166448 86828 166500 86834
rect 166448 86770 166500 86776
rect 166356 86760 166408 86766
rect 166356 86702 166408 86708
rect 167656 81190 167684 106286
rect 167748 84046 167776 114514
rect 167840 93362 167868 122810
rect 167920 113212 167972 113218
rect 167920 113154 167972 113160
rect 167828 93356 167880 93362
rect 167828 93298 167880 93304
rect 167932 90846 167960 113154
rect 168012 111784 168064 111790
rect 168010 111752 168012 111761
rect 168064 111752 168066 111761
rect 168010 111687 168066 111696
rect 168104 110424 168156 110430
rect 168104 110366 168156 110372
rect 168116 110129 168144 110366
rect 168102 110120 168158 110129
rect 168102 110055 168158 110064
rect 167920 90840 167972 90846
rect 167920 90782 167972 90788
rect 169036 88058 169064 143550
rect 169116 125656 169168 125662
rect 169116 125598 169168 125604
rect 169128 94110 169156 125598
rect 170416 122126 170444 395286
rect 177304 337476 177356 337482
rect 177304 337418 177356 337424
rect 171784 228608 171836 228614
rect 171784 228550 171836 228556
rect 170496 190596 170548 190602
rect 170496 190538 170548 190544
rect 170508 157350 170536 190538
rect 171796 181626 171824 228550
rect 173164 189100 173216 189106
rect 173164 189042 173216 189048
rect 171784 181620 171836 181626
rect 171784 181562 171836 181568
rect 171876 181008 171928 181014
rect 171876 180950 171928 180956
rect 170588 180872 170640 180878
rect 170588 180814 170640 180820
rect 170496 157344 170548 157350
rect 170496 157286 170548 157292
rect 170600 155922 170628 180814
rect 170680 176996 170732 177002
rect 170680 176938 170732 176944
rect 170692 169658 170720 176938
rect 170680 169652 170732 169658
rect 170680 169594 170732 169600
rect 171888 167006 171916 180950
rect 171876 167000 171928 167006
rect 171876 166942 171928 166948
rect 173176 157282 173204 189042
rect 173164 157276 173216 157282
rect 173164 157218 173216 157224
rect 170588 155916 170640 155922
rect 170588 155858 170640 155864
rect 173164 151972 173216 151978
rect 173164 151914 173216 151920
rect 171784 146328 171836 146334
rect 171784 146270 171836 146276
rect 170496 143676 170548 143682
rect 170496 143618 170548 143624
rect 170404 122120 170456 122126
rect 170404 122062 170456 122068
rect 170404 117360 170456 117366
rect 170404 117302 170456 117308
rect 169208 116000 169260 116006
rect 169208 115942 169260 115948
rect 169116 94104 169168 94110
rect 169116 94046 169168 94052
rect 169024 88052 169076 88058
rect 169024 87994 169076 88000
rect 169220 86698 169248 115942
rect 169300 110492 169352 110498
rect 169300 110434 169352 110440
rect 169208 86692 169260 86698
rect 169208 86634 169260 86640
rect 169312 84114 169340 110434
rect 170416 89622 170444 117302
rect 170508 90953 170536 143618
rect 170588 124228 170640 124234
rect 170588 124170 170640 124176
rect 170494 90944 170550 90953
rect 170494 90879 170550 90888
rect 170404 89616 170456 89622
rect 170404 89558 170456 89564
rect 170600 85270 170628 124170
rect 170680 107704 170732 107710
rect 170680 107646 170732 107652
rect 170588 85264 170640 85270
rect 170588 85206 170640 85212
rect 170402 84824 170458 84833
rect 170402 84759 170458 84768
rect 169300 84108 169352 84114
rect 169300 84050 169352 84056
rect 167736 84040 167788 84046
rect 167736 83982 167788 83988
rect 167644 81184 167696 81190
rect 167644 81126 167696 81132
rect 164884 3664 164936 3670
rect 164884 3606 164936 3612
rect 170416 3602 170444 84759
rect 170692 82686 170720 107646
rect 171796 93498 171824 146270
rect 171968 135312 172020 135318
rect 171968 135254 172020 135260
rect 171876 129804 171928 129810
rect 171876 129746 171928 129752
rect 171784 93492 171836 93498
rect 171784 93434 171836 93440
rect 170680 82680 170732 82686
rect 170680 82622 170732 82628
rect 171888 78538 171916 129746
rect 171980 85338 172008 135254
rect 172060 109064 172112 109070
rect 172060 109006 172112 109012
rect 172072 93906 172100 109006
rect 172060 93900 172112 93906
rect 172060 93842 172112 93848
rect 173176 90710 173204 151914
rect 176016 150476 176068 150482
rect 176016 150418 176068 150424
rect 174544 140820 174596 140826
rect 174544 140762 174596 140768
rect 173256 131164 173308 131170
rect 173256 131106 173308 131112
rect 173164 90704 173216 90710
rect 173164 90646 173216 90652
rect 171968 85332 172020 85338
rect 171968 85274 172020 85280
rect 173268 82618 173296 131106
rect 173440 104916 173492 104922
rect 173440 104858 173492 104864
rect 173348 102808 173400 102814
rect 173348 102750 173400 102756
rect 173360 92206 173388 102750
rect 173452 94761 173480 104858
rect 173438 94752 173494 94761
rect 173438 94687 173494 94696
rect 173348 92200 173400 92206
rect 173348 92142 173400 92148
rect 174556 83910 174584 140762
rect 174636 138032 174688 138038
rect 174636 137974 174688 137980
rect 174648 89418 174676 137974
rect 175924 133952 175976 133958
rect 175924 133894 175976 133900
rect 174820 116068 174872 116074
rect 174820 116010 174872 116016
rect 174728 107772 174780 107778
rect 174728 107714 174780 107720
rect 174636 89412 174688 89418
rect 174636 89354 174688 89360
rect 174544 83904 174596 83910
rect 174544 83846 174596 83852
rect 173256 82612 173308 82618
rect 173256 82554 173308 82560
rect 174740 78606 174768 107714
rect 174832 93226 174860 116010
rect 174820 93220 174872 93226
rect 174820 93162 174872 93168
rect 174728 78600 174780 78606
rect 174728 78542 174780 78548
rect 171876 78532 171928 78538
rect 171876 78474 171928 78480
rect 175936 77178 175964 133894
rect 176028 111790 176056 150418
rect 176108 120148 176160 120154
rect 176108 120090 176160 120096
rect 176016 111784 176068 111790
rect 176016 111726 176068 111732
rect 176016 106412 176068 106418
rect 176016 106354 176068 106360
rect 176028 79966 176056 106354
rect 176120 86630 176148 120090
rect 176108 86624 176160 86630
rect 176108 86566 176160 86572
rect 176016 79960 176068 79966
rect 176016 79902 176068 79908
rect 175924 77172 175976 77178
rect 175924 77114 175976 77120
rect 177316 76566 177344 337418
rect 177396 140072 177448 140078
rect 177396 140014 177448 140020
rect 177408 92138 177436 140014
rect 177488 118720 177540 118726
rect 177488 118662 177540 118668
rect 177396 92132 177448 92138
rect 177396 92074 177448 92080
rect 177500 85406 177528 118662
rect 177580 100768 177632 100774
rect 177580 100710 177632 100716
rect 177488 85400 177540 85406
rect 177488 85342 177540 85348
rect 177592 77246 177620 100710
rect 177580 77240 177632 77246
rect 177580 77182 177632 77188
rect 177304 76560 177356 76566
rect 177304 76502 177356 76508
rect 178696 35290 178724 396714
rect 186964 392624 187016 392630
rect 186964 392566 187016 392572
rect 184204 388136 184256 388142
rect 184204 388078 184256 388084
rect 180064 348424 180116 348430
rect 180064 348366 180116 348372
rect 178774 294264 178830 294273
rect 178774 294199 178830 294208
rect 178788 95198 178816 294199
rect 178868 153264 178920 153270
rect 178868 153206 178920 153212
rect 178776 95192 178828 95198
rect 178776 95134 178828 95140
rect 178880 90778 178908 153206
rect 178960 122936 179012 122942
rect 178960 122878 179012 122884
rect 178868 90772 178920 90778
rect 178868 90714 178920 90720
rect 178972 88126 179000 122878
rect 178960 88120 179012 88126
rect 178960 88062 179012 88068
rect 178776 83496 178828 83502
rect 178776 83438 178828 83444
rect 178684 35284 178736 35290
rect 178684 35226 178736 35232
rect 170404 3596 170456 3602
rect 170404 3538 170456 3544
rect 178788 3534 178816 83438
rect 180076 33114 180104 348366
rect 181444 238264 181496 238270
rect 181444 238206 181496 238212
rect 180156 127016 180208 127022
rect 180156 126958 180208 126964
rect 180168 81258 180196 126958
rect 180248 121508 180300 121514
rect 180248 121450 180300 121456
rect 180260 83978 180288 121450
rect 181456 95130 181484 238206
rect 182824 234116 182876 234122
rect 182824 234058 182876 234064
rect 181536 142180 181588 142186
rect 181536 142122 181588 142128
rect 181444 95124 181496 95130
rect 181444 95066 181496 95072
rect 181548 94042 181576 142122
rect 181536 94036 181588 94042
rect 181536 93978 181588 93984
rect 182836 89622 182864 234058
rect 182916 147688 182968 147694
rect 182916 147630 182968 147636
rect 182824 89616 182876 89622
rect 182824 89558 182876 89564
rect 182928 89350 182956 147630
rect 182916 89344 182968 89350
rect 182916 89286 182968 89292
rect 180248 83972 180300 83978
rect 180248 83914 180300 83920
rect 180156 81252 180208 81258
rect 180156 81194 180208 81200
rect 184216 79354 184244 388078
rect 184294 177304 184350 177313
rect 184294 177239 184350 177248
rect 184204 79348 184256 79354
rect 184204 79290 184256 79296
rect 184308 34474 184336 177239
rect 184572 151088 184624 151094
rect 184572 151030 184624 151036
rect 184584 150414 184612 151030
rect 184572 150408 184624 150414
rect 184572 150350 184624 150356
rect 185584 146396 185636 146402
rect 185584 146338 185636 146344
rect 184388 139460 184440 139466
rect 184388 139402 184440 139408
rect 184400 78470 184428 139402
rect 184480 110560 184532 110566
rect 184480 110502 184532 110508
rect 184492 90982 184520 110502
rect 184480 90976 184532 90982
rect 184480 90918 184532 90924
rect 185596 82550 185624 146338
rect 185676 118788 185728 118794
rect 185676 118730 185728 118736
rect 185688 93974 185716 118730
rect 185676 93968 185728 93974
rect 185676 93910 185728 93916
rect 185584 82544 185636 82550
rect 185584 82486 185636 82492
rect 184388 78464 184440 78470
rect 184388 78406 184440 78412
rect 184296 34468 184348 34474
rect 184296 34410 184348 34416
rect 180064 33108 180116 33114
rect 180064 33050 180116 33056
rect 186976 22846 187004 392566
rect 187056 301096 187108 301102
rect 187056 301038 187108 301044
rect 187068 254590 187096 301038
rect 187056 254584 187108 254590
rect 187056 254526 187108 254532
rect 187056 184476 187108 184482
rect 187056 184418 187108 184424
rect 187068 92478 187096 184418
rect 187148 132524 187200 132530
rect 187148 132466 187200 132472
rect 187056 92472 187108 92478
rect 187056 92414 187108 92420
rect 187160 84182 187188 132466
rect 187148 84176 187200 84182
rect 187148 84118 187200 84124
rect 186964 22840 187016 22846
rect 186964 22782 187016 22788
rect 188356 7750 188384 397530
rect 202144 397520 202196 397526
rect 202144 397462 202196 397468
rect 195244 394732 195296 394738
rect 195244 394674 195296 394680
rect 191104 362228 191156 362234
rect 191104 362170 191156 362176
rect 188434 294128 188490 294137
rect 188434 294063 188490 294072
rect 188448 93537 188476 294063
rect 189724 151904 189776 151910
rect 189724 151846 189776 151852
rect 188528 128376 188580 128382
rect 188528 128318 188580 128324
rect 188434 93528 188490 93537
rect 188434 93463 188490 93472
rect 188540 93158 188568 128318
rect 188620 104984 188672 104990
rect 188620 104926 188672 104932
rect 188528 93152 188580 93158
rect 188528 93094 188580 93100
rect 188632 89554 188660 104926
rect 189736 94178 189764 151846
rect 189724 94172 189776 94178
rect 189724 94114 189776 94120
rect 188620 89548 188672 89554
rect 188620 89490 188672 89496
rect 191116 13258 191144 362170
rect 192484 309868 192536 309874
rect 192484 309810 192536 309816
rect 191196 298376 191248 298382
rect 191196 298318 191248 298324
rect 191208 96626 191236 298318
rect 191288 153332 191340 153338
rect 191288 153274 191340 153280
rect 191196 96620 191248 96626
rect 191196 96562 191248 96568
rect 191300 93430 191328 153274
rect 191288 93424 191340 93430
rect 191288 93366 191340 93372
rect 192496 49706 192524 309810
rect 193864 302320 193916 302326
rect 193864 302262 193916 302268
rect 193876 95062 193904 302262
rect 193956 118856 194008 118862
rect 193956 118798 194008 118804
rect 193864 95056 193916 95062
rect 193864 94998 193916 95004
rect 193968 90914 193996 118798
rect 193956 90908 194008 90914
rect 193956 90850 194008 90856
rect 192484 49700 192536 49706
rect 192484 49642 192536 49648
rect 195256 36650 195284 394674
rect 196624 393984 196676 393990
rect 196624 393926 196676 393932
rect 195336 298784 195388 298790
rect 195336 298726 195388 298732
rect 195348 203590 195376 298726
rect 195336 203584 195388 203590
rect 195336 203526 195388 203532
rect 195336 190528 195388 190534
rect 195336 190470 195388 190476
rect 195348 160002 195376 190470
rect 195336 159996 195388 160002
rect 195336 159938 195388 159944
rect 195336 138100 195388 138106
rect 195336 138042 195388 138048
rect 195348 92410 195376 138042
rect 195428 113280 195480 113286
rect 195428 113222 195480 113228
rect 195336 92404 195388 92410
rect 195336 92346 195388 92352
rect 195440 88194 195468 113222
rect 195428 88188 195480 88194
rect 195428 88130 195480 88136
rect 196636 38078 196664 393926
rect 198096 389224 198148 389230
rect 198096 389166 198148 389172
rect 198004 325032 198056 325038
rect 198004 324974 198056 324980
rect 196716 303952 196768 303958
rect 196716 303894 196768 303900
rect 196728 192642 196756 303894
rect 196716 192636 196768 192642
rect 196716 192578 196768 192584
rect 196808 184408 196860 184414
rect 196808 184350 196860 184356
rect 196716 122120 196768 122126
rect 196716 122062 196768 122068
rect 196624 38072 196676 38078
rect 196624 38014 196676 38020
rect 195244 36644 195296 36650
rect 195244 36586 195296 36592
rect 196728 25702 196756 122062
rect 196820 92410 196848 184350
rect 196900 117428 196952 117434
rect 196900 117370 196952 117376
rect 196808 92404 196860 92410
rect 196808 92346 196860 92352
rect 196912 81394 196940 117370
rect 196900 81388 196952 81394
rect 196900 81330 196952 81336
rect 196716 25696 196768 25702
rect 196716 25638 196768 25644
rect 191104 13252 191156 13258
rect 191104 13194 191156 13200
rect 188344 7744 188396 7750
rect 188344 7686 188396 7692
rect 198016 4146 198044 324974
rect 198108 86193 198136 389166
rect 200764 387932 200816 387938
rect 200764 387874 200816 387880
rect 199384 192704 199436 192710
rect 199384 192646 199436 192652
rect 198188 121576 198240 121582
rect 198188 121518 198240 121524
rect 198094 86184 198150 86193
rect 198094 86119 198150 86128
rect 198200 82754 198228 121518
rect 199396 94994 199424 192646
rect 199476 124296 199528 124302
rect 199476 124238 199528 124244
rect 199384 94988 199436 94994
rect 199384 94930 199436 94936
rect 199488 89486 199516 124238
rect 199568 98116 199620 98122
rect 199568 98058 199620 98064
rect 199476 89480 199528 89486
rect 199476 89422 199528 89428
rect 198188 82748 198240 82754
rect 198188 82690 198240 82696
rect 199580 75886 199608 98058
rect 200776 91798 200804 387874
rect 200764 91792 200816 91798
rect 200764 91734 200816 91740
rect 202156 79422 202184 397462
rect 228364 391264 228416 391270
rect 228364 391206 228416 391212
rect 204904 388476 204956 388482
rect 204904 388418 204956 388424
rect 202234 292768 202290 292777
rect 202234 292703 202290 292712
rect 202248 181694 202276 292703
rect 203524 181756 203576 181762
rect 203524 181698 203576 181704
rect 202236 181688 202288 181694
rect 202236 181630 202288 181636
rect 202236 130416 202288 130422
rect 202236 130358 202288 130364
rect 202248 92274 202276 130358
rect 202328 125724 202380 125730
rect 202328 125666 202380 125672
rect 202236 92268 202288 92274
rect 202236 92210 202288 92216
rect 202234 90400 202290 90409
rect 202234 90335 202290 90344
rect 202144 79416 202196 79422
rect 202144 79358 202196 79364
rect 199568 75880 199620 75886
rect 199568 75822 199620 75828
rect 198004 4140 198056 4146
rect 198004 4082 198056 4088
rect 178776 3528 178828 3534
rect 178776 3470 178828 3476
rect 202248 3466 202276 90335
rect 202340 79898 202368 125666
rect 202328 79892 202380 79898
rect 202328 79834 202380 79840
rect 203536 67590 203564 181698
rect 203616 105052 203668 105058
rect 203616 104994 203668 105000
rect 203628 93673 203656 104994
rect 203614 93664 203670 93673
rect 203614 93599 203670 93608
rect 204916 80034 204944 388418
rect 206284 358828 206336 358834
rect 206284 358770 206336 358776
rect 204996 316736 205048 316742
rect 204996 316678 205048 316684
rect 204904 80028 204956 80034
rect 204904 79970 204956 79976
rect 203524 67584 203576 67590
rect 203524 67526 203576 67532
rect 205008 51882 205036 316678
rect 206296 82142 206324 358770
rect 213184 351212 213236 351218
rect 213184 351154 213236 351160
rect 209044 345704 209096 345710
rect 209044 345646 209096 345652
rect 207664 320952 207716 320958
rect 207664 320894 207716 320900
rect 206376 243024 206428 243030
rect 206376 242966 206428 242972
rect 206388 184414 206416 242966
rect 206376 184408 206428 184414
rect 206376 184350 206428 184356
rect 206376 182844 206428 182850
rect 206376 182786 206428 182792
rect 206388 94926 206416 182786
rect 206468 135380 206520 135386
rect 206468 135322 206520 135328
rect 206376 94920 206428 94926
rect 206376 94862 206428 94868
rect 206284 82136 206336 82142
rect 206284 82078 206336 82084
rect 206480 79830 206508 135322
rect 206560 103556 206612 103562
rect 206560 103498 206612 103504
rect 206572 94897 206600 103498
rect 206558 94888 206614 94897
rect 206558 94823 206614 94832
rect 207676 83570 207704 320894
rect 207664 83564 207716 83570
rect 207664 83506 207716 83512
rect 209056 80714 209084 345646
rect 211804 337408 211856 337414
rect 211804 337350 211856 337356
rect 209228 186380 209280 186386
rect 209228 186322 209280 186328
rect 209136 176180 209188 176186
rect 209136 176122 209188 176128
rect 209148 150346 209176 176122
rect 209240 171086 209268 186322
rect 209228 171080 209280 171086
rect 209228 171022 209280 171028
rect 209136 150340 209188 150346
rect 209136 150282 209188 150288
rect 209136 140888 209188 140894
rect 209136 140830 209188 140836
rect 209148 81326 209176 140830
rect 210424 136740 210476 136746
rect 210424 136682 210476 136688
rect 209228 102196 209280 102202
rect 209228 102138 209280 102144
rect 209240 89729 209268 102138
rect 210436 92342 210464 136682
rect 210516 120216 210568 120222
rect 210516 120158 210568 120164
rect 210424 92336 210476 92342
rect 210424 92278 210476 92284
rect 209226 89720 209282 89729
rect 209226 89655 209282 89664
rect 209136 81320 209188 81326
rect 209136 81262 209188 81268
rect 209044 80708 209096 80714
rect 209044 80650 209096 80656
rect 206468 79824 206520 79830
rect 206468 79766 206520 79772
rect 210528 78674 210556 120158
rect 211816 86290 211844 337350
rect 211896 176248 211948 176254
rect 211896 176190 211948 176196
rect 211908 149054 211936 176190
rect 211896 149048 211948 149054
rect 211896 148990 211948 148996
rect 211896 114640 211948 114646
rect 211896 114582 211948 114588
rect 211804 86284 211856 86290
rect 211804 86226 211856 86232
rect 211908 82822 211936 114582
rect 211988 99408 212040 99414
rect 211988 99350 212040 99356
rect 212000 91050 212028 99350
rect 211988 91044 212040 91050
rect 211988 90986 212040 90992
rect 213196 87650 213224 351154
rect 215944 347132 215996 347138
rect 215944 347074 215996 347080
rect 213276 306536 213328 306542
rect 213276 306478 213328 306484
rect 213288 188562 213316 306478
rect 214656 301028 214708 301034
rect 214656 300970 214708 300976
rect 214564 289876 214616 289882
rect 214564 289818 214616 289824
rect 213276 188556 213328 188562
rect 213276 188498 213328 188504
rect 214576 177342 214604 289818
rect 214668 192710 214696 300970
rect 214656 192704 214708 192710
rect 214656 192646 214708 192652
rect 214656 187740 214708 187746
rect 214656 187682 214708 187688
rect 214564 177336 214616 177342
rect 214564 177278 214616 177284
rect 213920 176792 213972 176798
rect 213920 176734 213972 176740
rect 213932 176225 213960 176734
rect 214012 176656 214064 176662
rect 214012 176598 214064 176604
rect 213918 176216 213974 176225
rect 213918 176151 213974 176160
rect 213368 175976 213420 175982
rect 213368 175918 213420 175924
rect 213274 175400 213330 175409
rect 213274 175335 213330 175344
rect 213288 155961 213316 175335
rect 213380 166161 213408 175918
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175137 213960 175170
rect 213918 175128 213974 175137
rect 213918 175063 213974 175072
rect 214024 174729 214052 176598
rect 214104 176044 214156 176050
rect 214104 175986 214156 175992
rect 214010 174720 214066 174729
rect 214010 174655 214066 174664
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173777 213960 173810
rect 214012 173800 214064 173806
rect 213918 173768 213974 173777
rect 214012 173742 214064 173748
rect 213918 173703 213974 173712
rect 214024 173369 214052 173742
rect 214010 173360 214066 173369
rect 214010 173295 214066 173304
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172009 213960 172450
rect 214116 172417 214144 175986
rect 214564 174548 214616 174554
rect 214564 174490 214616 174496
rect 214102 172408 214158 172417
rect 214102 172343 214158 172352
rect 213918 172000 213974 172009
rect 213918 171935 213974 171944
rect 213920 171080 213972 171086
rect 213918 171048 213920 171057
rect 213972 171048 213974 171057
rect 213918 170983 213974 170992
rect 214012 169720 214064 169726
rect 213918 169688 213974 169697
rect 214012 169662 214064 169668
rect 213918 169623 213920 169632
rect 213972 169623 213974 169632
rect 213920 169594 213972 169600
rect 214024 169425 214052 169662
rect 214010 169416 214066 169425
rect 214010 169351 214066 169360
rect 213920 168360 213972 168366
rect 213920 168302 213972 168308
rect 213932 168065 213960 168302
rect 214012 168292 214064 168298
rect 214012 168234 214064 168240
rect 213918 168056 213974 168065
rect 213918 167991 213974 168000
rect 214024 167929 214052 168234
rect 214010 167920 214066 167929
rect 214010 167855 214066 167864
rect 213920 167000 213972 167006
rect 213920 166942 213972 166948
rect 213932 166705 213960 166942
rect 213918 166696 213974 166705
rect 213918 166631 213974 166640
rect 213366 166152 213422 166161
rect 213366 166087 213422 166096
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165345 213960 165514
rect 214012 165504 214064 165510
rect 214012 165446 214064 165452
rect 213918 165336 213974 165345
rect 213918 165271 213974 165280
rect 214024 164801 214052 165446
rect 214010 164792 214066 164801
rect 214010 164727 214066 164736
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163985 213960 164154
rect 213918 163976 213974 163985
rect 213918 163911 213974 163920
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162625 213960 162794
rect 213918 162616 213974 162625
rect 213918 162551 213974 162560
rect 213920 161424 213972 161430
rect 213918 161392 213920 161401
rect 213972 161392 213974 161401
rect 213918 161327 213974 161336
rect 214576 160857 214604 174490
rect 214668 166977 214696 187682
rect 214748 184952 214800 184958
rect 214748 184894 214800 184900
rect 214760 170785 214788 184894
rect 214746 170776 214802 170785
rect 214746 170711 214802 170720
rect 214654 166968 214710 166977
rect 214654 166903 214710 166912
rect 214562 160848 214618 160857
rect 214562 160783 214618 160792
rect 214102 160712 214158 160721
rect 214102 160647 214158 160656
rect 214012 160064 214064 160070
rect 214012 160006 214064 160012
rect 213920 159996 213972 160002
rect 213920 159938 213972 159944
rect 213932 159905 213960 159938
rect 213918 159896 213974 159905
rect 213918 159831 213974 159840
rect 214024 159497 214052 160006
rect 214010 159488 214066 159497
rect 214010 159423 214066 159432
rect 213920 158704 213972 158710
rect 213918 158672 213920 158681
rect 213972 158672 213974 158681
rect 213918 158607 213974 158616
rect 214116 158137 214144 160647
rect 214102 158128 214158 158137
rect 214102 158063 214158 158072
rect 214012 157344 214064 157350
rect 213918 157312 213974 157321
rect 214012 157286 214064 157292
rect 213918 157247 213920 157256
rect 213972 157247 213974 157256
rect 213920 157218 213972 157224
rect 214024 156913 214052 157286
rect 214010 156904 214066 156913
rect 214010 156839 214066 156848
rect 213274 155952 213330 155961
rect 213274 155887 213330 155896
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155553 213960 155858
rect 213918 155544 213974 155553
rect 213918 155479 213974 155488
rect 214010 153912 214066 153921
rect 214010 153847 214066 153856
rect 213918 153368 213974 153377
rect 213918 153303 213920 153312
rect 213972 153303 213974 153312
rect 213920 153274 213972 153280
rect 214024 153270 214052 153847
rect 214012 153264 214064 153270
rect 214012 153206 214064 153212
rect 214010 152688 214066 152697
rect 214010 152623 214066 152632
rect 213918 152008 213974 152017
rect 214024 151978 214052 152623
rect 213918 151943 213974 151952
rect 214012 151972 214064 151978
rect 213932 151910 213960 151943
rect 214012 151914 214064 151920
rect 213920 151904 213972 151910
rect 213458 151872 213514 151881
rect 213920 151846 213972 151852
rect 213458 151807 213514 151816
rect 213368 145716 213420 145722
rect 213368 145658 213420 145664
rect 213274 142352 213330 142361
rect 213274 142287 213330 142296
rect 213184 87644 213236 87650
rect 213184 87586 213236 87592
rect 213288 86902 213316 142287
rect 213380 110430 213408 145658
rect 213472 142866 213500 151807
rect 215022 150784 215078 150793
rect 215022 150719 215078 150728
rect 213918 150648 213974 150657
rect 213918 150583 213974 150592
rect 213932 150482 213960 150583
rect 213920 150476 213972 150482
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 213920 150340 213972 150346
rect 213920 150282 213972 150288
rect 213932 150113 213960 150282
rect 213918 150104 213974 150113
rect 213918 150039 213974 150048
rect 214024 149569 214052 150350
rect 214010 149560 214066 149569
rect 214010 149495 214066 149504
rect 213920 149048 213972 149054
rect 213920 148990 213972 148996
rect 213932 148889 213960 148990
rect 213918 148880 213974 148889
rect 213918 148815 213974 148824
rect 213918 148064 213974 148073
rect 213918 147999 213974 148008
rect 213932 147694 213960 147999
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 214010 146704 214066 146713
rect 214010 146639 214066 146648
rect 213918 146432 213974 146441
rect 214024 146402 214052 146639
rect 213918 146367 213974 146376
rect 214012 146396 214064 146402
rect 213932 146334 213960 146367
rect 214012 146338 214064 146344
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 215036 145722 215064 150719
rect 215024 145716 215076 145722
rect 215024 145658 215076 145664
rect 214654 145344 214710 145353
rect 214654 145279 214710 145288
rect 214010 143984 214066 143993
rect 214010 143919 214066 143928
rect 213920 143676 213972 143682
rect 213920 143618 213972 143624
rect 213932 143585 213960 143618
rect 214024 143614 214052 143919
rect 214012 143608 214064 143614
rect 213918 143576 213974 143585
rect 214012 143550 214064 143556
rect 213918 143511 213974 143520
rect 213460 142860 213512 142866
rect 213460 142802 213512 142808
rect 213918 142760 213974 142769
rect 213918 142695 213974 142704
rect 213932 142186 213960 142695
rect 213920 142180 213972 142186
rect 213920 142122 213972 142128
rect 214010 141400 214066 141409
rect 214010 141335 214066 141344
rect 214024 140894 214052 141335
rect 214012 140888 214064 140894
rect 213918 140856 213974 140865
rect 214012 140830 214064 140836
rect 213918 140791 213920 140800
rect 213972 140791 213974 140800
rect 213920 140762 213972 140768
rect 214668 140078 214696 145279
rect 214656 140072 214708 140078
rect 214562 140040 214618 140049
rect 214656 140014 214708 140020
rect 214562 139975 214618 139984
rect 213918 139496 213974 139505
rect 213918 139431 213920 139440
rect 213972 139431 213974 139440
rect 213920 139402 213972 139408
rect 214010 138816 214066 138825
rect 214010 138751 214066 138760
rect 213918 138136 213974 138145
rect 213918 138071 213920 138080
rect 213972 138071 213974 138080
rect 213920 138042 213972 138048
rect 214024 138038 214052 138751
rect 214012 138032 214064 138038
rect 214012 137974 214064 137980
rect 213918 137456 213974 137465
rect 213918 137391 213974 137400
rect 213932 136678 213960 137391
rect 214010 136776 214066 136785
rect 214010 136711 214012 136720
rect 214064 136711 214066 136720
rect 214012 136682 214064 136688
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214010 136096 214066 136105
rect 214010 136031 214066 136040
rect 213918 135416 213974 135425
rect 213918 135351 213920 135360
rect 213972 135351 213974 135360
rect 213920 135322 213972 135328
rect 214024 135318 214052 136031
rect 214012 135312 214064 135318
rect 214012 135254 214064 135260
rect 213918 134056 213974 134065
rect 213918 133991 213974 134000
rect 213932 133958 213960 133991
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 213918 132560 213974 132569
rect 213918 132495 213920 132504
rect 213972 132495 213974 132504
rect 213920 132466 213972 132472
rect 213918 131200 213974 131209
rect 213918 131135 213920 131144
rect 213972 131135 213974 131144
rect 213920 131106 213972 131112
rect 213918 129840 213974 129849
rect 213918 129775 213920 129784
rect 213972 129775 213974 129784
rect 213920 129746 213972 129752
rect 213918 128888 213974 128897
rect 213918 128823 213974 128832
rect 213932 128382 213960 128823
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 213918 127120 213974 127129
rect 213918 127055 213974 127064
rect 213932 127022 213960 127055
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 214010 126168 214066 126177
rect 214010 126103 214066 126112
rect 213918 125760 213974 125769
rect 213918 125695 213920 125704
rect 213972 125695 213974 125704
rect 213920 125666 213972 125672
rect 214024 125662 214052 126103
rect 214012 125656 214064 125662
rect 214012 125598 214064 125604
rect 214010 124808 214066 124817
rect 214010 124743 214066 124752
rect 213918 124400 213974 124409
rect 213918 124335 213974 124344
rect 213932 124302 213960 124335
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 124743
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 214010 123584 214066 123593
rect 214010 123519 214066 123528
rect 213918 123176 213974 123185
rect 213918 123111 213974 123120
rect 213932 122942 213960 123111
rect 213920 122936 213972 122942
rect 213920 122878 213972 122884
rect 214024 122874 214052 123519
rect 214012 122868 214064 122874
rect 214012 122810 214064 122816
rect 214010 122224 214066 122233
rect 214010 122159 214066 122168
rect 214024 121582 214052 122159
rect 214012 121576 214064 121582
rect 213918 121544 213974 121553
rect 214012 121518 214064 121524
rect 213918 121479 213920 121488
rect 213972 121479 213974 121488
rect 213920 121450 213972 121456
rect 213918 120864 213974 120873
rect 213918 120799 213974 120808
rect 213932 120154 213960 120799
rect 214010 120320 214066 120329
rect 214010 120255 214066 120264
rect 214024 120222 214052 120255
rect 214012 120216 214064 120222
rect 214012 120158 214064 120164
rect 213920 120148 213972 120154
rect 213920 120090 213972 120096
rect 214010 119640 214066 119649
rect 214010 119575 214066 119584
rect 213918 118960 213974 118969
rect 213918 118895 213974 118904
rect 213932 118794 213960 118895
rect 214024 118862 214052 119575
rect 214102 119096 214158 119105
rect 214102 119031 214158 119040
rect 214012 118856 214064 118862
rect 214012 118798 214064 118804
rect 213920 118788 213972 118794
rect 213920 118730 213972 118736
rect 214116 118726 214144 119031
rect 214104 118720 214156 118726
rect 214104 118662 214156 118668
rect 214010 117600 214066 117609
rect 214010 117535 214066 117544
rect 214024 117434 214052 117535
rect 214012 117428 214064 117434
rect 214012 117370 214064 117376
rect 213920 117360 213972 117366
rect 213918 117328 213920 117337
rect 213972 117328 213974 117337
rect 213918 117263 213974 117272
rect 214010 116240 214066 116249
rect 214010 116175 214066 116184
rect 214024 116074 214052 116175
rect 214012 116068 214064 116074
rect 214012 116010 214064 116016
rect 213920 116000 213972 116006
rect 213918 115968 213920 115977
rect 213972 115968 213974 115977
rect 213918 115903 213974 115912
rect 214010 115016 214066 115025
rect 214010 114951 214066 114960
rect 214024 114646 214052 114951
rect 214012 114640 214064 114646
rect 213918 114608 213974 114617
rect 214012 114582 214064 114588
rect 213918 114543 213920 114552
rect 213972 114543 213974 114552
rect 213920 114514 213972 114520
rect 214010 113656 214066 113665
rect 214010 113591 214066 113600
rect 214024 113286 214052 113591
rect 214012 113280 214064 113286
rect 213918 113248 213974 113257
rect 214012 113222 214064 113228
rect 213918 113183 213920 113192
rect 213972 113183 213974 113192
rect 213920 113154 213972 113160
rect 213458 112296 213514 112305
rect 213458 112231 213514 112240
rect 213368 110424 213420 110430
rect 213368 110366 213420 110372
rect 213276 86896 213328 86902
rect 213276 86838 213328 86844
rect 213472 85474 213500 112231
rect 213918 111888 213974 111897
rect 213918 111823 213920 111832
rect 213972 111823 213974 111832
rect 213920 111794 213972 111800
rect 214010 110936 214066 110945
rect 214010 110871 214066 110880
rect 213920 110560 213972 110566
rect 213918 110528 213920 110537
rect 213972 110528 213974 110537
rect 214024 110498 214052 110871
rect 213918 110463 213974 110472
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 213918 109304 213974 109313
rect 213918 109239 213974 109248
rect 213932 109070 213960 109239
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108352 214066 108361
rect 214010 108287 214066 108296
rect 213918 107944 213974 107953
rect 213918 107879 213974 107888
rect 213932 107710 213960 107879
rect 214024 107778 214052 108287
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 106992 214066 107001
rect 214010 106927 214066 106936
rect 213918 106448 213974 106457
rect 213918 106383 213920 106392
rect 213972 106383 213974 106392
rect 213920 106354 213972 106360
rect 214024 106350 214052 106927
rect 214012 106344 214064 106350
rect 214012 106286 214064 106292
rect 214010 105768 214066 105777
rect 214010 105703 214066 105712
rect 213918 105088 213974 105097
rect 213918 105023 213920 105032
rect 213972 105023 213974 105032
rect 213920 104994 213972 105000
rect 214024 104990 214052 105703
rect 214102 105224 214158 105233
rect 214102 105159 214158 105168
rect 214012 104984 214064 104990
rect 214012 104926 214064 104932
rect 214116 104922 214144 105159
rect 214104 104916 214156 104922
rect 214104 104858 214156 104864
rect 213918 103864 213974 103873
rect 213918 103799 213974 103808
rect 213932 103562 213960 103799
rect 213920 103556 213972 103562
rect 213920 103498 213972 103504
rect 213918 102640 213974 102649
rect 213918 102575 213974 102584
rect 213932 102202 213960 102575
rect 213920 102196 213972 102202
rect 213920 102138 213972 102144
rect 214576 101425 214604 139975
rect 214746 135552 214802 135561
rect 214746 135487 214802 135496
rect 214760 130422 214788 135487
rect 214748 130416 214800 130422
rect 214748 130358 214800 130364
rect 214654 130112 214710 130121
rect 214654 130047 214710 130056
rect 214668 102814 214696 130047
rect 214746 109712 214802 109721
rect 214746 109647 214802 109656
rect 214656 102808 214708 102814
rect 214656 102750 214708 102756
rect 214562 101416 214618 101425
rect 214562 101351 214618 101360
rect 213918 100872 213974 100881
rect 213918 100807 213974 100816
rect 213932 100774 213960 100807
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214102 99784 214158 99793
rect 214102 99719 214158 99728
rect 214010 98424 214066 98433
rect 214010 98359 214066 98368
rect 213920 98116 213972 98122
rect 213920 98058 213972 98064
rect 213932 98025 213960 98058
rect 214024 98054 214052 98359
rect 214012 98048 214064 98054
rect 213918 98016 213974 98025
rect 214012 97990 214064 97996
rect 213918 97951 213974 97960
rect 214116 95946 214144 99719
rect 214286 99512 214342 99521
rect 214286 99447 214342 99456
rect 214300 99414 214328 99447
rect 214288 99408 214340 99414
rect 214288 99350 214340 99356
rect 214654 96656 214710 96665
rect 214654 96591 214710 96600
rect 214104 95940 214156 95946
rect 214104 95882 214156 95888
rect 214562 95840 214618 95849
rect 214562 95775 214618 95784
rect 214576 86970 214604 95775
rect 214668 88330 214696 96591
rect 214656 88324 214708 88330
rect 214656 88266 214708 88272
rect 214760 88262 214788 109647
rect 214838 101144 214894 101153
rect 214838 101079 214894 101088
rect 214852 89690 214880 101079
rect 214840 89684 214892 89690
rect 214840 89626 214892 89632
rect 214748 88256 214800 88262
rect 214748 88198 214800 88204
rect 214564 86964 214616 86970
rect 214564 86906 214616 86912
rect 213460 85468 213512 85474
rect 213460 85410 213512 85416
rect 211896 82816 211948 82822
rect 211896 82758 211948 82764
rect 210516 78668 210568 78674
rect 210516 78610 210568 78616
rect 204996 51876 205048 51882
rect 204996 51818 205048 51824
rect 215956 3466 215984 347074
rect 217324 322244 217376 322250
rect 217324 322186 217376 322192
rect 216036 308508 216088 308514
rect 216036 308450 216088 308456
rect 216048 4078 216076 308450
rect 216678 97064 216734 97073
rect 216678 96999 216734 97008
rect 216692 85542 216720 96999
rect 216680 85536 216732 85542
rect 216680 85478 216732 85484
rect 216036 4072 216088 4078
rect 216036 4014 216088 4020
rect 217336 3534 217364 322186
rect 221464 305108 221516 305114
rect 221464 305050 221516 305056
rect 220084 298308 220136 298314
rect 220084 298250 220136 298256
rect 220096 180169 220124 298250
rect 220176 292664 220228 292670
rect 220176 292606 220228 292612
rect 220188 183122 220216 292606
rect 221476 192778 221504 305050
rect 226984 300212 227036 300218
rect 226984 300154 227036 300160
rect 224316 296948 224368 296954
rect 224316 296890 224368 296896
rect 224224 291848 224276 291854
rect 224224 291790 224276 291796
rect 222844 288516 222896 288522
rect 222844 288458 222896 288464
rect 221464 192772 221516 192778
rect 221464 192714 221516 192720
rect 220176 183116 220228 183122
rect 220176 183058 220228 183064
rect 220082 180160 220138 180169
rect 220082 180095 220138 180104
rect 222856 177313 222884 288458
rect 222936 274712 222988 274718
rect 222936 274654 222988 274660
rect 222948 187270 222976 274654
rect 222936 187264 222988 187270
rect 222936 187206 222988 187212
rect 224236 180033 224264 291790
rect 224328 191350 224356 296890
rect 225604 295520 225656 295526
rect 225604 295462 225656 295468
rect 224316 191344 224368 191350
rect 224316 191286 224368 191292
rect 225616 184482 225644 295462
rect 225604 184476 225656 184482
rect 225604 184418 225656 184424
rect 226996 180198 227024 300154
rect 227076 244996 227128 245002
rect 227076 244938 227128 244944
rect 227088 185842 227116 244938
rect 227076 185836 227128 185842
rect 227076 185778 227128 185784
rect 226984 180192 227036 180198
rect 226984 180134 227036 180140
rect 224222 180024 224278 180033
rect 224222 179959 224278 179968
rect 228376 177449 228404 391206
rect 286324 386436 286376 386442
rect 286324 386378 286376 386384
rect 276664 378820 276716 378826
rect 276664 378762 276716 378768
rect 272522 369064 272578 369073
rect 272522 368999 272578 369008
rect 242164 327820 242216 327826
rect 242164 327762 242216 327768
rect 228456 309256 228508 309262
rect 228456 309198 228508 309204
rect 228362 177440 228418 177449
rect 228362 177375 228418 177384
rect 222842 177304 222898 177313
rect 222842 177239 222898 177248
rect 228468 175953 228496 309198
rect 240784 306468 240836 306474
rect 240784 306410 240836 306416
rect 233884 303884 233936 303890
rect 233884 303826 233936 303832
rect 232596 302388 232648 302394
rect 232596 302330 232648 302336
rect 229744 292596 229796 292602
rect 229744 292538 229796 292544
rect 229756 187338 229784 292538
rect 231216 291372 231268 291378
rect 231216 291314 231268 291320
rect 231124 269204 231176 269210
rect 231124 269146 231176 269152
rect 229744 187332 229796 187338
rect 229744 187274 229796 187280
rect 231136 177410 231164 269146
rect 231228 243710 231256 291314
rect 232504 260908 232556 260914
rect 232504 260850 232556 260856
rect 231216 243704 231268 243710
rect 231216 243646 231268 243652
rect 231308 242956 231360 242962
rect 231308 242898 231360 242904
rect 231320 198014 231348 242898
rect 231308 198008 231360 198014
rect 231308 197950 231360 197956
rect 232516 182850 232544 260850
rect 232608 243642 232636 302330
rect 232596 243636 232648 243642
rect 232596 243578 232648 243584
rect 232596 213240 232648 213246
rect 232596 213182 232648 213188
rect 232504 182844 232556 182850
rect 232504 182786 232556 182792
rect 232608 180334 232636 213182
rect 233896 199442 233924 303826
rect 238024 301504 238076 301510
rect 238024 301446 238076 301452
rect 236644 278860 236696 278866
rect 236644 278802 236696 278808
rect 233976 270564 234028 270570
rect 233976 270506 234028 270512
rect 233884 199436 233936 199442
rect 233884 199378 233936 199384
rect 233988 181762 234016 270506
rect 235264 247172 235316 247178
rect 235264 247114 235316 247120
rect 233976 181756 234028 181762
rect 233976 181698 234028 181704
rect 232596 180328 232648 180334
rect 232596 180270 232648 180276
rect 235276 179042 235304 247114
rect 236656 180402 236684 278802
rect 238036 213246 238064 301446
rect 238116 240236 238168 240242
rect 238116 240178 238168 240184
rect 238024 213240 238076 213246
rect 238024 213182 238076 213188
rect 238024 198076 238076 198082
rect 238024 198018 238076 198024
rect 236644 180396 236696 180402
rect 236644 180338 236696 180344
rect 235264 179036 235316 179042
rect 235264 178978 235316 178984
rect 238036 177585 238064 198018
rect 238128 178974 238156 240178
rect 239404 235408 239456 235414
rect 239404 235350 239456 235356
rect 238116 178968 238168 178974
rect 238116 178910 238168 178916
rect 238022 177576 238078 177585
rect 238022 177511 238078 177520
rect 231124 177404 231176 177410
rect 231124 177346 231176 177352
rect 239416 175982 239444 235350
rect 240796 183190 240824 306410
rect 240876 280288 240928 280294
rect 240876 280230 240928 280236
rect 240784 183184 240836 183190
rect 240784 183126 240836 183132
rect 240888 177478 240916 280230
rect 242176 181393 242204 327762
rect 265624 323672 265676 323678
rect 265624 323614 265676 323620
rect 246304 298240 246356 298246
rect 246304 298182 246356 298188
rect 244924 295452 244976 295458
rect 244924 295394 244976 295400
rect 243544 249824 243596 249830
rect 243544 249766 243596 249772
rect 242162 181384 242218 181393
rect 242162 181319 242218 181328
rect 243556 178022 243584 249766
rect 243544 178016 243596 178022
rect 243544 177958 243596 177964
rect 240876 177472 240928 177478
rect 240876 177414 240928 177420
rect 244936 176118 244964 295394
rect 245016 259480 245068 259486
rect 245016 259422 245068 259428
rect 244924 176112 244976 176118
rect 244924 176054 244976 176060
rect 245028 176050 245056 259422
rect 245384 183048 245436 183054
rect 245384 182990 245436 182996
rect 245396 177954 245424 182990
rect 245384 177948 245436 177954
rect 245384 177890 245436 177896
rect 246316 177546 246344 298182
rect 249800 296880 249852 296886
rect 249800 296822 249852 296828
rect 246396 281648 246448 281654
rect 246396 281590 246448 281596
rect 246408 180470 246436 281590
rect 249064 281580 249116 281586
rect 249064 281522 249116 281528
rect 246488 217388 246540 217394
rect 246488 217330 246540 217336
rect 246396 180464 246448 180470
rect 246396 180406 246448 180412
rect 246304 177540 246356 177546
rect 246304 177482 246356 177488
rect 246500 176633 246528 217330
rect 249076 190058 249104 281522
rect 249064 190052 249116 190058
rect 249064 189994 249116 190000
rect 249340 188488 249392 188494
rect 249340 188430 249392 188436
rect 247684 185700 247736 185706
rect 247684 185642 247736 185648
rect 247696 178673 247724 185642
rect 249064 180464 249116 180470
rect 249064 180406 249116 180412
rect 247682 178664 247738 178673
rect 247682 178599 247738 178608
rect 246486 176624 246542 176633
rect 246486 176559 246542 176568
rect 245016 176044 245068 176050
rect 245016 175986 245068 175992
rect 239404 175976 239456 175982
rect 228454 175944 228510 175953
rect 239404 175918 239456 175924
rect 228454 175879 228510 175888
rect 249076 174690 249104 180406
rect 249156 178016 249208 178022
rect 249156 177958 249208 177964
rect 249168 175273 249196 177958
rect 249248 177948 249300 177954
rect 249248 177890 249300 177896
rect 249154 175264 249210 175273
rect 249154 175199 249210 175208
rect 249154 174704 249210 174713
rect 249076 174662 249154 174690
rect 249154 174639 249210 174648
rect 249260 173369 249288 177890
rect 249352 175681 249380 188430
rect 249432 180396 249484 180402
rect 249432 180338 249484 180344
rect 249338 175672 249394 175681
rect 249338 175607 249394 175616
rect 249246 173360 249302 173369
rect 249246 173295 249302 173304
rect 249444 172825 249472 180338
rect 249430 172816 249486 172825
rect 249430 172751 249486 172760
rect 249812 168201 249840 296822
rect 251824 296812 251876 296818
rect 251824 296754 251876 296760
rect 251836 235414 251864 296754
rect 251916 272604 251968 272610
rect 251916 272546 251968 272552
rect 251928 238270 251956 272546
rect 252560 269136 252612 269142
rect 252560 269078 252612 269084
rect 251916 238264 251968 238270
rect 251916 238206 251968 238212
rect 251824 235408 251876 235414
rect 251824 235350 251876 235356
rect 251272 234048 251324 234054
rect 251272 233990 251324 233996
rect 251180 225684 251232 225690
rect 251180 225626 251232 225632
rect 249892 207800 249944 207806
rect 249892 207742 249944 207748
rect 249798 168192 249854 168201
rect 249798 168127 249854 168136
rect 249904 154465 249932 207742
rect 249984 199640 250036 199646
rect 249984 199582 250036 199588
rect 249996 160585 250024 199582
rect 250076 179036 250128 179042
rect 250076 178978 250128 178984
rect 250088 171465 250116 178978
rect 250074 171456 250130 171465
rect 250074 171391 250130 171400
rect 250444 162240 250496 162246
rect 250444 162182 250496 162188
rect 249982 160576 250038 160585
rect 249982 160511 250038 160520
rect 249890 154456 249946 154465
rect 249890 154391 249946 154400
rect 250456 144673 250484 162182
rect 250536 162172 250588 162178
rect 250536 162114 250588 162120
rect 250442 144664 250498 144673
rect 250442 144599 250498 144608
rect 249064 138032 249116 138038
rect 249064 137974 249116 137980
rect 246486 94480 246542 94489
rect 246486 94415 246542 94424
rect 232504 93152 232556 93158
rect 232504 93094 232556 93100
rect 232516 7682 232544 93094
rect 238024 91860 238076 91866
rect 238024 91802 238076 91808
rect 232504 7676 232556 7682
rect 232504 7618 232556 7624
rect 217324 3528 217376 3534
rect 217324 3470 217376 3476
rect 202236 3460 202288 3466
rect 202236 3402 202288 3408
rect 215944 3460 215996 3466
rect 215944 3402 215996 3408
rect 238036 3058 238064 91802
rect 246304 79416 246356 79422
rect 246304 79358 246356 79364
rect 243544 54596 243596 54602
rect 243544 54538 243596 54544
rect 240784 53168 240836 53174
rect 240784 53110 240836 53116
rect 240796 4078 240824 53110
rect 241520 51876 241572 51882
rect 241520 51818 241572 51824
rect 241532 16574 241560 51818
rect 241532 16546 241744 16574
rect 240508 4072 240560 4078
rect 240508 4014 240560 4020
rect 240784 4072 240836 4078
rect 240784 4014 240836 4020
rect 239312 3460 239364 3466
rect 239312 3402 239364 3408
rect 235816 3052 235868 3058
rect 235816 2994 235868 3000
rect 238024 3052 238076 3058
rect 238024 2994 238076 3000
rect 235828 480 235856 2994
rect 239324 480 239352 3402
rect 240520 480 240548 4014
rect 241716 480 241744 16546
rect 243556 10985 243584 54538
rect 244280 50584 244332 50590
rect 244280 50526 244332 50532
rect 244292 49706 244320 50526
rect 244280 49700 244332 49706
rect 244280 49642 244332 49648
rect 244292 16574 244320 49642
rect 246316 20670 246344 79358
rect 246394 77888 246450 77897
rect 246394 77823 246450 77832
rect 246408 57254 246436 77823
rect 246500 73914 246528 94415
rect 246488 73908 246540 73914
rect 246488 73850 246540 73856
rect 246396 57248 246448 57254
rect 246396 57190 246448 57196
rect 249076 51814 249104 137974
rect 250548 136649 250576 162114
rect 250628 159452 250680 159458
rect 250628 159394 250680 159400
rect 250640 144129 250668 159394
rect 250810 153776 250866 153785
rect 250810 153711 250866 153720
rect 250720 144220 250772 144226
rect 250720 144162 250772 144168
rect 250626 144120 250682 144129
rect 250626 144055 250682 144064
rect 250628 136672 250680 136678
rect 250534 136640 250590 136649
rect 250628 136614 250680 136620
rect 250534 136575 250590 136584
rect 250444 135312 250496 135318
rect 250444 135254 250496 135260
rect 249248 98048 249300 98054
rect 249248 97990 249300 97996
rect 249156 78056 249208 78062
rect 249156 77998 249208 78004
rect 249064 51808 249116 51814
rect 249064 51750 249116 51756
rect 246304 20664 246356 20670
rect 246304 20606 246356 20612
rect 249168 20602 249196 77998
rect 249260 50386 249288 97990
rect 249798 97064 249854 97073
rect 249798 96999 249854 97008
rect 249248 50380 249300 50386
rect 249248 50322 249300 50328
rect 249812 23458 249840 96999
rect 250456 45014 250484 135254
rect 250536 120216 250588 120222
rect 250536 120158 250588 120164
rect 250444 45008 250496 45014
rect 250444 44950 250496 44956
rect 250548 32502 250576 120158
rect 250640 54738 250668 136614
rect 250732 106049 250760 144162
rect 250824 141817 250852 153711
rect 251192 147937 251220 225626
rect 251284 157865 251312 233990
rect 251364 229900 251416 229906
rect 251364 229842 251416 229848
rect 251270 157856 251326 157865
rect 251270 157791 251326 157800
rect 251376 156369 251404 229842
rect 252468 172508 252520 172514
rect 252468 172450 252520 172456
rect 252376 172440 252428 172446
rect 252480 172417 252508 172450
rect 252376 172382 252428 172388
rect 252466 172408 252522 172417
rect 252388 171873 252416 172382
rect 252466 172343 252522 172352
rect 252374 171864 252430 171873
rect 252374 171799 252430 171808
rect 252376 171080 252428 171086
rect 252376 171022 252428 171028
rect 252388 170513 252416 171022
rect 252468 171012 252520 171018
rect 252468 170954 252520 170960
rect 252480 170921 252508 170954
rect 252466 170912 252522 170921
rect 252466 170847 252522 170856
rect 252374 170504 252430 170513
rect 252374 170439 252430 170448
rect 252468 170128 252520 170134
rect 252466 170096 252468 170105
rect 252520 170096 252522 170105
rect 252466 170031 252522 170040
rect 252468 169652 252520 169658
rect 252468 169594 252520 169600
rect 252376 169584 252428 169590
rect 252376 169526 252428 169532
rect 252388 168609 252416 169526
rect 252480 169153 252508 169594
rect 252466 169144 252522 169153
rect 252466 169079 252522 169088
rect 252374 168600 252430 168609
rect 252374 168535 252430 168544
rect 252376 168360 252428 168366
rect 252376 168302 252428 168308
rect 252388 167657 252416 168302
rect 252468 167952 252520 167958
rect 252468 167894 252520 167900
rect 252374 167648 252430 167657
rect 252374 167583 252430 167592
rect 252480 167249 252508 167894
rect 252466 167240 252522 167249
rect 252466 167175 252522 167184
rect 252466 166696 252522 166705
rect 252466 166631 252522 166640
rect 252480 166394 252508 166631
rect 252468 166388 252520 166394
rect 252468 166330 252520 166336
rect 252468 166116 252520 166122
rect 252468 166058 252520 166064
rect 252480 165753 252508 166058
rect 252466 165744 252522 165753
rect 252466 165679 252522 165688
rect 252284 165572 252336 165578
rect 252284 165514 252336 165520
rect 252296 164801 252324 165514
rect 252468 165504 252520 165510
rect 252468 165446 252520 165452
rect 252376 165436 252428 165442
rect 252376 165378 252428 165384
rect 252282 164792 252338 164801
rect 252282 164727 252338 164736
rect 252388 164393 252416 165378
rect 252480 165345 252508 165446
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 252374 164384 252430 164393
rect 252374 164319 252430 164328
rect 252376 164212 252428 164218
rect 252376 164154 252428 164160
rect 252284 164144 252336 164150
rect 252284 164086 252336 164092
rect 252296 163033 252324 164086
rect 252388 163441 252416 164154
rect 252468 164076 252520 164082
rect 252468 164018 252520 164024
rect 252480 163985 252508 164018
rect 252466 163976 252522 163985
rect 252466 163911 252522 163920
rect 252374 163432 252430 163441
rect 252374 163367 252430 163376
rect 252282 163024 252338 163033
rect 252282 162959 252338 162968
rect 252376 162852 252428 162858
rect 252376 162794 252428 162800
rect 252388 161537 252416 162794
rect 252468 162784 252520 162790
rect 252468 162726 252520 162732
rect 252480 162081 252508 162726
rect 252572 162489 252600 269078
rect 260840 256760 260892 256766
rect 260840 256702 260892 256708
rect 258080 252680 258132 252686
rect 258080 252622 258132 252628
rect 255412 227112 255464 227118
rect 255412 227054 255464 227060
rect 252652 209228 252704 209234
rect 252652 209170 252704 209176
rect 252558 162480 252614 162489
rect 252558 162415 252614 162424
rect 252466 162072 252522 162081
rect 252466 162007 252522 162016
rect 252374 161528 252430 161537
rect 252374 161463 252430 161472
rect 252468 161424 252520 161430
rect 252468 161366 252520 161372
rect 252480 160313 252508 161366
rect 252466 160304 252522 160313
rect 252466 160239 252522 160248
rect 252468 160064 252520 160070
rect 252468 160006 252520 160012
rect 251732 159996 251784 160002
rect 251732 159938 251784 159944
rect 251744 159633 251772 159938
rect 251730 159624 251786 159633
rect 251730 159559 251786 159568
rect 252480 158817 252508 160006
rect 252466 158808 252522 158817
rect 252466 158743 252522 158752
rect 252468 158704 252520 158710
rect 252468 158646 252520 158652
rect 252480 158273 252508 158646
rect 252466 158264 252522 158273
rect 252466 158199 252522 158208
rect 251824 158092 251876 158098
rect 251824 158034 251876 158040
rect 251362 156360 251418 156369
rect 251362 156295 251418 156304
rect 251178 147928 251234 147937
rect 251178 147863 251234 147872
rect 251456 147484 251508 147490
rect 251456 147426 251508 147432
rect 251468 146985 251496 147426
rect 251454 146976 251510 146985
rect 251454 146911 251510 146920
rect 251180 146124 251232 146130
rect 251180 146066 251232 146072
rect 251192 145081 251220 146066
rect 251178 145072 251234 145081
rect 251178 145007 251234 145016
rect 250810 141808 250866 141817
rect 250810 141743 250866 141752
rect 251180 141568 251232 141574
rect 251180 141510 251232 141516
rect 251192 140865 251220 141510
rect 251178 140856 251234 140865
rect 251178 140791 251234 140800
rect 251836 138553 251864 158034
rect 252468 157344 252520 157350
rect 252468 157286 252520 157292
rect 252480 156913 252508 157286
rect 252466 156904 252522 156913
rect 252466 156839 252522 156848
rect 252664 155961 252692 209170
rect 254216 203788 254268 203794
rect 254216 203730 254268 203736
rect 254032 196852 254084 196858
rect 254032 196794 254084 196800
rect 252836 193928 252888 193934
rect 252836 193870 252888 193876
rect 252744 182980 252796 182986
rect 252744 182922 252796 182928
rect 252650 155952 252706 155961
rect 252376 155916 252428 155922
rect 252650 155887 252706 155896
rect 252376 155858 252428 155864
rect 252388 155009 252416 155858
rect 252468 155848 252520 155854
rect 252468 155790 252520 155796
rect 252480 155417 252508 155790
rect 252466 155408 252522 155417
rect 252466 155343 252522 155352
rect 252374 155000 252430 155009
rect 252374 154935 252430 154944
rect 252468 154556 252520 154562
rect 252468 154498 252520 154504
rect 252100 154488 252152 154494
rect 252100 154430 252152 154436
rect 252112 153513 252140 154430
rect 252480 154057 252508 154498
rect 252466 154048 252522 154057
rect 252466 153983 252522 153992
rect 252098 153504 252154 153513
rect 252098 153439 252154 153448
rect 252284 153196 252336 153202
rect 252284 153138 252336 153144
rect 252296 153105 252324 153138
rect 252376 153128 252428 153134
rect 252282 153096 252338 153105
rect 252376 153070 252428 153076
rect 252282 153031 252338 153040
rect 252388 152153 252416 153070
rect 252468 153060 252520 153066
rect 252468 153002 252520 153008
rect 252480 152697 252508 153002
rect 252466 152688 252522 152697
rect 252466 152623 252522 152632
rect 252374 152144 252430 152153
rect 252374 152079 252430 152088
rect 252468 151768 252520 151774
rect 252466 151736 252468 151745
rect 252520 151736 252522 151745
rect 252466 151671 252522 151680
rect 252468 151496 252520 151502
rect 252468 151438 252520 151444
rect 252284 151292 252336 151298
rect 252284 151234 252336 151240
rect 252296 150793 252324 151234
rect 252480 151201 252508 151438
rect 252466 151192 252522 151201
rect 252466 151127 252522 151136
rect 252282 150784 252338 150793
rect 252282 150719 252338 150728
rect 252376 150408 252428 150414
rect 252376 150350 252428 150356
rect 252284 150272 252336 150278
rect 252284 150214 252336 150220
rect 252296 149841 252324 150214
rect 252282 149832 252338 149841
rect 252282 149767 252338 149776
rect 252388 149297 252416 150350
rect 252468 150340 252520 150346
rect 252468 150282 252520 150288
rect 252480 150249 252508 150282
rect 252466 150240 252522 150249
rect 252466 150175 252522 150184
rect 252374 149288 252430 149297
rect 252374 149223 252430 149232
rect 252468 149048 252520 149054
rect 252468 148990 252520 148996
rect 252376 148980 252428 148986
rect 252376 148922 252428 148928
rect 252388 148345 252416 148922
rect 252480 148889 252508 148990
rect 252466 148880 252522 148889
rect 252466 148815 252522 148824
rect 252374 148336 252430 148345
rect 252374 148271 252430 148280
rect 252376 147620 252428 147626
rect 252376 147562 252428 147568
rect 252388 146577 252416 147562
rect 252468 147552 252520 147558
rect 252466 147520 252468 147529
rect 252520 147520 252522 147529
rect 252466 147455 252522 147464
rect 252374 146568 252430 146577
rect 252374 146503 252430 146512
rect 252468 146260 252520 146266
rect 252468 146202 252520 146208
rect 252376 146192 252428 146198
rect 252376 146134 252428 146140
rect 252388 145625 252416 146134
rect 252480 146033 252508 146202
rect 252466 146024 252522 146033
rect 252466 145959 252522 145968
rect 252374 145616 252430 145625
rect 252374 145551 252430 145560
rect 252468 144900 252520 144906
rect 252468 144842 252520 144848
rect 252100 144356 252152 144362
rect 252100 144298 252152 144304
rect 252008 141432 252060 141438
rect 252008 141374 252060 141380
rect 251916 140004 251968 140010
rect 251916 139946 251968 139952
rect 251822 138544 251878 138553
rect 251822 138479 251878 138488
rect 251824 124908 251876 124914
rect 251824 124850 251876 124856
rect 251180 111784 251232 111790
rect 251180 111726 251232 111732
rect 251192 111217 251220 111726
rect 251178 111208 251234 111217
rect 251178 111143 251234 111152
rect 251732 110424 251784 110430
rect 251732 110366 251784 110372
rect 251744 109313 251772 110366
rect 251730 109304 251786 109313
rect 251730 109239 251786 109248
rect 250718 106040 250774 106049
rect 250718 105975 250774 105984
rect 251364 105664 251416 105670
rect 251364 105606 251416 105612
rect 251376 98025 251404 105606
rect 251732 102876 251784 102882
rect 251732 102818 251784 102824
rect 251744 101425 251772 102818
rect 251836 102785 251864 124850
rect 251928 120193 251956 139946
rect 252020 124817 252048 141374
rect 252112 131481 252140 144298
rect 252480 143721 252508 144842
rect 252466 143712 252522 143721
rect 252466 143647 252522 143656
rect 252468 143540 252520 143546
rect 252468 143482 252520 143488
rect 252376 143472 252428 143478
rect 252376 143414 252428 143420
rect 252388 142769 252416 143414
rect 252480 143177 252508 143482
rect 252466 143168 252522 143177
rect 252466 143103 252522 143112
rect 252374 142760 252430 142769
rect 252374 142695 252430 142704
rect 252756 142154 252784 182922
rect 252848 169561 252876 193870
rect 252834 169552 252890 169561
rect 252834 169487 252890 169496
rect 253296 163532 253348 163538
rect 253296 163474 253348 163480
rect 253204 152516 253256 152522
rect 253204 152458 253256 152464
rect 252572 142126 252784 142154
rect 252468 142112 252520 142118
rect 252468 142054 252520 142060
rect 252480 141409 252508 142054
rect 252466 141400 252522 141409
rect 252466 141335 252522 141344
rect 252468 140752 252520 140758
rect 252468 140694 252520 140700
rect 252376 140684 252428 140690
rect 252376 140626 252428 140632
rect 252388 139913 252416 140626
rect 252480 140457 252508 140694
rect 252466 140448 252522 140457
rect 252466 140383 252522 140392
rect 252374 139904 252430 139913
rect 252374 139839 252430 139848
rect 252572 139505 252600 142126
rect 252558 139496 252614 139505
rect 252558 139431 252614 139440
rect 252468 139392 252520 139398
rect 252468 139334 252520 139340
rect 252480 138961 252508 139334
rect 252466 138952 252522 138961
rect 252466 138887 252522 138896
rect 252466 138000 252522 138009
rect 252466 137935 252468 137944
rect 252520 137935 252522 137944
rect 252468 137906 252520 137912
rect 252192 137284 252244 137290
rect 252192 137226 252244 137232
rect 252098 131472 252154 131481
rect 252098 131407 252154 131416
rect 252100 124976 252152 124982
rect 252100 124918 252152 124924
rect 252006 124808 252062 124817
rect 252006 124743 252062 124752
rect 252112 121145 252140 124918
rect 252204 124409 252232 137226
rect 252284 136604 252336 136610
rect 252284 136546 252336 136552
rect 252296 135289 252324 136546
rect 252468 136536 252520 136542
rect 252468 136478 252520 136484
rect 252376 136468 252428 136474
rect 252376 136410 252428 136416
rect 252388 135697 252416 136410
rect 252480 136241 252508 136478
rect 252466 136232 252522 136241
rect 252466 136167 252522 136176
rect 252374 135688 252430 135697
rect 252374 135623 252430 135632
rect 252282 135280 252338 135289
rect 252282 135215 252338 135224
rect 252468 135244 252520 135250
rect 252468 135186 252520 135192
rect 252376 135176 252428 135182
rect 252376 135118 252428 135124
rect 252388 134337 252416 135118
rect 252480 134745 252508 135186
rect 252466 134736 252522 134745
rect 252466 134671 252522 134680
rect 252374 134328 252430 134337
rect 252374 134263 252430 134272
rect 252284 133884 252336 133890
rect 252284 133826 252336 133832
rect 252296 132841 252324 133826
rect 252376 133816 252428 133822
rect 252376 133758 252428 133764
rect 252466 133784 252522 133793
rect 252388 133385 252416 133758
rect 252466 133719 252468 133728
rect 252520 133719 252522 133728
rect 252468 133690 252520 133696
rect 252374 133376 252430 133385
rect 252374 133311 252430 133320
rect 252282 132832 252338 132841
rect 252282 132767 252338 132776
rect 252376 132456 252428 132462
rect 252376 132398 252428 132404
rect 252466 132424 252522 132433
rect 252388 131889 252416 132398
rect 252466 132359 252468 132368
rect 252520 132359 252522 132368
rect 252468 132330 252520 132336
rect 252374 131880 252430 131889
rect 252374 131815 252430 131824
rect 252376 131096 252428 131102
rect 252376 131038 252428 131044
rect 252284 131028 252336 131034
rect 252284 130970 252336 130976
rect 252296 130121 252324 130970
rect 252388 130937 252416 131038
rect 252468 130960 252520 130966
rect 252374 130928 252430 130937
rect 252468 130902 252520 130908
rect 252374 130863 252430 130872
rect 252480 130529 252508 130902
rect 252466 130520 252522 130529
rect 252466 130455 252522 130464
rect 252282 130112 252338 130121
rect 252282 130047 252338 130056
rect 252468 129736 252520 129742
rect 252468 129678 252520 129684
rect 252376 129668 252428 129674
rect 252376 129610 252428 129616
rect 252284 129600 252336 129606
rect 252284 129542 252336 129548
rect 252296 128625 252324 129542
rect 252388 129169 252416 129610
rect 252480 129577 252508 129678
rect 252466 129568 252522 129577
rect 252466 129503 252522 129512
rect 252374 129160 252430 129169
rect 252374 129095 252430 129104
rect 252282 128616 252338 128625
rect 252282 128551 252338 128560
rect 252468 128308 252520 128314
rect 252468 128250 252520 128256
rect 252284 128240 252336 128246
rect 252480 128217 252508 128250
rect 252284 128182 252336 128188
rect 252466 128208 252522 128217
rect 252296 127673 252324 128182
rect 252376 128172 252428 128178
rect 252466 128143 252522 128152
rect 252376 128114 252428 128120
rect 252282 127664 252338 127673
rect 252282 127599 252338 127608
rect 252388 127265 252416 128114
rect 252374 127256 252430 127265
rect 252374 127191 252430 127200
rect 252284 126948 252336 126954
rect 252284 126890 252336 126896
rect 252296 125769 252324 126890
rect 252468 126880 252520 126886
rect 252468 126822 252520 126828
rect 252376 126812 252428 126818
rect 252376 126754 252428 126760
rect 252388 126313 252416 126754
rect 252480 126721 252508 126822
rect 252466 126712 252522 126721
rect 252466 126647 252522 126656
rect 252374 126304 252430 126313
rect 252374 126239 252430 126248
rect 252282 125760 252338 125769
rect 252282 125695 252338 125704
rect 252468 125588 252520 125594
rect 252468 125530 252520 125536
rect 252480 125361 252508 125530
rect 252466 125352 252522 125361
rect 252466 125287 252522 125296
rect 252190 124400 252246 124409
rect 252190 124335 252246 124344
rect 252376 124160 252428 124166
rect 252376 124102 252428 124108
rect 252284 124024 252336 124030
rect 252284 123966 252336 123972
rect 252296 123049 252324 123966
rect 252388 123457 252416 124102
rect 252468 124092 252520 124098
rect 252468 124034 252520 124040
rect 252480 124001 252508 124034
rect 252466 123992 252522 124001
rect 252466 123927 252522 123936
rect 252374 123448 252430 123457
rect 252374 123383 252430 123392
rect 252282 123040 252338 123049
rect 252282 122975 252338 122984
rect 252468 122800 252520 122806
rect 252468 122742 252520 122748
rect 252376 122732 252428 122738
rect 252376 122674 252428 122680
rect 252284 122664 252336 122670
rect 252284 122606 252336 122612
rect 252296 121553 252324 122606
rect 252388 122097 252416 122674
rect 252480 122505 252508 122742
rect 252466 122496 252522 122505
rect 252466 122431 252522 122440
rect 252374 122088 252430 122097
rect 252374 122023 252430 122032
rect 252282 121544 252338 121553
rect 252282 121479 252338 121488
rect 252468 121440 252520 121446
rect 252468 121382 252520 121388
rect 252098 121136 252154 121145
rect 252098 121071 252154 121080
rect 252480 120601 252508 121382
rect 252466 120592 252522 120601
rect 252466 120527 252522 120536
rect 251914 120184 251970 120193
rect 251914 120119 251970 120128
rect 252008 120148 252060 120154
rect 252008 120090 252060 120096
rect 251916 116612 251968 116618
rect 251916 116554 251968 116560
rect 251928 107953 251956 116554
rect 251914 107944 251970 107953
rect 251914 107879 251970 107888
rect 252020 105097 252048 120090
rect 252284 120080 252336 120086
rect 252284 120022 252336 120028
rect 252296 119241 252324 120022
rect 252468 120012 252520 120018
rect 252468 119954 252520 119960
rect 252376 119876 252428 119882
rect 252376 119818 252428 119824
rect 252282 119232 252338 119241
rect 252282 119167 252338 119176
rect 252388 118833 252416 119818
rect 252480 119649 252508 119954
rect 252466 119640 252522 119649
rect 252466 119575 252522 119584
rect 252374 118824 252430 118833
rect 252374 118759 252430 118768
rect 252376 118652 252428 118658
rect 252376 118594 252428 118600
rect 252284 118584 252336 118590
rect 252284 118526 252336 118532
rect 252296 117337 252324 118526
rect 252388 117881 252416 118594
rect 252466 118280 252522 118289
rect 252466 118215 252522 118224
rect 252374 117872 252430 117881
rect 252374 117807 252430 117816
rect 252480 117706 252508 118215
rect 252468 117700 252520 117706
rect 252468 117642 252520 117648
rect 252282 117328 252338 117337
rect 252282 117263 252338 117272
rect 252468 117292 252520 117298
rect 252468 117234 252520 117240
rect 252376 117224 252428 117230
rect 252376 117166 252428 117172
rect 252388 115977 252416 117166
rect 252480 116385 252508 117234
rect 252466 116376 252522 116385
rect 252466 116311 252522 116320
rect 252374 115968 252430 115977
rect 252374 115903 252430 115912
rect 252468 115932 252520 115938
rect 252468 115874 252520 115880
rect 252376 115864 252428 115870
rect 252376 115806 252428 115812
rect 252284 115252 252336 115258
rect 252284 115194 252336 115200
rect 252296 113529 252324 115194
rect 252388 115025 252416 115806
rect 252480 115433 252508 115874
rect 252466 115424 252522 115433
rect 252466 115359 252522 115368
rect 252374 115016 252430 115025
rect 252374 114951 252430 114960
rect 252468 114504 252520 114510
rect 252466 114472 252468 114481
rect 252520 114472 252522 114481
rect 252466 114407 252522 114416
rect 253216 114073 253244 152458
rect 253308 141574 253336 163474
rect 253480 159384 253532 159390
rect 253480 159326 253532 159332
rect 253492 146130 253520 159326
rect 253940 155236 253992 155242
rect 253940 155178 253992 155184
rect 253952 153202 253980 155178
rect 253940 153196 253992 153202
rect 253940 153138 253992 153144
rect 254044 151774 254072 196794
rect 254124 176112 254176 176118
rect 254124 176054 254176 176060
rect 254136 160002 254164 176054
rect 254124 159996 254176 160002
rect 254124 159938 254176 159944
rect 254032 151768 254084 151774
rect 254032 151710 254084 151716
rect 254228 147490 254256 203730
rect 255424 154494 255452 227054
rect 255596 224324 255648 224330
rect 255596 224266 255648 224272
rect 255504 202292 255556 202298
rect 255504 202234 255556 202240
rect 255412 154488 255464 154494
rect 255412 154430 255464 154436
rect 255516 151298 255544 202234
rect 255608 151502 255636 224266
rect 256700 187332 256752 187338
rect 256700 187274 256752 187280
rect 256240 153876 256292 153882
rect 256240 153818 256292 153824
rect 255596 151496 255648 151502
rect 255596 151438 255648 151444
rect 255504 151292 255556 151298
rect 255504 151234 255556 151240
rect 255964 150544 256016 150550
rect 255964 150486 256016 150492
rect 254676 150476 254728 150482
rect 254676 150418 254728 150424
rect 254216 147484 254268 147490
rect 254216 147426 254268 147432
rect 253480 146124 253532 146130
rect 253480 146066 253532 146072
rect 253388 145580 253440 145586
rect 253388 145522 253440 145528
rect 253296 141568 253348 141574
rect 253296 141510 253348 141516
rect 253296 138100 253348 138106
rect 253296 138042 253348 138048
rect 253202 114064 253258 114073
rect 253202 113999 253258 114008
rect 252376 113824 252428 113830
rect 252376 113766 252428 113772
rect 252282 113520 252338 113529
rect 252282 113455 252338 113464
rect 252282 113112 252338 113121
rect 252282 113047 252284 113056
rect 252336 113047 252338 113056
rect 252284 113018 252336 113024
rect 252388 112713 252416 113766
rect 252468 113144 252520 113150
rect 252468 113086 252520 113092
rect 252374 112704 252430 112713
rect 252374 112639 252430 112648
rect 252284 112464 252336 112470
rect 252284 112406 252336 112412
rect 252296 105641 252324 112406
rect 252480 112169 252508 113086
rect 252466 112160 252522 112169
rect 252466 112095 252522 112104
rect 252374 111752 252430 111761
rect 252374 111687 252376 111696
rect 252428 111687 252430 111696
rect 252376 111658 252428 111664
rect 252468 111648 252520 111654
rect 252468 111590 252520 111596
rect 252480 110809 252508 111590
rect 252466 110800 252522 110809
rect 252466 110735 252522 110744
rect 252468 110356 252520 110362
rect 252468 110298 252520 110304
rect 252480 110265 252508 110298
rect 252466 110256 252522 110265
rect 252466 110191 252522 110200
rect 253204 109064 253256 109070
rect 253204 109006 253256 109012
rect 252376 108996 252428 109002
rect 252376 108938 252428 108944
rect 252388 108361 252416 108938
rect 252468 108928 252520 108934
rect 252466 108896 252468 108905
rect 252520 108896 252522 108905
rect 252466 108831 252522 108840
rect 252374 108352 252430 108361
rect 252374 108287 252430 108296
rect 252468 107636 252520 107642
rect 252468 107578 252520 107584
rect 252376 107568 252428 107574
rect 252480 107545 252508 107578
rect 252376 107510 252428 107516
rect 252466 107536 252522 107545
rect 252388 107001 252416 107510
rect 252466 107471 252522 107480
rect 252374 106992 252430 107001
rect 252374 106927 252430 106936
rect 252468 106956 252520 106962
rect 252468 106898 252520 106904
rect 252480 106593 252508 106898
rect 252466 106584 252522 106593
rect 252466 106519 252522 106528
rect 252282 105632 252338 105641
rect 252282 105567 252338 105576
rect 252376 105596 252428 105602
rect 252376 105538 252428 105544
rect 252006 105088 252062 105097
rect 252006 105023 252062 105032
rect 252284 104780 252336 104786
rect 252284 104722 252336 104728
rect 252296 104689 252324 104722
rect 252282 104680 252338 104689
rect 252282 104615 252338 104624
rect 252388 104145 252416 105538
rect 252468 104848 252520 104854
rect 252468 104790 252520 104796
rect 252374 104136 252430 104145
rect 252374 104071 252430 104080
rect 252480 103737 252508 104790
rect 252466 103728 252522 103737
rect 252466 103663 252522 103672
rect 252376 103488 252428 103494
rect 252376 103430 252428 103436
rect 251822 102776 251878 102785
rect 251822 102711 251878 102720
rect 252388 102241 252416 103430
rect 252466 103184 252522 103193
rect 252466 103119 252522 103128
rect 252480 102610 252508 103119
rect 252468 102604 252520 102610
rect 252468 102546 252520 102552
rect 252374 102232 252430 102241
rect 252374 102167 252430 102176
rect 252468 102128 252520 102134
rect 252468 102070 252520 102076
rect 252376 102060 252428 102066
rect 252376 102002 252428 102008
rect 252192 101448 252244 101454
rect 251730 101416 251786 101425
rect 252192 101390 252244 101396
rect 251730 101351 251786 101360
rect 251362 98016 251418 98025
rect 251362 97951 251418 97960
rect 252204 97617 252232 101390
rect 252388 100881 252416 102002
rect 252480 101833 252508 102070
rect 252466 101824 252522 101833
rect 252466 101759 252522 101768
rect 252374 100872 252430 100881
rect 252374 100807 252430 100816
rect 252284 100700 252336 100706
rect 252284 100642 252336 100648
rect 252296 99929 252324 100642
rect 252468 100632 252520 100638
rect 252468 100574 252520 100580
rect 252376 100564 252428 100570
rect 252376 100506 252428 100512
rect 252282 99920 252338 99929
rect 252282 99855 252338 99864
rect 252388 99521 252416 100506
rect 252480 100473 252508 100574
rect 252466 100464 252522 100473
rect 252466 100399 252522 100408
rect 252374 99512 252430 99521
rect 252374 99447 252430 99456
rect 252376 99340 252428 99346
rect 252376 99282 252428 99288
rect 252388 98569 252416 99282
rect 252468 99272 252520 99278
rect 252468 99214 252520 99220
rect 252480 98977 252508 99214
rect 252466 98968 252522 98977
rect 252466 98903 252522 98912
rect 252374 98560 252430 98569
rect 252374 98495 252430 98504
rect 252190 97608 252246 97617
rect 252190 97543 252246 97552
rect 252466 97336 252522 97345
rect 252466 97271 252522 97280
rect 252480 96665 252508 97271
rect 252466 96656 252522 96665
rect 252466 96591 252522 96600
rect 251178 96248 251234 96257
rect 251178 96183 251234 96192
rect 251192 91866 251220 96183
rect 251824 95260 251876 95266
rect 251824 95202 251876 95208
rect 251180 91860 251232 91866
rect 251180 91802 251232 91808
rect 251178 86184 251234 86193
rect 251178 86119 251234 86128
rect 250628 54732 250680 54738
rect 250628 54674 250680 54680
rect 250536 32496 250588 32502
rect 250536 32438 250588 32444
rect 249800 23452 249852 23458
rect 249800 23394 249852 23400
rect 249800 20664 249852 20670
rect 249800 20606 249852 20612
rect 250812 20664 250864 20670
rect 250812 20606 250864 20612
rect 248420 20596 248472 20602
rect 248420 20538 248472 20544
rect 249156 20596 249208 20602
rect 249156 20538 249208 20544
rect 246304 18692 246356 18698
rect 246304 18634 246356 18640
rect 246316 16574 246344 18634
rect 244292 16546 245240 16574
rect 246316 16546 246436 16574
rect 242898 10976 242954 10985
rect 242898 10911 242954 10920
rect 243542 10976 243598 10985
rect 243542 10911 243598 10920
rect 242912 3534 242940 10911
rect 242992 3596 243044 3602
rect 242992 3538 243044 3544
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 243004 2394 243032 3538
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 242912 2366 243032 2394
rect 242912 480 242940 2366
rect 244108 480 244136 3470
rect 245212 480 245240 16546
rect 246408 4146 246436 16546
rect 246396 4140 246448 4146
rect 246396 4082 246448 4088
rect 246408 480 246436 4082
rect 247592 3596 247644 3602
rect 247592 3538 247644 3544
rect 247604 480 247632 3538
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 20538
rect 249812 16574 249840 20606
rect 250824 20058 250852 20606
rect 250812 20052 250864 20058
rect 250812 19994 250864 20000
rect 249812 16546 250024 16574
rect 249996 480 250024 16546
rect 251192 3670 251220 86119
rect 251836 60042 251864 95202
rect 252480 91050 252508 96591
rect 252468 91044 252520 91050
rect 252468 90986 252520 90992
rect 252480 89758 252508 90986
rect 251916 89752 251968 89758
rect 251916 89694 251968 89700
rect 252468 89752 252520 89758
rect 252468 89694 252520 89700
rect 251928 66230 251956 89694
rect 251916 66224 251968 66230
rect 251916 66166 251968 66172
rect 251824 60036 251876 60042
rect 251824 59978 251876 59984
rect 251272 57248 251324 57254
rect 251272 57190 251324 57196
rect 251180 3664 251232 3670
rect 251180 3606 251232 3612
rect 251284 3482 251312 57190
rect 252560 21616 252612 21622
rect 252560 21558 252612 21564
rect 252572 6914 252600 21558
rect 253216 13190 253244 109006
rect 253308 50522 253336 138042
rect 253400 111790 253428 145522
rect 254584 139460 254636 139466
rect 254584 139402 254636 139408
rect 253388 111784 253440 111790
rect 253388 111726 253440 111732
rect 253388 91792 253440 91798
rect 253388 91734 253440 91740
rect 253296 50516 253348 50522
rect 253296 50458 253348 50464
rect 253400 22098 253428 91734
rect 253388 22092 253440 22098
rect 253388 22034 253440 22040
rect 253400 21622 253428 22034
rect 253388 21616 253440 21622
rect 253388 21558 253440 21564
rect 253204 13184 253256 13190
rect 253204 13126 253256 13132
rect 254596 10334 254624 139402
rect 254688 110430 254716 150418
rect 254860 146532 254912 146538
rect 254860 146474 254912 146480
rect 254768 142180 254820 142186
rect 254768 142122 254820 142128
rect 254676 110424 254728 110430
rect 254676 110366 254728 110372
rect 254780 102882 254808 142122
rect 254872 120154 254900 146474
rect 254860 120148 254912 120154
rect 254860 120090 254912 120096
rect 255976 110362 256004 150486
rect 256148 148368 256200 148374
rect 256148 148310 256200 148316
rect 256056 147688 256108 147694
rect 256056 147630 256108 147636
rect 255964 110356 256016 110362
rect 255964 110298 256016 110304
rect 256068 107574 256096 147630
rect 256160 113082 256188 148310
rect 256252 121446 256280 153818
rect 256712 148986 256740 187274
rect 256884 181756 256936 181762
rect 256884 181698 256936 181704
rect 256792 180328 256844 180334
rect 256792 180270 256844 180276
rect 256804 150278 256832 180270
rect 256896 172446 256924 181698
rect 256884 172440 256936 172446
rect 256884 172382 256936 172388
rect 258092 167958 258120 252622
rect 259460 238196 259512 238202
rect 259460 238138 259512 238144
rect 258172 189916 258224 189922
rect 258172 189858 258224 189864
rect 258080 167952 258132 167958
rect 258080 167894 258132 167900
rect 257344 167068 257396 167074
rect 257344 167010 257396 167016
rect 256792 150272 256844 150278
rect 256792 150214 256844 150220
rect 256700 148980 256752 148986
rect 256700 148922 256752 148928
rect 257356 129606 257384 167010
rect 258184 159390 258212 189858
rect 258356 178968 258408 178974
rect 258356 178910 258408 178916
rect 258264 177404 258316 177410
rect 258264 177346 258316 177352
rect 258276 162246 258304 177346
rect 258368 166394 258396 178910
rect 258356 166388 258408 166394
rect 258356 166330 258408 166336
rect 258724 165640 258776 165646
rect 258724 165582 258776 165588
rect 258264 162240 258316 162246
rect 258264 162182 258316 162188
rect 258172 159384 258224 159390
rect 258172 159326 258224 159332
rect 257436 151836 257488 151842
rect 257436 151778 257488 151784
rect 257344 129600 257396 129606
rect 257344 129542 257396 129548
rect 256240 121440 256292 121446
rect 256240 121382 256292 121388
rect 257344 120216 257396 120222
rect 257344 120158 257396 120164
rect 256148 113076 256200 113082
rect 256148 113018 256200 113024
rect 256056 107568 256108 107574
rect 256056 107510 256108 107516
rect 256148 106344 256200 106350
rect 256148 106286 256200 106292
rect 255964 103556 256016 103562
rect 255964 103498 256016 103504
rect 254768 102876 254820 102882
rect 254768 102818 254820 102824
rect 254676 76560 254728 76566
rect 254676 76502 254728 76508
rect 254688 58002 254716 76502
rect 254676 57996 254728 58002
rect 254676 57938 254728 57944
rect 254584 10328 254636 10334
rect 254584 10270 254636 10276
rect 252572 6886 253520 6914
rect 252376 3664 252428 3670
rect 252376 3606 252428 3612
rect 251192 3454 251312 3482
rect 251192 480 251220 3454
rect 252388 480 252416 3606
rect 253492 480 253520 6886
rect 254688 480 254716 57938
rect 255976 26926 256004 103498
rect 256160 68406 256188 106286
rect 256148 68400 256200 68406
rect 256148 68342 256200 68348
rect 256056 35284 256108 35290
rect 256056 35226 256108 35232
rect 255964 26920 256016 26926
rect 255964 26862 256016 26868
rect 256068 13734 256096 35226
rect 255872 13728 255924 13734
rect 255872 13670 255924 13676
rect 256056 13728 256108 13734
rect 256056 13670 256108 13676
rect 255884 480 255912 13670
rect 257356 11830 257384 120158
rect 257448 111722 257476 151778
rect 257528 146396 257580 146402
rect 257528 146338 257580 146344
rect 257436 111716 257488 111722
rect 257436 111658 257488 111664
rect 257436 109132 257488 109138
rect 257436 109074 257488 109080
rect 257448 18766 257476 109074
rect 257540 104786 257568 146338
rect 258736 128178 258764 165582
rect 259000 160132 259052 160138
rect 259000 160074 259052 160080
rect 258816 157412 258868 157418
rect 258816 157354 258868 157360
rect 258724 128172 258776 128178
rect 258724 128114 258776 128120
rect 258724 120284 258776 120290
rect 258724 120226 258776 120232
rect 257528 104780 257580 104786
rect 257528 104722 257580 104728
rect 257436 18760 257488 18766
rect 257436 18702 257488 18708
rect 258736 14618 258764 120226
rect 258828 117706 258856 157354
rect 258906 140040 258962 140049
rect 259012 140010 259040 160074
rect 259472 158098 259500 238138
rect 259644 200932 259696 200938
rect 259644 200874 259696 200880
rect 259552 198144 259604 198150
rect 259552 198086 259604 198092
rect 259564 166122 259592 198086
rect 259656 170134 259684 200874
rect 259736 180260 259788 180266
rect 259736 180202 259788 180208
rect 259644 170128 259696 170134
rect 259644 170070 259696 170076
rect 259552 166116 259604 166122
rect 259552 166058 259604 166064
rect 259748 159458 259776 180202
rect 260288 164280 260340 164286
rect 260288 164222 260340 164228
rect 259736 159452 259788 159458
rect 259736 159394 259788 159400
rect 260196 158772 260248 158778
rect 260196 158714 260248 158720
rect 259460 158092 259512 158098
rect 259460 158034 259512 158040
rect 258906 139975 258962 139984
rect 259000 140004 259052 140010
rect 258816 117700 258868 117706
rect 258816 117642 258868 117648
rect 258920 102610 258948 139975
rect 259000 139946 259052 139952
rect 260104 136740 260156 136746
rect 260104 136682 260156 136688
rect 259000 133204 259052 133210
rect 259000 133146 259052 133152
rect 259012 106962 259040 133146
rect 259000 106956 259052 106962
rect 259000 106898 259052 106904
rect 258908 102604 258960 102610
rect 258908 102546 258960 102552
rect 258816 102196 258868 102202
rect 258816 102138 258868 102144
rect 258828 62898 258856 102138
rect 260116 65686 260144 136682
rect 260208 119882 260236 158714
rect 260300 137290 260328 164222
rect 260852 144906 260880 256702
rect 263600 244316 263652 244322
rect 263600 244258 263652 244264
rect 263612 242894 263640 244258
rect 263600 242888 263652 242894
rect 263600 242830 263652 242836
rect 263600 207732 263652 207738
rect 263600 207674 263652 207680
rect 262312 199708 262364 199714
rect 262312 199650 262364 199656
rect 260932 195492 260984 195498
rect 260932 195434 260984 195440
rect 260944 162178 260972 195434
rect 261116 183184 261168 183190
rect 261116 183126 261168 183132
rect 261024 177540 261076 177546
rect 261024 177482 261076 177488
rect 260932 162172 260984 162178
rect 260932 162114 260984 162120
rect 261036 158710 261064 177482
rect 261128 171018 261156 183126
rect 262220 175976 262272 175982
rect 262220 175918 262272 175924
rect 262232 171086 262260 175918
rect 262220 171080 262272 171086
rect 262220 171022 262272 171028
rect 261116 171012 261168 171018
rect 261116 170954 261168 170960
rect 262324 168366 262352 199650
rect 262496 177472 262548 177478
rect 262496 177414 262548 177420
rect 262404 176044 262456 176050
rect 262404 175986 262456 175992
rect 262312 168360 262364 168366
rect 262312 168302 262364 168308
rect 261668 162920 261720 162926
rect 261668 162862 261720 162868
rect 261484 161492 261536 161498
rect 261484 161434 261536 161440
rect 261024 158704 261076 158710
rect 261024 158646 261076 158652
rect 260840 144900 260892 144906
rect 260840 144842 260892 144848
rect 260288 137284 260340 137290
rect 260288 137226 260340 137232
rect 261496 122670 261524 161434
rect 261576 155984 261628 155990
rect 261576 155926 261628 155932
rect 261484 122664 261536 122670
rect 261484 122606 261536 122612
rect 260196 119876 260248 119882
rect 260196 119818 260248 119824
rect 261588 117230 261616 155926
rect 261680 124030 261708 162862
rect 262416 157350 262444 175986
rect 262404 157344 262456 157350
rect 262404 157286 262456 157292
rect 262508 142118 262536 177414
rect 262864 169788 262916 169794
rect 262864 169730 262916 169736
rect 262496 142112 262548 142118
rect 262496 142054 262548 142060
rect 262876 130966 262904 169730
rect 263048 160200 263100 160206
rect 263048 160142 263100 160148
rect 262956 140820 263008 140826
rect 262956 140762 263008 140768
rect 262864 130960 262916 130966
rect 262864 130902 262916 130908
rect 261668 124024 261720 124030
rect 261668 123966 261720 123972
rect 261576 117224 261628 117230
rect 261576 117166 261628 117172
rect 262968 105670 262996 140762
rect 263060 124982 263088 160142
rect 263612 139398 263640 207674
rect 264980 206372 265032 206378
rect 264980 206314 265032 206320
rect 263692 203720 263744 203726
rect 263692 203662 263744 203668
rect 263704 165442 263732 203662
rect 263784 184340 263836 184346
rect 263784 184282 263836 184288
rect 263796 169658 263824 184282
rect 264244 172576 264296 172582
rect 264244 172518 264296 172524
rect 263784 169652 263836 169658
rect 263784 169594 263836 169600
rect 263692 165436 263744 165442
rect 263692 165378 263744 165384
rect 263600 139392 263652 139398
rect 263600 139334 263652 139340
rect 264256 133754 264284 172518
rect 264428 164892 264480 164898
rect 264428 164834 264480 164840
rect 264336 154624 264388 154630
rect 264336 154566 264388 154572
rect 264244 133748 264296 133754
rect 264244 133690 264296 133696
rect 264244 128376 264296 128382
rect 264244 128318 264296 128324
rect 263048 124976 263100 124982
rect 263048 124918 263100 124924
rect 262956 105664 263008 105670
rect 262956 105606 263008 105612
rect 261484 104916 261536 104922
rect 261484 104858 261536 104864
rect 260104 65680 260156 65686
rect 259550 65648 259606 65657
rect 260104 65622 260156 65628
rect 259550 65583 259552 65592
rect 259604 65583 259606 65592
rect 259552 65554 259604 65560
rect 258816 62892 258868 62898
rect 258816 62834 258868 62840
rect 260840 60308 260892 60314
rect 260840 60250 260892 60256
rect 259368 58744 259420 58750
rect 259368 58686 259420 58692
rect 259380 58002 259408 58686
rect 259368 57996 259420 58002
rect 259368 57938 259420 57944
rect 259460 22840 259512 22846
rect 259460 22782 259512 22788
rect 258724 14612 258776 14618
rect 258724 14554 258776 14560
rect 257436 13252 257488 13258
rect 257436 13194 257488 13200
rect 257344 11824 257396 11830
rect 257344 11766 257396 11772
rect 257448 5506 257476 13194
rect 258446 10976 258502 10985
rect 258446 10911 258448 10920
rect 258500 10911 258502 10920
rect 259368 10940 259420 10946
rect 258448 10882 258500 10888
rect 259368 10882 259420 10888
rect 259380 10334 259408 10882
rect 259368 10328 259420 10334
rect 259368 10270 259420 10276
rect 257068 5500 257120 5506
rect 257068 5442 257120 5448
rect 257436 5500 257488 5506
rect 257436 5442 257488 5448
rect 257080 480 257108 5442
rect 259380 3505 259408 10270
rect 259472 3602 259500 22782
rect 260852 16574 260880 60250
rect 261496 60110 261524 104858
rect 261576 82136 261628 82142
rect 261576 82078 261628 82084
rect 261588 60722 261616 82078
rect 263506 81560 263562 81569
rect 263506 81495 263562 81504
rect 261576 60716 261628 60722
rect 261576 60658 261628 60664
rect 261588 60314 261616 60658
rect 261576 60308 261628 60314
rect 261576 60250 261628 60256
rect 261484 60104 261536 60110
rect 261484 60046 261536 60052
rect 260852 16546 261800 16574
rect 260746 11792 260802 11801
rect 260746 11727 260802 11736
rect 259460 3596 259512 3602
rect 259460 3538 259512 3544
rect 260656 3596 260708 3602
rect 260656 3538 260708 3544
rect 258262 3496 258318 3505
rect 258262 3431 258318 3440
rect 259366 3496 259422 3505
rect 259366 3431 259422 3440
rect 258276 480 258304 3431
rect 259458 3360 259514 3369
rect 259458 3295 259514 3304
rect 259472 480 259500 3295
rect 260668 480 260696 3538
rect 260760 3369 260788 11727
rect 260746 3360 260802 3369
rect 260746 3295 260802 3304
rect 261772 480 261800 16546
rect 263520 3505 263548 81495
rect 263598 56536 263654 56545
rect 263598 56471 263654 56480
rect 263612 55962 263640 56471
rect 263600 55956 263652 55962
rect 263600 55898 263652 55904
rect 263612 3670 263640 55898
rect 264256 42158 264284 128318
rect 264348 115870 264376 154566
rect 264440 126818 264468 164834
rect 264992 155854 265020 206314
rect 265164 189984 265216 189990
rect 265164 189926 265216 189932
rect 265072 182912 265124 182918
rect 265072 182854 265124 182860
rect 265084 162790 265112 182854
rect 265176 169590 265204 189926
rect 265164 169584 265216 169590
rect 265164 169526 265216 169532
rect 265072 162784 265124 162790
rect 265072 162726 265124 162732
rect 264980 155848 265032 155854
rect 264980 155790 265032 155796
rect 264428 126812 264480 126818
rect 264428 126754 264480 126760
rect 264336 115864 264388 115870
rect 264336 115806 264388 115812
rect 264336 106412 264388 106418
rect 264336 106354 264388 106360
rect 264348 57322 264376 106354
rect 265636 62082 265664 323614
rect 266360 299600 266412 299606
rect 266360 299542 266412 299548
rect 265808 167680 265860 167686
rect 265808 167622 265860 167628
rect 265716 158840 265768 158846
rect 265716 158782 265768 158788
rect 265728 120018 265756 158782
rect 265820 129674 265848 167622
rect 266372 165510 266400 299542
rect 267740 273284 267792 273290
rect 267740 273226 267792 273232
rect 266452 199572 266504 199578
rect 266452 199514 266504 199520
rect 266360 165504 266412 165510
rect 266360 165446 266412 165452
rect 266464 162858 266492 199514
rect 267004 174140 267056 174146
rect 267004 174082 267056 174088
rect 266452 162852 266504 162858
rect 266452 162794 266504 162800
rect 267016 136474 267044 174082
rect 267752 172514 267780 273226
rect 270500 263696 270552 263702
rect 270500 263638 270552 263644
rect 269120 245676 269172 245682
rect 269120 245618 269172 245624
rect 267832 211948 267884 211954
rect 267832 211890 267884 211896
rect 267740 172508 267792 172514
rect 267740 172450 267792 172456
rect 267096 168428 267148 168434
rect 267096 168370 267148 168376
rect 267004 136468 267056 136474
rect 267004 136410 267056 136416
rect 267108 131034 267136 168370
rect 267280 149116 267332 149122
rect 267280 149058 267332 149064
rect 267188 144288 267240 144294
rect 267188 144230 267240 144236
rect 267096 131028 267148 131034
rect 267096 130970 267148 130976
rect 265808 129668 265860 129674
rect 265808 129610 265860 129616
rect 265716 120012 265768 120018
rect 265716 119954 265768 119960
rect 265716 117564 265768 117570
rect 265716 117506 265768 117512
rect 264980 62076 265032 62082
rect 264980 62018 265032 62024
rect 265624 62076 265676 62082
rect 265624 62018 265676 62024
rect 264336 57316 264388 57322
rect 264336 57258 264388 57264
rect 264244 42152 264296 42158
rect 264244 42094 264296 42100
rect 263692 24200 263744 24206
rect 263690 24168 263692 24177
rect 263744 24168 263746 24177
rect 263690 24103 263746 24112
rect 264610 11792 264666 11801
rect 264610 11727 264666 11736
rect 263600 3664 263652 3670
rect 263600 3606 263652 3612
rect 262954 3496 263010 3505
rect 262954 3431 263010 3440
rect 263506 3496 263562 3505
rect 263506 3431 263562 3440
rect 262968 480 262996 3431
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 354 264234 480
rect 264624 354 264652 11727
rect 264122 326 264652 354
rect 264992 354 265020 62018
rect 265728 29714 265756 117506
rect 267004 116000 267056 116006
rect 267004 115942 267056 115948
rect 265716 29708 265768 29714
rect 265716 29650 265768 29656
rect 267016 24138 267044 115942
rect 267200 107642 267228 144230
rect 267292 116618 267320 149058
rect 267844 146198 267872 211890
rect 267924 191276 267976 191282
rect 267924 191218 267976 191224
rect 267936 163538 267964 191218
rect 268016 183116 268068 183122
rect 268016 183058 268068 183064
rect 267924 163532 267976 163538
rect 267924 163474 267976 163480
rect 268028 155242 268056 183058
rect 268568 169856 268620 169862
rect 268568 169798 268620 169804
rect 268384 163532 268436 163538
rect 268384 163474 268436 163480
rect 268016 155236 268068 155242
rect 268016 155178 268068 155184
rect 267832 146192 267884 146198
rect 267832 146134 267884 146140
rect 267372 130416 267424 130422
rect 267372 130358 267424 130364
rect 267280 116612 267332 116618
rect 267280 116554 267332 116560
rect 267188 107636 267240 107642
rect 267188 107578 267240 107584
rect 267384 99278 267412 130358
rect 268396 126886 268424 163474
rect 268476 153264 268528 153270
rect 268476 153206 268528 153212
rect 268384 126880 268436 126886
rect 268384 126822 268436 126828
rect 268488 115258 268516 153206
rect 268580 144362 268608 169798
rect 268568 144356 268620 144362
rect 268568 144298 268620 144304
rect 269132 143478 269160 245618
rect 269212 202224 269264 202230
rect 269212 202166 269264 202172
rect 269224 160070 269252 202166
rect 269304 184476 269356 184482
rect 269304 184418 269356 184424
rect 269316 164082 269344 184418
rect 269764 166320 269816 166326
rect 269764 166262 269816 166268
rect 269304 164076 269356 164082
rect 269304 164018 269356 164024
rect 269212 160064 269264 160070
rect 269212 160006 269264 160012
rect 269120 143472 269172 143478
rect 269120 143414 269172 143420
rect 268568 135924 268620 135930
rect 268568 135866 268620 135872
rect 268476 115252 268528 115258
rect 268476 115194 268528 115200
rect 268384 114572 268436 114578
rect 268384 114514 268436 114520
rect 267372 99272 267424 99278
rect 267372 99214 267424 99220
rect 267096 96688 267148 96694
rect 267096 96630 267148 96636
rect 267108 53106 267136 96630
rect 267646 81424 267702 81433
rect 267646 81359 267702 81368
rect 267096 53100 267148 53106
rect 267096 53042 267148 53048
rect 267004 24132 267056 24138
rect 267004 24074 267056 24080
rect 267660 3505 267688 81359
rect 267740 62892 267792 62898
rect 267740 62834 267792 62840
rect 267752 58041 267780 62834
rect 267738 58032 267794 58041
rect 267738 57967 267794 57976
rect 268396 17270 268424 114514
rect 268476 107908 268528 107914
rect 268476 107850 268528 107856
rect 268488 56030 268516 107850
rect 268580 100570 268608 135866
rect 269776 128246 269804 166262
rect 270512 164150 270540 263638
rect 271880 196784 271932 196790
rect 271880 196726 271932 196732
rect 270684 185836 270736 185842
rect 270684 185778 270736 185784
rect 270592 177336 270644 177342
rect 270592 177278 270644 177284
rect 270500 164144 270552 164150
rect 270500 164086 270552 164092
rect 270604 143546 270632 177278
rect 270696 155922 270724 185778
rect 271144 172644 271196 172650
rect 271144 172586 271196 172592
rect 270684 155916 270736 155922
rect 270684 155858 270736 155864
rect 270592 143540 270644 143546
rect 270592 143482 270644 143488
rect 271156 135182 271184 172586
rect 271236 156052 271288 156058
rect 271236 155994 271288 156000
rect 271144 135176 271196 135182
rect 271144 135118 271196 135124
rect 269764 128240 269816 128246
rect 269764 128182 269816 128188
rect 269856 127016 269908 127022
rect 269856 126958 269908 126964
rect 269764 111852 269816 111858
rect 269764 111794 269816 111800
rect 268568 100564 268620 100570
rect 268568 100506 268620 100512
rect 268476 56024 268528 56030
rect 268476 55966 268528 55972
rect 269118 47560 269174 47569
rect 269118 47495 269120 47504
rect 269172 47495 269174 47504
rect 269120 47466 269172 47472
rect 268384 17264 268436 17270
rect 268384 17206 268436 17212
rect 268382 12336 268438 12345
rect 268382 12271 268438 12280
rect 266542 3496 266598 3505
rect 266542 3431 266598 3440
rect 267646 3496 267702 3505
rect 267646 3431 267702 3440
rect 266556 480 266584 3431
rect 267740 3392 267792 3398
rect 267740 3334 267792 3340
rect 267752 480 267780 3334
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 264122 -960 264234 326
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 12271
rect 269776 4826 269804 111794
rect 269868 47598 269896 126958
rect 271248 117298 271276 155994
rect 271892 146266 271920 196726
rect 271972 190052 272024 190058
rect 271972 189994 272024 190000
rect 271984 161430 272012 189994
rect 271972 161424 272024 161430
rect 271972 161366 272024 161372
rect 271880 146260 271932 146266
rect 271880 146202 271932 146208
rect 271420 139528 271472 139534
rect 271420 139470 271472 139476
rect 271236 117292 271288 117298
rect 271236 117234 271288 117240
rect 271144 116068 271196 116074
rect 271144 116010 271196 116016
rect 269856 47592 269908 47598
rect 269856 47534 269908 47540
rect 270590 27024 270646 27033
rect 270590 26959 270646 26968
rect 270604 26926 270632 26959
rect 270592 26920 270644 26926
rect 270592 26862 270644 26868
rect 270314 11792 270370 11801
rect 270314 11727 270370 11736
rect 269764 4820 269816 4826
rect 269764 4762 269816 4768
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 354 270122 480
rect 270328 354 270356 11727
rect 271156 7614 271184 116010
rect 271328 103624 271380 103630
rect 271328 103566 271380 103572
rect 271236 100972 271288 100978
rect 271236 100914 271288 100920
rect 271248 46238 271276 100914
rect 271340 61402 271368 103566
rect 271432 101454 271460 139470
rect 271512 119400 271564 119406
rect 271512 119342 271564 119348
rect 271524 104854 271552 119342
rect 271512 104848 271564 104854
rect 271512 104790 271564 104796
rect 271420 101448 271472 101454
rect 271420 101390 271472 101396
rect 272536 64870 272564 368999
rect 273904 311228 273956 311234
rect 273904 311170 273956 311176
rect 273260 210520 273312 210526
rect 273260 210462 273312 210468
rect 273272 164218 273300 210462
rect 273352 195356 273404 195362
rect 273352 195298 273404 195304
rect 273260 164212 273312 164218
rect 273260 164154 273312 164160
rect 272708 161560 272760 161566
rect 272708 161502 272760 161508
rect 272720 122738 272748 161502
rect 273364 154562 273392 195298
rect 273352 154556 273404 154562
rect 273352 154498 273404 154504
rect 272708 122732 272760 122738
rect 272708 122674 272760 122680
rect 272616 121508 272668 121514
rect 272616 121450 272668 121456
rect 272524 64864 272576 64870
rect 272524 64806 272576 64812
rect 272536 63578 272564 64806
rect 271880 63572 271932 63578
rect 271880 63514 271932 63520
rect 272524 63572 272576 63578
rect 272524 63514 272576 63520
rect 271328 61396 271380 61402
rect 271328 61338 271380 61344
rect 271236 46232 271288 46238
rect 271236 46174 271288 46180
rect 271236 17264 271288 17270
rect 271236 17206 271288 17212
rect 271144 7608 271196 7614
rect 271144 7550 271196 7556
rect 271248 3602 271276 17206
rect 271892 16574 271920 63514
rect 272628 38010 272656 121450
rect 273258 41304 273314 41313
rect 273258 41239 273314 41248
rect 272616 38004 272668 38010
rect 272616 37946 272668 37952
rect 271892 16546 272472 16574
rect 271786 12744 271842 12753
rect 271786 12679 271842 12688
rect 271236 3596 271288 3602
rect 271236 3538 271288 3544
rect 271800 3505 271828 12679
rect 271234 3496 271290 3505
rect 271234 3431 271290 3440
rect 271786 3496 271842 3505
rect 271786 3431 271842 3440
rect 271248 480 271276 3431
rect 272444 480 272472 16546
rect 270010 326 270356 354
rect 270010 -960 270122 326
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 354 273300 41239
rect 273916 3942 273944 311170
rect 275284 305720 275336 305726
rect 275284 305662 275336 305668
rect 274640 188556 274692 188562
rect 274640 188498 274692 188504
rect 273996 171148 274048 171154
rect 273996 171090 274048 171096
rect 274008 132394 274036 171090
rect 274088 155236 274140 155242
rect 274088 155178 274140 155184
rect 273996 132388 274048 132394
rect 273996 132330 274048 132336
rect 273996 129804 274048 129810
rect 273996 129746 274048 129752
rect 274008 40798 274036 129746
rect 274100 118590 274128 155178
rect 274652 147558 274680 188498
rect 274732 187264 274784 187270
rect 274732 187206 274784 187212
rect 274744 153134 274772 187206
rect 274732 153128 274784 153134
rect 274732 153070 274784 153076
rect 274640 147552 274692 147558
rect 274640 147494 274692 147500
rect 274180 142860 274232 142866
rect 274180 142802 274232 142808
rect 274088 118584 274140 118590
rect 274088 118526 274140 118532
rect 274192 103494 274220 142802
rect 274180 103488 274232 103494
rect 274180 103430 274232 103436
rect 274088 102264 274140 102270
rect 274088 102206 274140 102212
rect 273996 40792 274048 40798
rect 273996 40734 274048 40740
rect 274100 31142 274128 102206
rect 274178 71088 274234 71097
rect 274178 71023 274234 71032
rect 274192 41313 274220 71023
rect 274178 41304 274234 41313
rect 274178 41239 274234 41248
rect 274088 31136 274140 31142
rect 274088 31078 274140 31084
rect 274640 25696 274692 25702
rect 274640 25638 274692 25644
rect 273904 3936 273956 3942
rect 273904 3878 273956 3884
rect 274652 3398 274680 25638
rect 275296 4010 275324 305662
rect 276020 298172 276072 298178
rect 276020 298114 276072 298120
rect 275560 149184 275612 149190
rect 275560 149126 275612 149132
rect 275376 133952 275428 133958
rect 275376 133894 275428 133900
rect 275388 28286 275416 133894
rect 275572 108934 275600 149126
rect 276032 140690 276060 298114
rect 276112 222896 276164 222902
rect 276112 222838 276164 222844
rect 276124 165578 276152 222838
rect 276204 191344 276256 191350
rect 276204 191286 276256 191292
rect 276112 165572 276164 165578
rect 276112 165514 276164 165520
rect 276216 153066 276244 191286
rect 276204 153060 276256 153066
rect 276204 153002 276256 153008
rect 276020 140684 276072 140690
rect 276020 140626 276072 140632
rect 275560 108928 275612 108934
rect 275560 108870 275612 108876
rect 275468 107772 275520 107778
rect 275468 107714 275520 107720
rect 275480 54670 275508 107714
rect 276020 87644 276072 87650
rect 276020 87586 276072 87592
rect 276032 87038 276060 87586
rect 276020 87032 276072 87038
rect 276020 86974 276072 86980
rect 275468 54664 275520 54670
rect 275468 54606 275520 54612
rect 276676 42702 276704 378762
rect 283562 367704 283618 367713
rect 283562 367639 283618 367648
rect 280804 355360 280856 355366
rect 280804 355302 280856 355308
rect 278044 342916 278096 342922
rect 278044 342858 278096 342864
rect 277400 235408 277452 235414
rect 277400 235350 277452 235356
rect 276756 157480 276808 157486
rect 276756 157422 276808 157428
rect 276768 149705 276796 157422
rect 276754 149696 276810 149705
rect 276754 149631 276810 149640
rect 276848 146464 276900 146470
rect 276848 146406 276900 146412
rect 276756 128444 276808 128450
rect 276756 128386 276808 128392
rect 276020 42696 276072 42702
rect 276020 42638 276072 42644
rect 276664 42696 276716 42702
rect 276664 42638 276716 42644
rect 275376 28280 275428 28286
rect 275376 28222 275428 28228
rect 276032 16574 276060 42638
rect 276768 25634 276796 128386
rect 276860 112470 276888 146406
rect 277412 137970 277440 235350
rect 277492 192704 277544 192710
rect 277492 192646 277544 192652
rect 277504 140758 277532 192646
rect 277492 140752 277544 140758
rect 277492 140694 277544 140700
rect 277400 137964 277452 137970
rect 277400 137906 277452 137912
rect 276940 125656 276992 125662
rect 276940 125598 276992 125604
rect 276848 112464 276900 112470
rect 276848 112406 276900 112412
rect 276848 87032 276900 87038
rect 276848 86974 276900 86980
rect 276756 25628 276808 25634
rect 276756 25570 276808 25576
rect 276032 16546 276704 16574
rect 274824 4004 274876 4010
rect 274824 3946 274876 3952
rect 275284 4004 275336 4010
rect 275284 3946 275336 3952
rect 274640 3392 274692 3398
rect 274640 3334 274692 3340
rect 274836 480 274864 3946
rect 276020 3528 276072 3534
rect 276020 3470 276072 3476
rect 276032 480 276060 3470
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 16546
rect 276860 3534 276888 86974
rect 276952 68474 276980 125598
rect 277400 91792 277452 91798
rect 277400 91734 277452 91740
rect 277412 87038 277440 91734
rect 278056 87650 278084 342858
rect 279424 307080 279476 307086
rect 279424 307022 279476 307028
rect 278780 235340 278832 235346
rect 278780 235282 278832 235288
rect 278228 168496 278280 168502
rect 278228 168438 278280 168444
rect 278136 131164 278188 131170
rect 278136 131106 278188 131112
rect 278044 87644 278096 87650
rect 278044 87586 278096 87592
rect 277400 87032 277452 87038
rect 277400 86974 277452 86980
rect 278044 80708 278096 80714
rect 278044 80650 278096 80656
rect 276940 68468 276992 68474
rect 276940 68410 276992 68416
rect 278056 30326 278084 80650
rect 277400 30320 277452 30326
rect 277400 30262 277452 30268
rect 278044 30320 278096 30326
rect 278044 30262 278096 30268
rect 277412 16574 277440 30262
rect 278148 19990 278176 131106
rect 278240 129742 278268 168438
rect 278792 147626 278820 235282
rect 278780 147620 278832 147626
rect 278780 147562 278832 147568
rect 278318 137320 278374 137329
rect 278318 137255 278374 137264
rect 278228 129736 278280 129742
rect 278228 129678 278280 129684
rect 278228 124228 278280 124234
rect 278228 124170 278280 124176
rect 278240 93158 278268 124170
rect 278332 109002 278360 137255
rect 278320 108996 278372 109002
rect 278320 108938 278372 108944
rect 278320 96756 278372 96762
rect 278320 96698 278372 96704
rect 278228 93152 278280 93158
rect 278228 93094 278280 93100
rect 278332 39370 278360 96698
rect 279436 66230 279464 307022
rect 280160 192772 280212 192778
rect 280160 192714 280212 192720
rect 280172 150346 280200 192714
rect 280160 150340 280212 150346
rect 280160 150282 280212 150288
rect 279608 118856 279660 118862
rect 279608 118798 279660 118804
rect 279516 110492 279568 110498
rect 279516 110434 279568 110440
rect 279424 66224 279476 66230
rect 279424 66166 279476 66172
rect 279436 65482 279464 66166
rect 278780 65476 278832 65482
rect 278780 65418 278832 65424
rect 279424 65476 279476 65482
rect 279424 65418 279476 65424
rect 278320 39364 278372 39370
rect 278320 39306 278372 39312
rect 278136 19984 278188 19990
rect 278136 19926 278188 19932
rect 278792 16574 278820 65418
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 276848 3528 276900 3534
rect 276848 3470 276900 3476
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 279528 15978 279556 110434
rect 279620 65550 279648 118798
rect 279608 65544 279660 65550
rect 279608 65486 279660 65492
rect 280160 44192 280212 44198
rect 280160 44134 280212 44140
rect 280172 16574 280200 44134
rect 280816 40050 280844 355302
rect 280894 330440 280950 330449
rect 280894 330375 280950 330384
rect 280908 45558 280936 330375
rect 282184 329112 282236 329118
rect 282184 329054 282236 329060
rect 281540 220108 281592 220114
rect 281540 220050 281592 220056
rect 281080 149728 281132 149734
rect 281080 149670 281132 149676
rect 280988 114640 281040 114646
rect 280988 114582 281040 114588
rect 280896 45552 280948 45558
rect 280896 45494 280948 45500
rect 280908 44198 280936 45494
rect 280896 44192 280948 44198
rect 280896 44134 280948 44140
rect 280804 40044 280856 40050
rect 280804 39986 280856 39992
rect 280804 28280 280856 28286
rect 280804 28222 280856 28228
rect 280172 16546 280752 16574
rect 279516 15972 279568 15978
rect 279516 15914 279568 15920
rect 280724 480 280752 16546
rect 280816 4010 280844 28222
rect 281000 21418 281028 114582
rect 281092 111654 281120 149670
rect 281552 149054 281580 220050
rect 281540 149048 281592 149054
rect 281540 148990 281592 148996
rect 281080 111648 281132 111654
rect 281080 111590 281132 111596
rect 281080 98116 281132 98122
rect 281080 98058 281132 98064
rect 281092 64190 281120 98058
rect 281080 64184 281132 64190
rect 281080 64126 281132 64132
rect 282196 31142 282224 329054
rect 282276 313948 282328 313954
rect 282276 313890 282328 313896
rect 282184 31136 282236 31142
rect 282184 31078 282236 31084
rect 280988 21412 281040 21418
rect 280988 21354 281040 21360
rect 280804 4004 280856 4010
rect 280804 3946 280856 3952
rect 282196 3330 282224 31078
rect 282288 6866 282316 313890
rect 282460 134020 282512 134026
rect 282460 133962 282512 133968
rect 282368 104984 282420 104990
rect 282368 104926 282420 104932
rect 282380 9042 282408 104926
rect 282472 58818 282500 133962
rect 282460 58812 282512 58818
rect 282460 58754 282512 58760
rect 283576 12442 283604 367639
rect 284944 327752 284996 327758
rect 284944 327694 284996 327700
rect 284300 253972 284352 253978
rect 284300 253914 284352 253920
rect 283748 160744 283800 160750
rect 283748 160686 283800 160692
rect 283760 126954 283788 160686
rect 284312 150414 284340 253914
rect 284300 150408 284352 150414
rect 284300 150350 284352 150356
rect 283748 126948 283800 126954
rect 283748 126890 283800 126896
rect 283656 125724 283708 125730
rect 283656 125666 283708 125672
rect 283104 12436 283156 12442
rect 283104 12378 283156 12384
rect 283564 12436 283616 12442
rect 283564 12378 283616 12384
rect 282368 9036 282420 9042
rect 282368 8978 282420 8984
rect 282276 6860 282328 6866
rect 282276 6802 282328 6808
rect 282184 3324 282236 3330
rect 282184 3266 282236 3272
rect 282288 3210 282316 6802
rect 281920 3182 282316 3210
rect 281920 480 281948 3182
rect 283116 480 283144 12378
rect 283668 6186 283696 125666
rect 283748 117428 283800 117434
rect 283748 117370 283800 117376
rect 283760 32434 283788 117370
rect 284390 49056 284446 49065
rect 284390 48991 284392 49000
rect 284444 48991 284446 49000
rect 284392 48962 284444 48968
rect 284956 46306 284984 327694
rect 285036 172712 285088 172718
rect 285036 172654 285088 172660
rect 285048 135250 285076 172654
rect 285220 156120 285272 156126
rect 285220 156062 285272 156068
rect 285036 135244 285088 135250
rect 285036 135186 285088 135192
rect 285128 132524 285180 132530
rect 285128 132466 285180 132472
rect 285036 127084 285088 127090
rect 285036 127026 285088 127032
rect 284944 46300 284996 46306
rect 284944 46242 284996 46248
rect 283748 32428 283800 32434
rect 283748 32370 283800 32376
rect 284956 9654 284984 46242
rect 285048 44878 285076 127026
rect 285140 62830 285168 132466
rect 285232 115938 285260 156062
rect 285220 115932 285272 115938
rect 285220 115874 285272 115880
rect 285220 99408 285272 99414
rect 285220 99350 285272 99356
rect 285128 62824 285180 62830
rect 285128 62766 285180 62772
rect 285232 48958 285260 99350
rect 286336 67561 286364 386378
rect 287704 385144 287756 385150
rect 287704 385086 287756 385092
rect 286416 171216 286468 171222
rect 286416 171158 286468 171164
rect 286428 133822 286456 171158
rect 286600 154692 286652 154698
rect 286600 154634 286652 154640
rect 286416 133816 286468 133822
rect 286416 133758 286468 133764
rect 286508 132592 286560 132598
rect 286508 132534 286560 132540
rect 286416 124296 286468 124302
rect 286416 124238 286468 124244
rect 286322 67552 286378 67561
rect 286322 67487 286378 67496
rect 285220 48952 285272 48958
rect 285220 48894 285272 48900
rect 285036 44872 285088 44878
rect 285036 44814 285088 44820
rect 286428 24274 286456 124238
rect 286520 61470 286548 132534
rect 286612 114510 286640 154634
rect 286600 114504 286652 114510
rect 286600 114446 286652 114452
rect 286600 103692 286652 103698
rect 286600 103634 286652 103640
rect 286508 61464 286560 61470
rect 286508 61406 286560 61412
rect 286612 43450 286640 103634
rect 286966 67552 287022 67561
rect 286966 67487 287022 67496
rect 286600 43444 286652 43450
rect 286600 43386 286652 43392
rect 286416 24268 286468 24274
rect 286416 24210 286468 24216
rect 286416 15972 286468 15978
rect 286416 15914 286468 15920
rect 285586 11792 285642 11801
rect 285586 11727 285642 11736
rect 284944 9648 284996 9654
rect 284944 9590 284996 9596
rect 283656 6180 283708 6186
rect 283656 6122 283708 6128
rect 285600 3505 285628 11727
rect 284298 3496 284354 3505
rect 284298 3431 284354 3440
rect 285586 3496 285642 3505
rect 286428 3466 286456 15914
rect 285586 3431 285642 3440
rect 286416 3460 286468 3466
rect 284312 480 284340 3431
rect 286416 3402 286468 3408
rect 285404 3324 285456 3330
rect 285404 3266 285456 3272
rect 285416 480 285444 3266
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 354 286682 480
rect 286980 354 287008 67487
rect 287716 3874 287744 385086
rect 289096 177342 289124 402970
rect 358820 401668 358872 401674
rect 358820 401610 358872 401616
rect 357440 400240 357492 400246
rect 357440 400182 357492 400188
rect 308404 385076 308456 385082
rect 308404 385018 308456 385024
rect 295984 380180 296036 380186
rect 295984 380122 296036 380128
rect 293222 336016 293278 336025
rect 293222 335951 293278 335960
rect 291844 334620 291896 334626
rect 291844 334562 291896 334568
rect 289174 177440 289230 177449
rect 289174 177375 289230 177384
rect 289084 177336 289136 177342
rect 289084 177278 289136 177284
rect 287888 167136 287940 167142
rect 287888 167078 287940 167084
rect 287900 128314 287928 167078
rect 287980 141500 288032 141506
rect 287980 141442 288032 141448
rect 287888 128308 287940 128314
rect 287888 128250 287940 128256
rect 287796 127152 287848 127158
rect 287796 127094 287848 127100
rect 287808 15910 287836 127094
rect 287992 102066 288020 141442
rect 289084 131232 289136 131238
rect 289084 131174 289136 131180
rect 287980 102060 288032 102066
rect 287980 102002 288032 102008
rect 287888 100836 287940 100842
rect 287888 100778 287940 100784
rect 287900 35222 287928 100778
rect 287888 35216 287940 35222
rect 287888 35158 287940 35164
rect 288440 34468 288492 34474
rect 288440 34410 288492 34416
rect 288452 16574 288480 34410
rect 289096 33794 289124 131174
rect 289188 82142 289216 177375
rect 289268 169924 289320 169930
rect 289268 169866 289320 169872
rect 289280 132462 289308 169866
rect 290556 169040 290608 169046
rect 290556 168982 290608 168988
rect 289360 142248 289412 142254
rect 289360 142190 289412 142196
rect 289268 132456 289320 132462
rect 289268 132398 289320 132404
rect 289268 102332 289320 102338
rect 289268 102274 289320 102280
rect 289176 82136 289228 82142
rect 289176 82078 289228 82084
rect 289084 33788 289136 33794
rect 289084 33730 289136 33736
rect 289280 25566 289308 102274
rect 289372 100638 289400 142190
rect 290568 131102 290596 168982
rect 290648 143608 290700 143614
rect 290648 143550 290700 143556
rect 290556 131096 290608 131102
rect 290556 131038 290608 131044
rect 290464 129872 290516 129878
rect 290464 129814 290516 129820
rect 289360 100632 289412 100638
rect 289360 100574 289412 100580
rect 289820 67584 289872 67590
rect 289820 67526 289872 67532
rect 289728 35216 289780 35222
rect 289728 35158 289780 35164
rect 289740 34474 289768 35158
rect 289728 34468 289780 34474
rect 289728 34410 289780 34416
rect 289268 25560 289320 25566
rect 289268 25502 289320 25508
rect 288452 16546 289032 16574
rect 287796 15904 287848 15910
rect 287796 15846 287848 15852
rect 287796 9648 287848 9654
rect 287796 9590 287848 9596
rect 287704 3868 287756 3874
rect 287704 3810 287756 3816
rect 287808 480 287836 9590
rect 289004 480 289032 16546
rect 286570 326 287008 354
rect 286570 -960 286682 326
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 354 289860 67526
rect 290476 22778 290504 129814
rect 290556 113212 290608 113218
rect 290556 113154 290608 113160
rect 290568 66910 290596 113154
rect 290660 102134 290688 143550
rect 290648 102128 290700 102134
rect 290648 102070 290700 102076
rect 291108 68400 291160 68406
rect 291108 68342 291160 68348
rect 291120 67590 291148 68342
rect 291108 67584 291160 67590
rect 291108 67526 291160 67532
rect 290556 66904 290608 66910
rect 290556 66846 290608 66852
rect 291856 33046 291884 334562
rect 292028 158908 292080 158914
rect 292028 158850 292080 158856
rect 291936 129940 291988 129946
rect 291936 129882 291988 129888
rect 291844 33040 291896 33046
rect 291844 32982 291896 32988
rect 291856 31822 291884 32982
rect 291200 31816 291252 31822
rect 291200 31758 291252 31764
rect 291844 31816 291896 31822
rect 291844 31758 291896 31764
rect 290464 22772 290516 22778
rect 290464 22714 290516 22720
rect 291212 16574 291240 31758
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 291948 4894 291976 129882
rect 292040 120086 292068 158850
rect 292120 144968 292172 144974
rect 292120 144910 292172 144916
rect 292028 120080 292080 120086
rect 292028 120022 292080 120028
rect 292028 110560 292080 110566
rect 292028 110502 292080 110508
rect 292040 51746 292068 110502
rect 292132 105602 292160 144910
rect 292120 105596 292172 105602
rect 292120 105538 292172 105544
rect 293236 69766 293264 335951
rect 294604 305652 294656 305658
rect 294604 305594 294656 305600
rect 293408 150612 293460 150618
rect 293408 150554 293460 150560
rect 293316 116136 293368 116142
rect 293316 116078 293368 116084
rect 293224 69760 293276 69766
rect 293224 69702 293276 69708
rect 292028 51740 292080 51746
rect 292028 51682 292080 51688
rect 292580 36644 292632 36650
rect 292580 36586 292632 36592
rect 291936 4888 291988 4894
rect 291936 4830 291988 4836
rect 292592 480 292620 36586
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 69702
rect 293328 36582 293356 116078
rect 293420 111081 293448 150554
rect 293406 111072 293462 111081
rect 293406 111007 293462 111016
rect 293316 36576 293368 36582
rect 293316 36518 293368 36524
rect 293960 4820 294012 4826
rect 293960 4762 294012 4768
rect 293972 3942 294000 4762
rect 294616 4078 294644 305594
rect 294696 164348 294748 164354
rect 294696 164290 294748 164296
rect 294708 141438 294736 164290
rect 294696 141432 294748 141438
rect 294696 141374 294748 141380
rect 294880 138168 294932 138174
rect 294880 138110 294932 138116
rect 294696 131300 294748 131306
rect 294696 131242 294748 131248
rect 294604 4072 294656 4078
rect 294604 4014 294656 4020
rect 293960 3936 294012 3942
rect 293960 3878 294012 3884
rect 294708 2106 294736 131242
rect 294788 110628 294840 110634
rect 294788 110570 294840 110576
rect 294800 2174 294828 110570
rect 294892 53242 294920 138110
rect 295996 89010 296024 380122
rect 301502 370560 301558 370569
rect 301502 370495 301558 370504
rect 297364 347812 297416 347818
rect 297364 347754 297416 347760
rect 296076 161628 296128 161634
rect 296076 161570 296128 161576
rect 296088 122806 296116 161570
rect 296076 122800 296128 122806
rect 296076 122742 296128 122748
rect 296260 121576 296312 121582
rect 296260 121518 296312 121524
rect 296076 114708 296128 114714
rect 296076 114650 296128 114656
rect 295984 89004 296036 89010
rect 295984 88946 296036 88952
rect 294880 53236 294932 53242
rect 294880 53178 294932 53184
rect 295340 38072 295392 38078
rect 295340 38014 295392 38020
rect 295352 16574 295380 38014
rect 295352 16546 295656 16574
rect 294880 4820 294932 4826
rect 294880 4762 294932 4768
rect 294788 2168 294840 2174
rect 294788 2110 294840 2116
rect 294696 2100 294748 2106
rect 294696 2042 294748 2048
rect 294892 480 294920 4762
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 296088 8974 296116 114650
rect 296168 99476 296220 99482
rect 296168 99418 296220 99424
rect 296180 37942 296208 99418
rect 296272 69698 296300 121518
rect 297376 77246 297404 347754
rect 300124 264988 300176 264994
rect 300124 264930 300176 264936
rect 297456 174004 297508 174010
rect 297456 173946 297508 173952
rect 297468 136542 297496 173946
rect 298928 162988 298980 162994
rect 298928 162930 298980 162936
rect 297456 136536 297508 136542
rect 297456 136478 297508 136484
rect 298836 135380 298888 135386
rect 298836 135322 298888 135328
rect 297456 134564 297508 134570
rect 297456 134506 297508 134512
rect 297468 125594 297496 134506
rect 297456 125588 297508 125594
rect 297456 125530 297508 125536
rect 297548 124364 297600 124370
rect 297548 124306 297600 124312
rect 297456 111920 297508 111926
rect 297456 111862 297508 111868
rect 297364 77240 297416 77246
rect 297364 77182 297416 77188
rect 297364 71188 297416 71194
rect 297364 71130 297416 71136
rect 296260 69692 296312 69698
rect 296260 69634 296312 69640
rect 297376 40050 297404 71130
rect 297468 44946 297496 111862
rect 297560 71126 297588 124306
rect 298744 122936 298796 122942
rect 298744 122878 298796 122884
rect 297640 122868 297692 122874
rect 297640 122810 297692 122816
rect 297652 73846 297680 122810
rect 297640 73840 297692 73846
rect 297640 73782 297692 73788
rect 297548 71120 297600 71126
rect 297548 71062 297600 71068
rect 297456 44940 297508 44946
rect 297456 44882 297508 44888
rect 298192 43444 298244 43450
rect 298192 43386 298244 43392
rect 298204 43353 298232 43386
rect 298190 43344 298246 43353
rect 298190 43279 298246 43288
rect 296720 40044 296772 40050
rect 296720 39986 296772 39992
rect 297364 40044 297416 40050
rect 297364 39986 297416 39992
rect 296168 37936 296220 37942
rect 296168 37878 296220 37884
rect 296732 16574 296760 39986
rect 296732 16546 297312 16574
rect 296076 8968 296128 8974
rect 296076 8910 296128 8916
rect 297284 480 297312 16546
rect 298756 11762 298784 122878
rect 298848 43518 298876 135322
rect 298940 124098 298968 162930
rect 299112 152584 299164 152590
rect 299112 152526 299164 152532
rect 298928 124092 298980 124098
rect 298928 124034 298980 124040
rect 299020 118788 299072 118794
rect 299020 118730 299072 118736
rect 298928 111988 298980 111994
rect 298928 111930 298980 111936
rect 298940 47666 298968 111930
rect 299032 75206 299060 118730
rect 299124 113150 299152 152526
rect 299112 113144 299164 113150
rect 299112 113086 299164 113092
rect 300136 96558 300164 264930
rect 300216 157548 300268 157554
rect 300216 157490 300268 157496
rect 300228 118658 300256 157490
rect 300400 121644 300452 121650
rect 300400 121586 300452 121592
rect 300216 118652 300268 118658
rect 300216 118594 300268 118600
rect 300308 107704 300360 107710
rect 300308 107646 300360 107652
rect 300216 100904 300268 100910
rect 300216 100846 300268 100852
rect 300124 96552 300176 96558
rect 300124 96494 300176 96500
rect 299020 75200 299072 75206
rect 299020 75142 299072 75148
rect 300124 75200 300176 75206
rect 300124 75142 300176 75148
rect 298928 47660 298980 47666
rect 298928 47602 298980 47608
rect 298836 43512 298888 43518
rect 298836 43454 298888 43460
rect 299662 39400 299718 39409
rect 299662 39335 299664 39344
rect 299716 39335 299718 39344
rect 299664 39306 299716 39312
rect 299386 11792 299442 11801
rect 298744 11756 298796 11762
rect 299386 11727 299442 11736
rect 298744 11698 298796 11704
rect 299400 3505 299428 11727
rect 300136 9625 300164 75142
rect 300228 40730 300256 100846
rect 300320 50454 300348 107646
rect 300412 75274 300440 121586
rect 300400 75268 300452 75274
rect 300400 75210 300452 75216
rect 300308 50448 300360 50454
rect 300308 50390 300360 50396
rect 300216 40724 300268 40730
rect 300216 40666 300268 40672
rect 301516 16590 301544 370495
rect 305644 365016 305696 365022
rect 305644 364958 305696 364964
rect 304264 309188 304316 309194
rect 304264 309130 304316 309136
rect 304276 184249 304304 309130
rect 304356 213308 304408 213314
rect 304356 213250 304408 213256
rect 304262 184240 304318 184249
rect 304262 184175 304318 184184
rect 304368 175817 304396 213250
rect 304354 175808 304410 175817
rect 304354 175743 304410 175752
rect 302884 174072 302936 174078
rect 302884 174014 302936 174020
rect 301596 153332 301648 153338
rect 301596 153274 301648 153280
rect 301608 113830 301636 153274
rect 301872 140956 301924 140962
rect 301872 140898 301924 140904
rect 301596 113824 301648 113830
rect 301596 113766 301648 113772
rect 301688 113280 301740 113286
rect 301688 113222 301740 113228
rect 301596 106480 301648 106486
rect 301596 106422 301648 106428
rect 301504 16584 301556 16590
rect 301504 16526 301556 16532
rect 300766 11792 300822 11801
rect 300766 11727 300822 11736
rect 300122 9616 300178 9625
rect 300122 9551 300178 9560
rect 300674 9616 300730 9625
rect 300674 9551 300730 9560
rect 299662 3632 299718 3641
rect 299662 3567 299718 3576
rect 298466 3496 298522 3505
rect 298466 3431 298522 3440
rect 299386 3496 299442 3505
rect 299386 3431 299442 3440
rect 298480 480 298508 3431
rect 299676 480 299704 3567
rect 300688 3482 300716 9551
rect 300780 3641 300808 11727
rect 300766 3632 300822 3641
rect 300766 3567 300822 3576
rect 300688 3454 300808 3482
rect 300780 480 300808 3454
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 354 301544 16526
rect 301608 6254 301636 106422
rect 301700 18630 301728 113222
rect 301884 100706 301912 140898
rect 302896 136610 302924 174014
rect 304448 171284 304500 171290
rect 304448 171226 304500 171232
rect 304356 163056 304408 163062
rect 304356 162998 304408 163004
rect 303620 146328 303672 146334
rect 303620 146270 303672 146276
rect 303632 144226 303660 146270
rect 303620 144220 303672 144226
rect 303620 144162 303672 144168
rect 302976 143676 303028 143682
rect 302976 143618 303028 143624
rect 302884 136604 302936 136610
rect 302884 136546 302936 136552
rect 302988 124914 303016 143618
rect 303252 140888 303304 140894
rect 303252 140830 303304 140836
rect 302976 124908 303028 124914
rect 302976 124850 303028 124856
rect 303068 124432 303120 124438
rect 303068 124374 303120 124380
rect 302884 109200 302936 109206
rect 302884 109142 302936 109148
rect 301872 100700 301924 100706
rect 301872 100642 301924 100648
rect 301780 99544 301832 99550
rect 301780 99486 301832 99492
rect 301792 42090 301820 99486
rect 301780 42084 301832 42090
rect 301780 42026 301832 42032
rect 302238 40760 302294 40769
rect 302238 40695 302240 40704
rect 302292 40695 302294 40704
rect 302240 40666 302292 40672
rect 301688 18624 301740 18630
rect 301688 18566 301740 18572
rect 302896 17338 302924 109142
rect 302976 98184 303028 98190
rect 302976 98126 303028 98132
rect 302988 31074 303016 98126
rect 303080 60178 303108 124374
rect 303160 105052 303212 105058
rect 303160 104994 303212 105000
rect 303068 60172 303120 60178
rect 303068 60114 303120 60120
rect 303172 58682 303200 104994
rect 303264 99346 303292 140830
rect 304264 135448 304316 135454
rect 304264 135390 304316 135396
rect 303252 99340 303304 99346
rect 303252 99282 303304 99288
rect 303620 79348 303672 79354
rect 303620 79290 303672 79296
rect 303160 58676 303212 58682
rect 303160 58618 303212 58624
rect 302976 31068 303028 31074
rect 302976 31010 303028 31016
rect 302884 17332 302936 17338
rect 302884 17274 302936 17280
rect 303632 16574 303660 79290
rect 304276 49094 304304 135390
rect 304368 124166 304396 162998
rect 304460 133890 304488 171226
rect 304448 133884 304500 133890
rect 304448 133826 304500 133832
rect 304356 124160 304408 124166
rect 304356 124102 304408 124108
rect 304356 117360 304408 117366
rect 304356 117302 304408 117308
rect 304264 49088 304316 49094
rect 304264 49030 304316 49036
rect 304368 39438 304396 117302
rect 304448 100768 304500 100774
rect 304448 100710 304500 100716
rect 304460 72486 304488 100710
rect 304448 72480 304500 72486
rect 304448 72422 304500 72428
rect 304356 39432 304408 39438
rect 304356 39374 304408 39380
rect 303632 16546 303936 16574
rect 303526 11792 303582 11801
rect 303526 11727 303582 11736
rect 301596 6248 301648 6254
rect 301596 6190 301648 6196
rect 301934 354 302046 480
rect 301516 326 302046 354
rect 301934 -960 302046 326
rect 303130 354 303242 480
rect 303540 354 303568 11727
rect 303130 326 303568 354
rect 303908 354 303936 16546
rect 305656 9654 305684 364958
rect 307024 363656 307076 363662
rect 307024 363598 307076 363604
rect 305736 344344 305788 344350
rect 305736 344286 305788 344292
rect 305748 180334 305776 344286
rect 305736 180328 305788 180334
rect 305736 180270 305788 180276
rect 305734 174040 305790 174049
rect 305734 173975 305790 173984
rect 305748 130422 305776 173975
rect 306562 172272 306618 172281
rect 306562 172207 306618 172216
rect 306576 171222 306604 172207
rect 306564 171216 306616 171222
rect 306564 171158 306616 171164
rect 307036 170134 307064 363598
rect 307390 175264 307446 175273
rect 307390 175199 307446 175208
rect 307404 174049 307432 175199
rect 307482 174856 307538 174865
rect 307482 174791 307538 174800
rect 307390 174040 307446 174049
rect 307496 174010 307524 174791
rect 307666 174448 307722 174457
rect 307666 174383 307722 174392
rect 307680 174146 307708 174383
rect 307668 174140 307720 174146
rect 307668 174082 307720 174088
rect 307576 174072 307628 174078
rect 307574 174040 307576 174049
rect 307628 174040 307630 174049
rect 307390 173975 307446 173984
rect 307484 174004 307536 174010
rect 307574 173975 307630 173984
rect 307484 173946 307536 173952
rect 307574 173632 307630 173641
rect 307574 173567 307630 173576
rect 307482 173224 307538 173233
rect 307482 173159 307538 173168
rect 307496 172650 307524 173159
rect 307588 172718 307616 173567
rect 307576 172712 307628 172718
rect 307576 172654 307628 172660
rect 307666 172680 307722 172689
rect 307484 172644 307536 172650
rect 307666 172615 307722 172624
rect 307484 172586 307536 172592
rect 307680 172582 307708 172615
rect 307668 172576 307720 172582
rect 307668 172518 307720 172524
rect 307666 171864 307722 171873
rect 307666 171799 307722 171808
rect 307298 171456 307354 171465
rect 307298 171391 307354 171400
rect 307312 171154 307340 171391
rect 307680 171290 307708 171799
rect 307668 171284 307720 171290
rect 307668 171226 307720 171232
rect 307300 171148 307352 171154
rect 307300 171090 307352 171096
rect 307298 171048 307354 171057
rect 307298 170983 307354 170992
rect 307114 170232 307170 170241
rect 307114 170167 307170 170176
rect 307024 170128 307076 170134
rect 307024 170070 307076 170076
rect 307128 169046 307156 170167
rect 307312 169930 307340 170983
rect 307574 170640 307630 170649
rect 307574 170575 307630 170584
rect 307300 169924 307352 169930
rect 307300 169866 307352 169872
rect 307588 169862 307616 170575
rect 307576 169856 307628 169862
rect 307576 169798 307628 169804
rect 307666 169824 307722 169833
rect 307666 169759 307668 169768
rect 307720 169759 307722 169768
rect 307668 169730 307720 169736
rect 307482 169280 307538 169289
rect 307482 169215 307538 169224
rect 307116 169040 307168 169046
rect 307116 168982 307168 168988
rect 307496 168434 307524 169215
rect 307666 168872 307722 168881
rect 307666 168807 307722 168816
rect 307680 168502 307708 168807
rect 307668 168496 307720 168502
rect 307574 168464 307630 168473
rect 307484 168428 307536 168434
rect 307668 168438 307720 168444
rect 307574 168399 307630 168408
rect 307484 168370 307536 168376
rect 307482 168056 307538 168065
rect 307482 167991 307538 168000
rect 307496 167074 307524 167991
rect 307588 167686 307616 168399
rect 307576 167680 307628 167686
rect 307576 167622 307628 167628
rect 307666 167648 307722 167657
rect 307666 167583 307722 167592
rect 307574 167240 307630 167249
rect 307574 167175 307630 167184
rect 307484 167068 307536 167074
rect 307484 167010 307536 167016
rect 306746 166832 306802 166841
rect 306746 166767 306802 166776
rect 306760 165646 306788 166767
rect 307482 166424 307538 166433
rect 307482 166359 307538 166368
rect 306748 165640 306800 165646
rect 306748 165582 306800 165588
rect 307390 165472 307446 165481
rect 307390 165407 307446 165416
rect 307206 165064 307262 165073
rect 307206 164999 307262 165008
rect 307114 163024 307170 163033
rect 307114 162959 307170 162968
rect 307128 162926 307156 162959
rect 307116 162920 307168 162926
rect 307116 162862 307168 162868
rect 307114 159624 307170 159633
rect 307114 159559 307170 159568
rect 306746 159080 306802 159089
rect 306746 159015 306802 159024
rect 306760 158778 306788 159015
rect 307128 158914 307156 159559
rect 307116 158908 307168 158914
rect 307116 158850 307168 158856
rect 306748 158772 306800 158778
rect 306748 158714 306800 158720
rect 306562 158264 306618 158273
rect 306562 158199 306618 158208
rect 306576 157554 306604 158199
rect 306564 157548 306616 157554
rect 306564 157490 306616 157496
rect 306562 155680 306618 155689
rect 306562 155615 306618 155624
rect 306576 154630 306604 155615
rect 306564 154624 306616 154630
rect 306564 154566 306616 154572
rect 306930 154456 306986 154465
rect 306930 154391 306986 154400
rect 306746 154048 306802 154057
rect 306746 153983 306802 153992
rect 306654 151872 306710 151881
rect 306654 151807 306710 151816
rect 306668 149734 306696 151807
rect 306656 149728 306708 149734
rect 306656 149670 306708 149676
rect 306760 148374 306788 153983
rect 306944 153270 306972 154391
rect 306932 153264 306984 153270
rect 306932 153206 306984 153212
rect 307114 152688 307170 152697
rect 307114 152623 307170 152632
rect 306838 152280 306894 152289
rect 306838 152215 306894 152224
rect 306748 148368 306800 148374
rect 306748 148310 306800 148316
rect 306562 145888 306618 145897
rect 306562 145823 306618 145832
rect 306576 144974 306604 145823
rect 306852 145586 306880 152215
rect 307128 151842 307156 152623
rect 307116 151836 307168 151842
rect 307116 151778 307168 151784
rect 307114 148472 307170 148481
rect 307114 148407 307170 148416
rect 307022 148064 307078 148073
rect 307022 147999 307078 148008
rect 306840 145580 306892 145586
rect 306840 145522 306892 145528
rect 306564 144968 306616 144974
rect 306564 144910 306616 144916
rect 306562 144664 306618 144673
rect 306562 144599 306618 144608
rect 306576 143682 306604 144599
rect 307036 144158 307064 147999
rect 307128 147694 307156 148407
rect 307116 147688 307168 147694
rect 307116 147630 307168 147636
rect 307024 144152 307076 144158
rect 307024 144094 307076 144100
rect 306564 143676 306616 143682
rect 306564 143618 306616 143624
rect 306562 143032 306618 143041
rect 306562 142967 306618 142976
rect 306576 141506 306604 142967
rect 306930 142080 306986 142089
rect 306930 142015 306986 142024
rect 306564 141500 306616 141506
rect 306564 141442 306616 141448
rect 306944 140962 306972 142015
rect 307022 141672 307078 141681
rect 307022 141607 307078 141616
rect 306932 140956 306984 140962
rect 306932 140898 306984 140904
rect 306562 140448 306618 140457
rect 306562 140383 306618 140392
rect 306576 139534 306604 140383
rect 306564 139528 306616 139534
rect 306564 139470 306616 139476
rect 306562 139088 306618 139097
rect 306562 139023 306618 139032
rect 306576 138038 306604 139023
rect 306930 138680 306986 138689
rect 306930 138615 306986 138624
rect 306944 138174 306972 138615
rect 306932 138168 306984 138174
rect 306932 138110 306984 138116
rect 306564 138032 306616 138038
rect 306564 137974 306616 137980
rect 306562 136232 306618 136241
rect 306562 136167 306618 136176
rect 306576 135318 306604 136167
rect 307036 135930 307064 141607
rect 307114 137456 307170 137465
rect 307114 137391 307170 137400
rect 307128 136746 307156 137391
rect 307116 136740 307168 136746
rect 307116 136682 307168 136688
rect 307024 135924 307076 135930
rect 307024 135866 307076 135872
rect 306564 135312 306616 135318
rect 306564 135254 306616 135260
rect 307114 135280 307170 135289
rect 307114 135215 307170 135224
rect 307022 134056 307078 134065
rect 307022 133991 307078 134000
rect 306930 133648 306986 133657
rect 306930 133583 306986 133592
rect 306562 133240 306618 133249
rect 306562 133175 306618 133184
rect 306576 132530 306604 133175
rect 306944 132598 306972 133583
rect 306932 132592 306984 132598
rect 306932 132534 306984 132540
rect 306564 132524 306616 132530
rect 306564 132466 306616 132472
rect 305736 130416 305788 130422
rect 305736 130358 305788 130364
rect 306930 128888 306986 128897
rect 306930 128823 306986 128832
rect 306944 128450 306972 128823
rect 306932 128444 306984 128450
rect 306932 128386 306984 128392
rect 306746 122088 306802 122097
rect 306746 122023 306802 122032
rect 306760 121514 306788 122023
rect 306748 121508 306800 121514
rect 306748 121450 306800 121456
rect 306562 120048 306618 120057
rect 306562 119983 306618 119992
rect 305734 118960 305790 118969
rect 305734 118895 305790 118904
rect 305748 14550 305776 118895
rect 306576 118862 306604 119983
rect 306564 118856 306616 118862
rect 306564 118798 306616 118804
rect 305826 117600 305882 117609
rect 305826 117535 305882 117544
rect 305736 14544 305788 14550
rect 305736 14486 305788 14492
rect 305840 13122 305868 117535
rect 306562 114472 306618 114481
rect 306562 114407 306618 114416
rect 306576 113286 306604 114407
rect 306564 113280 306616 113286
rect 306564 113222 306616 113228
rect 306746 111072 306802 111081
rect 306746 111007 306802 111016
rect 306760 110634 306788 111007
rect 306748 110628 306800 110634
rect 306748 110570 306800 110576
rect 306930 109848 306986 109857
rect 306930 109783 306986 109792
rect 306944 109138 306972 109783
rect 306932 109132 306984 109138
rect 306932 109074 306984 109080
rect 305918 107944 305974 107953
rect 305918 107879 305974 107888
rect 305932 71058 305960 107879
rect 306746 106856 306802 106865
rect 306746 106791 306802 106800
rect 306760 106350 306788 106791
rect 306748 106344 306800 106350
rect 306748 106286 306800 106292
rect 306746 105496 306802 105505
rect 306746 105431 306802 105440
rect 306760 104922 306788 105431
rect 306748 104916 306800 104922
rect 306748 104858 306800 104864
rect 306930 104272 306986 104281
rect 306930 104207 306986 104216
rect 306746 103864 306802 103873
rect 306746 103799 306802 103808
rect 306760 103562 306788 103799
rect 306944 103630 306972 104207
rect 306932 103624 306984 103630
rect 306932 103566 306984 103572
rect 306748 103556 306800 103562
rect 306748 103498 306800 103504
rect 306562 102504 306618 102513
rect 306562 102439 306618 102448
rect 306576 102338 306604 102439
rect 306564 102332 306616 102338
rect 306564 102274 306616 102280
rect 306562 102096 306618 102105
rect 306562 102031 306618 102040
rect 306576 100910 306604 102031
rect 306564 100904 306616 100910
rect 306564 100846 306616 100852
rect 305920 71052 305972 71058
rect 305920 70994 305972 71000
rect 307036 68338 307064 133991
rect 307128 83502 307156 135215
rect 307220 134570 307248 164999
rect 307298 161664 307354 161673
rect 307298 161599 307354 161608
rect 307312 161498 307340 161599
rect 307300 161492 307352 161498
rect 307300 161434 307352 161440
rect 307298 160848 307354 160857
rect 307298 160783 307354 160792
rect 307312 153882 307340 160783
rect 307404 160750 307432 165407
rect 307496 163538 307524 166359
rect 307588 166326 307616 167175
rect 307680 167142 307708 167583
rect 307668 167136 307720 167142
rect 307668 167078 307720 167084
rect 307576 166320 307628 166326
rect 307576 166262 307628 166268
rect 307666 165880 307722 165889
rect 307666 165815 307722 165824
rect 307680 164898 307708 165815
rect 307668 164892 307720 164898
rect 307668 164834 307720 164840
rect 307574 164656 307630 164665
rect 307574 164591 307630 164600
rect 307588 164354 307616 164591
rect 307576 164348 307628 164354
rect 307576 164290 307628 164296
rect 307668 164280 307720 164286
rect 307666 164248 307668 164257
rect 307720 164248 307722 164257
rect 307666 164183 307722 164192
rect 307574 163840 307630 163849
rect 307574 163775 307630 163784
rect 307484 163532 307536 163538
rect 307484 163474 307536 163480
rect 307588 162994 307616 163775
rect 307666 163432 307722 163441
rect 307666 163367 307722 163376
rect 307680 163062 307708 163367
rect 307668 163056 307720 163062
rect 307668 162998 307720 163004
rect 307576 162988 307628 162994
rect 307576 162930 307628 162936
rect 307574 162480 307630 162489
rect 307574 162415 307630 162424
rect 307588 161634 307616 162415
rect 307666 162072 307722 162081
rect 307666 162007 307722 162016
rect 307576 161628 307628 161634
rect 307576 161570 307628 161576
rect 307680 161566 307708 162007
rect 307668 161560 307720 161566
rect 307668 161502 307720 161508
rect 307574 161256 307630 161265
rect 307574 161191 307630 161200
rect 307392 160744 307444 160750
rect 307392 160686 307444 160692
rect 307588 160206 307616 161191
rect 307666 160440 307722 160449
rect 307666 160375 307722 160384
rect 307576 160200 307628 160206
rect 307576 160142 307628 160148
rect 307680 160138 307708 160375
rect 307668 160132 307720 160138
rect 307668 160074 307720 160080
rect 307666 160032 307722 160041
rect 307666 159967 307722 159976
rect 307680 158846 307708 159967
rect 307668 158840 307720 158846
rect 307668 158782 307720 158788
rect 307574 158672 307630 158681
rect 307574 158607 307630 158616
rect 307390 157856 307446 157865
rect 307390 157791 307446 157800
rect 307404 155242 307432 157791
rect 307588 157418 307616 158607
rect 307668 157480 307720 157486
rect 307666 157448 307668 157457
rect 307720 157448 307722 157457
rect 307576 157412 307628 157418
rect 307666 157383 307722 157392
rect 307576 157354 307628 157360
rect 307482 157040 307538 157049
rect 307482 156975 307538 156984
rect 307496 156058 307524 156975
rect 307574 156632 307630 156641
rect 307574 156567 307630 156576
rect 307484 156052 307536 156058
rect 307484 155994 307536 156000
rect 307588 155990 307616 156567
rect 307666 156224 307722 156233
rect 307666 156159 307722 156168
rect 307680 156126 307708 156159
rect 307668 156120 307720 156126
rect 307668 156062 307720 156068
rect 307576 155984 307628 155990
rect 307576 155926 307628 155932
rect 307666 155272 307722 155281
rect 307392 155236 307444 155242
rect 307666 155207 307722 155216
rect 307392 155178 307444 155184
rect 307482 154864 307538 154873
rect 307482 154799 307538 154808
rect 307300 153876 307352 153882
rect 307300 153818 307352 153824
rect 307496 152522 307524 154799
rect 307680 154698 307708 155207
rect 307668 154692 307720 154698
rect 307668 154634 307720 154640
rect 307666 153640 307722 153649
rect 307666 153575 307722 153584
rect 307680 153338 307708 153575
rect 307668 153332 307720 153338
rect 307668 153274 307720 153280
rect 307666 153232 307722 153241
rect 307666 153167 307722 153176
rect 307680 152590 307708 153167
rect 307668 152584 307720 152590
rect 307668 152526 307720 152532
rect 307484 152516 307536 152522
rect 307484 152458 307536 152464
rect 307482 151464 307538 151473
rect 307482 151399 307538 151408
rect 307496 150550 307524 151399
rect 307666 151056 307722 151065
rect 307666 150991 307722 151000
rect 307574 150648 307630 150657
rect 307680 150618 307708 150991
rect 307574 150583 307630 150592
rect 307668 150612 307720 150618
rect 307484 150544 307536 150550
rect 307484 150486 307536 150492
rect 307588 150482 307616 150583
rect 307668 150554 307720 150560
rect 307576 150476 307628 150482
rect 307576 150418 307628 150424
rect 307574 150240 307630 150249
rect 307574 150175 307630 150184
rect 307588 149190 307616 150175
rect 307666 149288 307722 149297
rect 307666 149223 307722 149232
rect 307576 149184 307628 149190
rect 307576 149126 307628 149132
rect 307680 149122 307708 149223
rect 307668 149116 307720 149122
rect 307668 149058 307720 149064
rect 307390 148880 307446 148889
rect 307390 148815 307446 148824
rect 307298 145480 307354 145489
rect 307298 145415 307354 145424
rect 307208 134564 307260 134570
rect 307208 134506 307260 134512
rect 307312 122834 307340 145415
rect 307404 144294 307432 148815
rect 307482 147656 307538 147665
rect 307482 147591 307538 147600
rect 307496 146334 307524 147591
rect 307574 147248 307630 147257
rect 307574 147183 307630 147192
rect 307588 146470 307616 147183
rect 307666 146840 307722 146849
rect 307666 146775 307722 146784
rect 307680 146538 307708 146775
rect 307668 146532 307720 146538
rect 307668 146474 307720 146480
rect 307576 146464 307628 146470
rect 307576 146406 307628 146412
rect 307666 146432 307722 146441
rect 307666 146367 307668 146376
rect 307720 146367 307722 146376
rect 307668 146338 307720 146344
rect 307484 146328 307536 146334
rect 307484 146270 307536 146276
rect 307392 144288 307444 144294
rect 307392 144230 307444 144236
rect 307482 144256 307538 144265
rect 307482 144191 307538 144200
rect 307392 144152 307444 144158
rect 307392 144094 307444 144100
rect 307404 133210 307432 144094
rect 307496 142866 307524 144191
rect 307666 143848 307722 143857
rect 307666 143783 307722 143792
rect 307680 143614 307708 143783
rect 307668 143608 307720 143614
rect 307668 143550 307720 143556
rect 307574 143440 307630 143449
rect 307574 143375 307630 143384
rect 307484 142860 307536 142866
rect 307484 142802 307536 142808
rect 307588 142186 307616 143375
rect 307666 142488 307722 142497
rect 307666 142423 307722 142432
rect 307680 142254 307708 142423
rect 307668 142248 307720 142254
rect 307668 142190 307720 142196
rect 307576 142180 307628 142186
rect 307576 142122 307628 142128
rect 307574 141264 307630 141273
rect 307574 141199 307630 141208
rect 307588 140894 307616 141199
rect 307576 140888 307628 140894
rect 307576 140830 307628 140836
rect 307666 140856 307722 140865
rect 307666 140791 307668 140800
rect 307720 140791 307722 140800
rect 307668 140762 307720 140768
rect 307666 139632 307722 139641
rect 307666 139567 307722 139576
rect 307680 139466 307708 139567
rect 307668 139460 307720 139466
rect 307668 139402 307720 139408
rect 307666 138272 307722 138281
rect 307666 138207 307722 138216
rect 307680 138106 307708 138207
rect 307668 138100 307720 138106
rect 307668 138042 307720 138048
rect 307666 137864 307722 137873
rect 307666 137799 307722 137808
rect 307680 136678 307708 137799
rect 307668 136672 307720 136678
rect 307482 136640 307538 136649
rect 307668 136614 307720 136620
rect 307482 136575 307538 136584
rect 307496 135454 307524 136575
rect 307666 135688 307722 135697
rect 307666 135623 307722 135632
rect 307484 135448 307536 135454
rect 307484 135390 307536 135396
rect 307680 135386 307708 135623
rect 307668 135380 307720 135386
rect 307668 135322 307720 135328
rect 307574 134872 307630 134881
rect 307574 134807 307630 134816
rect 307588 134026 307616 134807
rect 307666 134464 307722 134473
rect 307666 134399 307722 134408
rect 307576 134020 307628 134026
rect 307576 133962 307628 133968
rect 307680 133958 307708 134399
rect 307668 133952 307720 133958
rect 307668 133894 307720 133900
rect 307392 133204 307444 133210
rect 307392 133146 307444 133152
rect 307482 132288 307538 132297
rect 307482 132223 307538 132232
rect 307496 131306 307524 132223
rect 307574 131880 307630 131889
rect 307574 131815 307630 131824
rect 307484 131300 307536 131306
rect 307484 131242 307536 131248
rect 307588 131238 307616 131815
rect 307666 131472 307722 131481
rect 307666 131407 307722 131416
rect 307576 131232 307628 131238
rect 307576 131174 307628 131180
rect 307680 131170 307708 131407
rect 307668 131164 307720 131170
rect 307668 131106 307720 131112
rect 307482 131064 307538 131073
rect 307482 130999 307538 131008
rect 307496 129878 307524 130999
rect 307574 129976 307630 129985
rect 307574 129911 307630 129920
rect 307668 129940 307720 129946
rect 307484 129872 307536 129878
rect 307484 129814 307536 129820
rect 307588 129810 307616 129911
rect 307668 129882 307720 129888
rect 307680 129849 307708 129882
rect 307666 129840 307722 129849
rect 307576 129804 307628 129810
rect 307666 129775 307722 129784
rect 307576 129746 307628 129752
rect 307666 129296 307722 129305
rect 307666 129231 307722 129240
rect 307680 128382 307708 129231
rect 307668 128376 307720 128382
rect 307668 128318 307720 128324
rect 307482 128072 307538 128081
rect 307482 128007 307538 128016
rect 307496 127090 307524 128007
rect 307574 127664 307630 127673
rect 307574 127599 307630 127608
rect 307484 127084 307536 127090
rect 307484 127026 307536 127032
rect 307588 127022 307616 127599
rect 307666 127256 307722 127265
rect 307666 127191 307722 127200
rect 307680 127158 307708 127191
rect 307668 127152 307720 127158
rect 307668 127094 307720 127100
rect 307576 127016 307628 127022
rect 307576 126958 307628 126964
rect 307574 126848 307630 126857
rect 307574 126783 307630 126792
rect 307588 125730 307616 126783
rect 307666 125760 307722 125769
rect 307576 125724 307628 125730
rect 307666 125695 307722 125704
rect 307576 125666 307628 125672
rect 307680 125662 307708 125695
rect 307668 125656 307720 125662
rect 307668 125598 307720 125604
rect 307482 125488 307538 125497
rect 307482 125423 307538 125432
rect 307496 124302 307524 125423
rect 307574 125080 307630 125089
rect 307574 125015 307630 125024
rect 307588 124370 307616 125015
rect 307666 124672 307722 124681
rect 307666 124607 307722 124616
rect 307680 124438 307708 124607
rect 307668 124432 307720 124438
rect 307668 124374 307720 124380
rect 307576 124364 307628 124370
rect 307576 124306 307628 124312
rect 307484 124296 307536 124302
rect 307484 124238 307536 124244
rect 307666 124264 307722 124273
rect 307666 124199 307668 124208
rect 307720 124199 307722 124208
rect 307668 124170 307720 124176
rect 307574 123448 307630 123457
rect 307574 123383 307630 123392
rect 307588 122874 307616 123383
rect 307666 123040 307722 123049
rect 307666 122975 307722 122984
rect 307680 122942 307708 122975
rect 307668 122936 307720 122942
rect 307668 122878 307720 122884
rect 307220 122806 307340 122834
rect 307576 122868 307628 122874
rect 307576 122810 307628 122816
rect 307220 119406 307248 122806
rect 307574 122496 307630 122505
rect 307574 122431 307630 122440
rect 307588 121650 307616 122431
rect 307666 121680 307722 121689
rect 307576 121644 307628 121650
rect 307666 121615 307722 121624
rect 307576 121586 307628 121592
rect 307680 121582 307708 121615
rect 307668 121576 307720 121582
rect 307668 121518 307720 121524
rect 307298 121272 307354 121281
rect 307298 121207 307354 121216
rect 307312 120290 307340 121207
rect 307574 120864 307630 120873
rect 307574 120799 307630 120808
rect 307300 120284 307352 120290
rect 307300 120226 307352 120232
rect 307588 120154 307616 120799
rect 307666 120456 307722 120465
rect 307666 120391 307722 120400
rect 307680 120222 307708 120391
rect 307668 120216 307720 120222
rect 307668 120158 307720 120164
rect 307576 120148 307628 120154
rect 307576 120090 307628 120096
rect 307666 119640 307722 119649
rect 307666 119575 307722 119584
rect 307208 119400 307260 119406
rect 307208 119342 307260 119348
rect 307680 118794 307708 119575
rect 307668 118788 307720 118794
rect 307668 118730 307720 118736
rect 307574 118688 307630 118697
rect 307574 118623 307630 118632
rect 307298 118280 307354 118289
rect 307298 118215 307354 118224
rect 307312 117366 307340 118215
rect 307588 117434 307616 118623
rect 307668 117564 307720 117570
rect 307668 117506 307720 117512
rect 307680 117473 307708 117506
rect 307666 117464 307722 117473
rect 307576 117428 307628 117434
rect 307666 117399 307722 117408
rect 307576 117370 307628 117376
rect 307300 117360 307352 117366
rect 307300 117302 307352 117308
rect 307482 117056 307538 117065
rect 307482 116991 307538 117000
rect 307496 116006 307524 116991
rect 307574 116648 307630 116657
rect 307574 116583 307630 116592
rect 307588 116074 307616 116583
rect 307666 116240 307722 116249
rect 307666 116175 307722 116184
rect 307680 116142 307708 116175
rect 307668 116136 307720 116142
rect 307668 116078 307720 116084
rect 307576 116068 307628 116074
rect 307576 116010 307628 116016
rect 307484 116000 307536 116006
rect 307484 115942 307536 115948
rect 307298 115696 307354 115705
rect 307298 115631 307354 115640
rect 307312 114578 307340 115631
rect 307574 115288 307630 115297
rect 307574 115223 307630 115232
rect 307588 114714 307616 115223
rect 307666 114880 307722 114889
rect 307666 114815 307722 114824
rect 307576 114708 307628 114714
rect 307576 114650 307628 114656
rect 307680 114646 307708 114815
rect 307668 114640 307720 114646
rect 307668 114582 307720 114588
rect 307300 114572 307352 114578
rect 307300 114514 307352 114520
rect 307666 113248 307722 113257
rect 307666 113183 307668 113192
rect 307720 113183 307722 113192
rect 307668 113154 307720 113160
rect 307482 112704 307538 112713
rect 307482 112639 307538 112648
rect 307496 111858 307524 112639
rect 307574 112296 307630 112305
rect 307574 112231 307630 112240
rect 307588 111926 307616 112231
rect 307668 111988 307720 111994
rect 307668 111930 307720 111936
rect 307576 111920 307628 111926
rect 307680 111897 307708 111930
rect 307576 111862 307628 111868
rect 307666 111888 307722 111897
rect 307484 111852 307536 111858
rect 307666 111823 307722 111832
rect 307484 111794 307536 111800
rect 307298 111480 307354 111489
rect 307298 111415 307354 111424
rect 307312 110566 307340 111415
rect 307666 110664 307722 110673
rect 307666 110599 307722 110608
rect 307300 110560 307352 110566
rect 307300 110502 307352 110508
rect 307680 110498 307708 110599
rect 307668 110492 307720 110498
rect 307668 110434 307720 110440
rect 307574 110256 307630 110265
rect 307574 110191 307630 110200
rect 307588 109206 307616 110191
rect 307666 109304 307722 109313
rect 307666 109239 307722 109248
rect 307576 109200 307628 109206
rect 307576 109142 307628 109148
rect 307680 109070 307708 109239
rect 307668 109064 307720 109070
rect 307668 109006 307720 109012
rect 307482 108896 307538 108905
rect 307482 108831 307538 108840
rect 307496 107914 307524 108831
rect 307484 107908 307536 107914
rect 307484 107850 307536 107856
rect 307574 107808 307630 107817
rect 307574 107743 307630 107752
rect 307668 107772 307720 107778
rect 307588 107710 307616 107743
rect 307668 107714 307720 107720
rect 307576 107704 307628 107710
rect 307680 107681 307708 107714
rect 307576 107646 307628 107652
rect 307666 107672 307722 107681
rect 307666 107607 307722 107616
rect 307666 107264 307722 107273
rect 307666 107199 307722 107208
rect 307680 106486 307708 107199
rect 307668 106480 307720 106486
rect 307482 106448 307538 106457
rect 307668 106422 307720 106428
rect 307482 106383 307484 106392
rect 307536 106383 307538 106392
rect 307484 106354 307536 106360
rect 307574 105904 307630 105913
rect 307574 105839 307630 105848
rect 307588 105058 307616 105839
rect 307666 105088 307722 105097
rect 307576 105052 307628 105058
rect 307666 105023 307722 105032
rect 307576 104994 307628 105000
rect 307680 104990 307708 105023
rect 307668 104984 307720 104990
rect 307668 104926 307720 104932
rect 307482 104680 307538 104689
rect 307482 104615 307538 104624
rect 307496 103698 307524 104615
rect 307484 103692 307536 103698
rect 307484 103634 307536 103640
rect 307574 103456 307630 103465
rect 307574 103391 307630 103400
rect 307588 102202 307616 103391
rect 307666 103048 307722 103057
rect 307666 102983 307722 102992
rect 307680 102270 307708 102983
rect 307668 102264 307720 102270
rect 307668 102206 307720 102212
rect 307576 102196 307628 102202
rect 307576 102138 307628 102144
rect 307482 101688 307538 101697
rect 307482 101623 307538 101632
rect 307496 100774 307524 101623
rect 307574 101280 307630 101289
rect 307574 101215 307630 101224
rect 307588 100842 307616 101215
rect 307668 100972 307720 100978
rect 307668 100914 307720 100920
rect 307680 100881 307708 100914
rect 307666 100872 307722 100881
rect 307576 100836 307628 100842
rect 307666 100807 307722 100816
rect 307576 100778 307628 100784
rect 307484 100768 307536 100774
rect 307484 100710 307536 100716
rect 307482 100464 307538 100473
rect 307482 100399 307538 100408
rect 307496 99550 307524 100399
rect 307574 100056 307630 100065
rect 307574 99991 307630 100000
rect 307484 99544 307536 99550
rect 307484 99486 307536 99492
rect 307588 99482 307616 99991
rect 307666 99648 307722 99657
rect 307666 99583 307722 99592
rect 307576 99476 307628 99482
rect 307576 99418 307628 99424
rect 307680 99414 307708 99583
rect 307668 99408 307720 99414
rect 307668 99350 307720 99356
rect 307574 99104 307630 99113
rect 307574 99039 307630 99048
rect 307298 98288 307354 98297
rect 307298 98223 307354 98232
rect 307312 98054 307340 98223
rect 307588 98122 307616 99039
rect 307666 98696 307722 98705
rect 307666 98631 307722 98640
rect 307680 98190 307708 98631
rect 307668 98184 307720 98190
rect 307668 98126 307720 98132
rect 307576 98116 307628 98122
rect 307576 98058 307628 98064
rect 307300 98048 307352 98054
rect 307300 97990 307352 97996
rect 307206 97880 307262 97889
rect 307206 97815 307262 97824
rect 307116 83496 307168 83502
rect 307116 83438 307168 83444
rect 307024 68332 307076 68338
rect 307024 68274 307076 68280
rect 307220 54534 307248 97815
rect 307574 97472 307630 97481
rect 307574 97407 307630 97416
rect 307390 97064 307446 97073
rect 307390 96999 307446 97008
rect 307404 55894 307432 96999
rect 307588 96694 307616 97407
rect 307668 96756 307720 96762
rect 307668 96698 307720 96704
rect 307576 96688 307628 96694
rect 307680 96665 307708 96698
rect 307576 96630 307628 96636
rect 307666 96656 307722 96665
rect 307666 96591 307722 96600
rect 307666 96248 307722 96257
rect 307666 96183 307722 96192
rect 307680 95266 307708 96183
rect 307668 95260 307720 95266
rect 307668 95202 307720 95208
rect 307392 55888 307444 55894
rect 307392 55830 307444 55836
rect 307208 54528 307260 54534
rect 307208 54470 307260 54476
rect 307760 37256 307812 37262
rect 307760 37198 307812 37204
rect 305828 13116 305880 13122
rect 305828 13058 305880 13064
rect 305644 9648 305696 9654
rect 305644 9590 305696 9596
rect 305656 6914 305684 9590
rect 306748 7608 306800 7614
rect 306748 7550 306800 7556
rect 305564 6886 305684 6914
rect 305564 480 305592 6886
rect 306760 480 306788 7550
rect 307772 3534 307800 37198
rect 308416 3942 308444 385018
rect 308496 356108 308548 356114
rect 308496 356050 308548 356056
rect 308508 87718 308536 356050
rect 337382 349752 337438 349761
rect 337382 349687 337438 349696
rect 309784 338836 309836 338842
rect 309784 338778 309836 338784
rect 309140 333260 309192 333266
rect 309140 333202 309192 333208
rect 308588 170128 308640 170134
rect 308588 170070 308640 170076
rect 308496 87712 308548 87718
rect 308496 87654 308548 87660
rect 308496 83632 308548 83638
rect 308496 83574 308548 83580
rect 308508 37262 308536 83574
rect 308496 37256 308548 37262
rect 308496 37198 308548 37204
rect 308600 6798 308628 170070
rect 309152 101833 309180 333202
rect 309322 114064 309378 114073
rect 309322 113999 309378 114008
rect 309336 113121 309364 113999
rect 309322 113112 309378 113121
rect 309322 113047 309378 113056
rect 309138 101824 309194 101833
rect 309138 101759 309194 101768
rect 308588 6792 308640 6798
rect 308588 6734 308640 6740
rect 308404 3936 308456 3942
rect 308404 3878 308456 3884
rect 307760 3528 307812 3534
rect 307760 3470 307812 3476
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 303130 -960 303242 326
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 354 308026 480
rect 308600 354 308628 6734
rect 309796 4010 309824 338778
rect 320824 336796 320876 336802
rect 320824 336738 320876 336744
rect 315304 303816 315356 303822
rect 315304 303758 315356 303764
rect 313922 293992 313978 294001
rect 313922 293927 313978 293936
rect 311164 293276 311216 293282
rect 311164 293218 311216 293224
rect 311176 180266 311204 293218
rect 312544 266484 312596 266490
rect 312544 266426 312596 266432
rect 311164 180260 311216 180266
rect 311164 180202 311216 180208
rect 312556 175982 312584 266426
rect 312636 204944 312688 204950
rect 312636 204886 312688 204892
rect 312648 177449 312676 204886
rect 312634 177440 312690 177449
rect 313936 177410 313964 293927
rect 314016 228540 314068 228546
rect 314016 228482 314068 228488
rect 314028 180470 314056 228482
rect 314108 214736 314160 214742
rect 314108 214678 314160 214684
rect 314016 180464 314068 180470
rect 314016 180406 314068 180412
rect 314120 177546 314148 214678
rect 314108 177540 314160 177546
rect 314108 177482 314160 177488
rect 312634 177375 312690 177384
rect 313924 177404 313976 177410
rect 313924 177346 313976 177352
rect 315316 176050 315344 303758
rect 318064 303748 318116 303754
rect 318064 303690 318116 303696
rect 316684 277432 316736 277438
rect 316684 277374 316736 277380
rect 315396 216028 315448 216034
rect 315396 215970 315448 215976
rect 315408 176118 315436 215970
rect 316696 182918 316724 277374
rect 316776 252612 316828 252618
rect 316776 252554 316828 252560
rect 316684 182912 316736 182918
rect 316684 182854 316736 182860
rect 316788 180402 316816 252554
rect 316776 180396 316828 180402
rect 316776 180338 316828 180344
rect 318076 178673 318104 303690
rect 319444 278792 319496 278798
rect 319444 278734 319496 278740
rect 318156 243704 318208 243710
rect 318156 243646 318208 243652
rect 318062 178664 318118 178673
rect 318062 178599 318118 178608
rect 318168 177478 318196 243646
rect 318248 199504 318300 199510
rect 318248 199446 318300 199452
rect 318156 177472 318208 177478
rect 318156 177414 318208 177420
rect 316038 176760 316094 176769
rect 316038 176695 316094 176704
rect 315396 176112 315448 176118
rect 315396 176054 315448 176060
rect 315304 176044 315356 176050
rect 315304 175986 315356 175992
rect 312544 175976 312596 175982
rect 316052 175930 316080 176695
rect 318260 175953 318288 199446
rect 318340 185632 318392 185638
rect 318340 185574 318392 185580
rect 318352 177614 318380 185574
rect 318340 177608 318392 177614
rect 318340 177550 318392 177556
rect 312544 175918 312596 175924
rect 316020 175902 316080 175930
rect 318246 175944 318302 175953
rect 318246 175879 318302 175888
rect 319456 175642 319484 278734
rect 320836 267034 320864 336738
rect 325700 302252 325752 302258
rect 325700 302194 325752 302200
rect 322940 284436 322992 284442
rect 322940 284378 322992 284384
rect 320824 267028 320876 267034
rect 320824 266970 320876 266976
rect 321560 264240 321612 264246
rect 321560 264182 321612 264188
rect 321284 184272 321336 184278
rect 321284 184214 321336 184220
rect 319444 175636 319496 175642
rect 319444 175578 319496 175584
rect 321296 172689 321324 184214
rect 321468 175636 321520 175642
rect 321468 175578 321520 175584
rect 321480 175273 321508 175578
rect 321466 175264 321522 175273
rect 321466 175199 321522 175208
rect 321282 172680 321338 172689
rect 321282 172615 321338 172624
rect 321572 141953 321600 264182
rect 321652 240780 321704 240786
rect 321652 240722 321704 240728
rect 321558 141944 321614 141953
rect 321558 141879 321614 141888
rect 321664 119921 321692 240722
rect 321744 195424 321796 195430
rect 321744 195366 321796 195372
rect 321650 119912 321706 119921
rect 321650 119847 321706 119856
rect 321756 104553 321784 195366
rect 321836 187128 321888 187134
rect 321836 187070 321888 187076
rect 321848 170649 321876 187070
rect 321834 170640 321890 170649
rect 321834 170575 321890 170584
rect 322952 160177 322980 284378
rect 323032 260228 323084 260234
rect 323032 260170 323084 260176
rect 322938 160168 322994 160177
rect 322938 160103 322994 160112
rect 323044 137873 323072 260170
rect 323124 209160 323176 209166
rect 323124 209102 323176 209108
rect 323030 137864 323086 137873
rect 323030 137799 323086 137808
rect 323136 121689 323164 209102
rect 324320 188352 324372 188358
rect 324320 188294 324372 188300
rect 323216 178900 323268 178906
rect 323216 178842 323268 178848
rect 323228 147801 323256 178842
rect 324332 174049 324360 188294
rect 324412 178832 324464 178838
rect 324412 178774 324464 178780
rect 324318 174040 324374 174049
rect 324318 173975 324374 173984
rect 324320 173868 324372 173874
rect 324320 173810 324372 173816
rect 324332 173233 324360 173810
rect 324318 173224 324374 173233
rect 324318 173159 324374 173168
rect 324320 171080 324372 171086
rect 324320 171022 324372 171028
rect 324332 170921 324360 171022
rect 324318 170912 324374 170921
rect 324318 170847 324374 170856
rect 324320 168360 324372 168366
rect 324320 168302 324372 168308
rect 324332 167113 324360 168302
rect 324424 167793 324452 178774
rect 324504 178764 324556 178770
rect 324504 178706 324556 178712
rect 324516 168609 324544 178706
rect 324502 168600 324558 168609
rect 324502 168535 324558 168544
rect 324410 167784 324466 167793
rect 324410 167719 324466 167728
rect 324318 167104 324374 167113
rect 324318 167039 324374 167048
rect 324320 167000 324372 167006
rect 324320 166942 324372 166948
rect 324332 166297 324360 166942
rect 324318 166288 324374 166297
rect 324318 166223 324374 166232
rect 324412 165572 324464 165578
rect 324412 165514 324464 165520
rect 324320 165504 324372 165510
rect 324318 165472 324320 165481
rect 324372 165472 324374 165481
rect 324318 165407 324374 165416
rect 324424 164801 324452 165514
rect 324410 164792 324466 164801
rect 324410 164727 324466 164736
rect 324412 164212 324464 164218
rect 324412 164154 324464 164160
rect 324320 164144 324372 164150
rect 324320 164086 324372 164092
rect 324332 163985 324360 164086
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324424 163169 324452 164154
rect 324410 163160 324466 163169
rect 324410 163095 324466 163104
rect 324320 162852 324372 162858
rect 324320 162794 324372 162800
rect 324332 162489 324360 162794
rect 324412 162784 324464 162790
rect 324412 162726 324464 162732
rect 324318 162480 324374 162489
rect 324318 162415 324374 162424
rect 324424 161673 324452 162726
rect 324410 161664 324466 161673
rect 324410 161599 324466 161608
rect 324320 161424 324372 161430
rect 324320 161366 324372 161372
rect 324332 160857 324360 161366
rect 324318 160848 324374 160857
rect 324318 160783 324374 160792
rect 324320 160064 324372 160070
rect 324320 160006 324372 160012
rect 324332 159361 324360 160006
rect 324318 159352 324374 159361
rect 324318 159287 324374 159296
rect 324412 158704 324464 158710
rect 324412 158646 324464 158652
rect 324320 158636 324372 158642
rect 324320 158578 324372 158584
rect 324332 158545 324360 158578
rect 324318 158536 324374 158545
rect 324318 158471 324374 158480
rect 324424 157865 324452 158646
rect 324410 157856 324466 157865
rect 324410 157791 324466 157800
rect 324320 157344 324372 157350
rect 324320 157286 324372 157292
rect 324332 157049 324360 157286
rect 324318 157040 324374 157049
rect 324318 156975 324374 156984
rect 324320 156868 324372 156874
rect 324320 156810 324372 156816
rect 324332 156369 324360 156810
rect 324318 156360 324374 156369
rect 324318 156295 324374 156304
rect 324412 155916 324464 155922
rect 324412 155858 324464 155864
rect 324320 155848 324372 155854
rect 324320 155790 324372 155796
rect 324332 155553 324360 155790
rect 324318 155544 324374 155553
rect 324318 155479 324374 155488
rect 324424 154737 324452 155858
rect 324410 154728 324466 154737
rect 324410 154663 324466 154672
rect 324412 154488 324464 154494
rect 324412 154430 324464 154436
rect 324320 154352 324372 154358
rect 324320 154294 324372 154300
rect 324332 154057 324360 154294
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 324424 153241 324452 154430
rect 324410 153232 324466 153241
rect 324320 153196 324372 153202
rect 324410 153167 324466 153176
rect 324320 153138 324372 153144
rect 324332 152425 324360 153138
rect 324318 152416 324374 152425
rect 324318 152351 324374 152360
rect 324320 151768 324372 151774
rect 324318 151736 324320 151745
rect 324372 151736 324374 151745
rect 324318 151671 324374 151680
rect 324412 151700 324464 151706
rect 324412 151642 324464 151648
rect 324424 150929 324452 151642
rect 324410 150920 324466 150929
rect 324410 150855 324466 150864
rect 324320 150408 324372 150414
rect 324320 150350 324372 150356
rect 324332 150113 324360 150350
rect 324318 150104 324374 150113
rect 324318 150039 324374 150048
rect 324320 149796 324372 149802
rect 324320 149738 324372 149744
rect 324332 149433 324360 149738
rect 324318 149424 324374 149433
rect 324318 149359 324374 149368
rect 324320 149048 324372 149054
rect 324320 148990 324372 148996
rect 324332 148617 324360 148990
rect 324318 148608 324374 148617
rect 324318 148543 324374 148552
rect 323214 147792 323270 147801
rect 323214 147727 323270 147736
rect 324320 147620 324372 147626
rect 324320 147562 324372 147568
rect 324332 147121 324360 147562
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 325712 146962 325740 302194
rect 331864 299532 331916 299538
rect 331864 299474 331916 299480
rect 328460 288448 328512 288454
rect 328460 288390 328512 288396
rect 325792 287088 325844 287094
rect 325792 287030 325844 287036
rect 325804 147082 325832 287030
rect 327080 262268 327132 262274
rect 327080 262210 327132 262216
rect 325884 210588 325936 210594
rect 325884 210530 325936 210536
rect 325792 147076 325844 147082
rect 325792 147018 325844 147024
rect 325712 146934 325832 146962
rect 325700 146872 325752 146878
rect 325700 146814 325752 146820
rect 324318 146296 324374 146305
rect 324318 146231 324320 146240
rect 324372 146231 324374 146240
rect 324320 146202 324372 146208
rect 324412 146192 324464 146198
rect 324412 146134 324464 146140
rect 324424 145489 324452 146134
rect 324410 145480 324466 145489
rect 324410 145415 324466 145424
rect 324320 144900 324372 144906
rect 324320 144842 324372 144848
rect 324332 143993 324360 144842
rect 324318 143984 324374 143993
rect 324318 143919 324374 143928
rect 324320 143472 324372 143478
rect 324320 143414 324372 143420
rect 324332 143177 324360 143414
rect 324318 143168 324374 143177
rect 324318 143103 324374 143112
rect 325606 142488 325662 142497
rect 325712 142474 325740 146814
rect 325662 142446 325740 142474
rect 325606 142423 325662 142432
rect 324320 142112 324372 142118
rect 324320 142054 324372 142060
rect 324332 140865 324360 142054
rect 324318 140856 324374 140865
rect 324318 140791 324374 140800
rect 324320 140752 324372 140758
rect 324320 140694 324372 140700
rect 324332 140185 324360 140694
rect 324318 140176 324374 140185
rect 324318 140111 324374 140120
rect 324412 139392 324464 139398
rect 324318 139360 324374 139369
rect 324412 139334 324464 139340
rect 324318 139295 324320 139304
rect 324372 139295 324374 139304
rect 324320 139266 324372 139272
rect 324424 138553 324452 139334
rect 324410 138544 324466 138553
rect 324410 138479 324466 138488
rect 324320 137964 324372 137970
rect 324320 137906 324372 137912
rect 324332 137057 324360 137906
rect 324318 137048 324374 137057
rect 324318 136983 324374 136992
rect 324320 136604 324372 136610
rect 324320 136546 324372 136552
rect 324332 136377 324360 136546
rect 324318 136368 324374 136377
rect 324318 136303 324374 136312
rect 325606 136096 325662 136105
rect 325804 136082 325832 146934
rect 325662 136054 325832 136082
rect 325606 136031 325662 136040
rect 324320 133884 324372 133890
rect 324320 133826 324372 133832
rect 324332 133249 324360 133826
rect 324318 133240 324374 133249
rect 324318 133175 324374 133184
rect 324964 132524 325016 132530
rect 324964 132466 325016 132472
rect 324412 132456 324464 132462
rect 324318 132424 324374 132433
rect 324412 132398 324464 132404
rect 324318 132359 324320 132368
rect 324372 132359 324374 132368
rect 324320 132330 324372 132336
rect 324424 131753 324452 132398
rect 324410 131744 324466 131753
rect 324410 131679 324466 131688
rect 324320 131096 324372 131102
rect 324320 131038 324372 131044
rect 324332 130937 324360 131038
rect 324412 131028 324464 131034
rect 324412 130970 324464 130976
rect 324318 130928 324374 130937
rect 324318 130863 324374 130872
rect 324424 130121 324452 130970
rect 324410 130112 324466 130121
rect 324410 130047 324466 130056
rect 324320 129736 324372 129742
rect 324320 129678 324372 129684
rect 324332 129441 324360 129678
rect 324412 129668 324464 129674
rect 324412 129610 324464 129616
rect 324318 129432 324374 129441
rect 324318 129367 324374 129376
rect 324424 128625 324452 129610
rect 324410 128616 324466 128625
rect 324410 128551 324466 128560
rect 324320 128308 324372 128314
rect 324320 128250 324372 128256
rect 324332 127809 324360 128250
rect 324412 128240 324464 128246
rect 324412 128182 324464 128188
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324424 127129 324452 128182
rect 324410 127120 324466 127129
rect 324410 127055 324466 127064
rect 324320 125588 324372 125594
rect 324320 125530 324372 125536
rect 324332 125497 324360 125530
rect 324412 125520 324464 125526
rect 324318 125488 324374 125497
rect 324412 125462 324464 125468
rect 324318 125423 324374 125432
rect 324424 124817 324452 125462
rect 324410 124808 324466 124817
rect 324410 124743 324466 124752
rect 324320 124160 324372 124166
rect 324320 124102 324372 124108
rect 324332 124001 324360 124102
rect 324318 123992 324374 124001
rect 324318 123927 324374 123936
rect 324976 123185 325004 132466
rect 324962 123176 325018 123185
rect 324962 123111 325018 123120
rect 324320 122800 324372 122806
rect 324320 122742 324372 122748
rect 324332 122505 324360 122742
rect 324318 122496 324374 122505
rect 324318 122431 324374 122440
rect 323122 121680 323178 121689
rect 323122 121615 323178 121624
rect 324320 121440 324372 121446
rect 324320 121382 324372 121388
rect 324332 120873 324360 121382
rect 324412 121372 324464 121378
rect 324412 121314 324464 121320
rect 324318 120864 324374 120873
rect 324318 120799 324374 120808
rect 324424 120193 324452 121314
rect 324410 120184 324466 120193
rect 324410 120119 324466 120128
rect 324320 118652 324372 118658
rect 324320 118594 324372 118600
rect 324332 118561 324360 118594
rect 324412 118584 324464 118590
rect 324318 118552 324374 118561
rect 324412 118526 324464 118532
rect 324318 118487 324374 118496
rect 324424 117881 324452 118526
rect 324410 117872 324466 117881
rect 324410 117807 324466 117816
rect 324320 117292 324372 117298
rect 324320 117234 324372 117240
rect 324332 116385 324360 117234
rect 324318 116376 324374 116385
rect 324318 116311 324374 116320
rect 324320 115932 324372 115938
rect 324320 115874 324372 115880
rect 324332 115569 324360 115874
rect 324412 115864 324464 115870
rect 324412 115806 324464 115812
rect 324318 115560 324374 115569
rect 324318 115495 324374 115504
rect 324424 114753 324452 115806
rect 324410 114744 324466 114753
rect 324410 114679 324466 114688
rect 324320 114436 324372 114442
rect 324320 114378 324372 114384
rect 321834 113656 321890 113665
rect 321834 113591 321890 113600
rect 321742 104544 321798 104553
rect 321742 104479 321798 104488
rect 321742 102232 321798 102241
rect 321742 102167 321798 102176
rect 321650 101144 321706 101153
rect 321650 101079 321706 101088
rect 321374 99648 321430 99657
rect 321374 99583 321430 99592
rect 321388 95130 321416 99583
rect 321466 97336 321522 97345
rect 321466 97271 321522 97280
rect 321480 96558 321508 97271
rect 321558 96656 321614 96665
rect 321558 96591 321614 96600
rect 321468 96552 321520 96558
rect 321468 96494 321520 96500
rect 321572 95198 321600 96591
rect 321560 95192 321612 95198
rect 321560 95134 321612 95140
rect 321376 95124 321428 95130
rect 321376 95066 321428 95072
rect 321664 94994 321692 101079
rect 321652 94988 321704 94994
rect 321652 94930 321704 94936
rect 320824 94512 320876 94518
rect 320824 94454 320876 94460
rect 311900 90432 311952 90438
rect 311898 90400 311900 90409
rect 311952 90400 311954 90409
rect 311898 90335 311954 90344
rect 315304 89004 315356 89010
rect 315304 88946 315356 88952
rect 316684 89004 316736 89010
rect 316684 88946 316736 88952
rect 309876 80708 309928 80714
rect 309876 80650 309928 80656
rect 309888 6798 309916 80650
rect 310518 78024 310574 78033
rect 310518 77959 310520 77968
rect 310572 77959 310574 77968
rect 310520 77930 310572 77936
rect 309968 29640 310020 29646
rect 309968 29582 310020 29588
rect 309980 6798 310008 29582
rect 315316 13802 315344 88946
rect 316132 33108 316184 33114
rect 316132 33050 316184 33056
rect 314660 13796 314712 13802
rect 314660 13738 314712 13744
rect 315304 13796 315356 13802
rect 315304 13738 315356 13744
rect 312634 11792 312690 11801
rect 312634 11727 312690 11736
rect 311438 11656 311494 11665
rect 311438 11591 311494 11600
rect 309876 6792 309928 6798
rect 309876 6734 309928 6740
rect 309968 6792 310020 6798
rect 309968 6734 310020 6740
rect 309784 4004 309836 4010
rect 309784 3946 309836 3952
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309060 480 309088 3470
rect 307914 326 308628 354
rect 307914 -960 308026 326
rect 309018 -960 309130 480
rect 309980 354 310008 6734
rect 311452 480 311480 11591
rect 312648 480 312676 11727
rect 313832 3460 313884 3466
rect 313832 3402 313884 3408
rect 313844 480 313872 3402
rect 310214 354 310326 480
rect 309980 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314672 354 314700 13738
rect 316144 3534 316172 33050
rect 316696 3874 316724 88946
rect 319444 84856 319496 84862
rect 319444 84798 319496 84804
rect 317420 82136 317472 82142
rect 317420 82078 317472 82084
rect 316776 44872 316828 44878
rect 316776 44814 316828 44820
rect 316788 33114 316816 44814
rect 316776 33108 316828 33114
rect 316776 33050 316828 33056
rect 317432 16574 317460 82078
rect 318890 43480 318946 43489
rect 318890 43415 318946 43424
rect 317432 16546 318104 16574
rect 316224 3868 316276 3874
rect 316224 3810 316276 3816
rect 316684 3868 316736 3874
rect 316684 3810 316736 3816
rect 316132 3528 316184 3534
rect 316132 3470 316184 3476
rect 316236 480 316264 3810
rect 317328 3528 317380 3534
rect 317328 3470 317380 3476
rect 317340 480 317368 3470
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 318904 3466 318932 43415
rect 319456 16574 319484 84798
rect 320088 43512 320140 43518
rect 320086 43480 320088 43489
rect 320140 43480 320142 43489
rect 320086 43415 320142 43424
rect 320836 16574 320864 94454
rect 321756 92478 321784 102167
rect 321848 94926 321876 113591
rect 324332 113257 324360 114378
rect 324318 113248 324374 113257
rect 324318 113183 324374 113192
rect 325896 113174 325924 210530
rect 325976 187196 326028 187202
rect 325976 187138 326028 187144
rect 325988 154358 326016 187138
rect 326066 178664 326122 178673
rect 326066 178599 326122 178608
rect 326080 171329 326108 178599
rect 326066 171320 326122 171329
rect 326066 171255 326122 171264
rect 325976 154352 326028 154358
rect 325976 154294 326028 154300
rect 327092 132530 327120 262210
rect 327264 251252 327316 251258
rect 327264 251194 327316 251200
rect 327172 221604 327224 221610
rect 327172 221546 327224 221552
rect 327080 132524 327132 132530
rect 327080 132466 327132 132472
rect 324320 113144 324372 113150
rect 324320 113086 324372 113092
rect 325712 113146 325924 113174
rect 324332 112441 324360 113086
rect 324318 112432 324374 112441
rect 324318 112367 324374 112376
rect 322938 111752 322994 111761
rect 322938 111687 322994 111696
rect 321926 102776 321982 102785
rect 321926 102711 321982 102720
rect 321836 94920 321888 94926
rect 321836 94862 321888 94868
rect 321744 92472 321796 92478
rect 321744 92414 321796 92420
rect 321940 92410 321968 102711
rect 322952 95062 322980 111687
rect 324320 110424 324372 110430
rect 324320 110366 324372 110372
rect 324332 109449 324360 110366
rect 324318 109440 324374 109449
rect 324318 109375 324374 109384
rect 324320 108996 324372 109002
rect 324320 108938 324372 108944
rect 324332 108633 324360 108938
rect 324318 108624 324374 108633
rect 324318 108559 324374 108568
rect 325606 107808 325662 107817
rect 325712 107794 325740 113146
rect 325662 107766 325740 107794
rect 325606 107743 325662 107752
rect 327184 105874 327212 221546
rect 327276 149802 327304 251194
rect 327356 188420 327408 188426
rect 327356 188362 327408 188368
rect 327368 156874 327396 188362
rect 327356 156868 327408 156874
rect 327356 156810 327408 156816
rect 327264 149796 327316 149802
rect 327264 149738 327316 149744
rect 328472 140758 328500 288390
rect 328552 244928 328604 244934
rect 328552 244870 328604 244876
rect 328460 140752 328512 140758
rect 328460 140694 328512 140700
rect 328564 125594 328592 244870
rect 331220 240168 331272 240174
rect 331220 240110 331272 240116
rect 328644 225616 328696 225622
rect 328644 225558 328696 225564
rect 328656 154494 328684 225558
rect 329932 213376 329984 213382
rect 329932 213318 329984 213324
rect 328736 196716 328788 196722
rect 328736 196658 328788 196664
rect 328644 154488 328696 154494
rect 328644 154430 328696 154436
rect 328748 131034 328776 196658
rect 329840 177608 329892 177614
rect 329840 177550 329892 177556
rect 329852 168366 329880 177550
rect 329840 168360 329892 168366
rect 329840 168302 329892 168308
rect 329944 136610 329972 213318
rect 330116 210452 330168 210458
rect 330116 210394 330168 210400
rect 330024 176112 330076 176118
rect 330024 176054 330076 176060
rect 330036 165510 330064 176054
rect 330024 165504 330076 165510
rect 330024 165446 330076 165452
rect 329932 136604 329984 136610
rect 329932 136546 329984 136552
rect 328736 131028 328788 131034
rect 328736 130970 328788 130976
rect 330128 128246 330156 210394
rect 331232 129674 331260 240110
rect 331312 229832 331364 229838
rect 331312 229774 331364 229780
rect 331220 129668 331272 129674
rect 331220 129610 331272 129616
rect 331324 128314 331352 229774
rect 331496 180464 331548 180470
rect 331496 180406 331548 180412
rect 331404 175976 331456 175982
rect 331404 175918 331456 175924
rect 331416 158642 331444 175918
rect 331508 164150 331536 180406
rect 331876 178770 331904 299474
rect 333980 295384 334032 295390
rect 333980 295326 334032 295332
rect 332600 238060 332652 238066
rect 332600 238002 332652 238008
rect 331864 178764 331916 178770
rect 331864 178706 331916 178712
rect 331496 164144 331548 164150
rect 331496 164086 331548 164092
rect 331404 158636 331456 158642
rect 331404 158578 331456 158584
rect 332612 151706 332640 238002
rect 333336 224256 333388 224262
rect 333336 224198 333388 224204
rect 333244 180328 333296 180334
rect 333244 180270 333296 180276
rect 332692 177540 332744 177546
rect 332692 177482 332744 177488
rect 332600 151700 332652 151706
rect 332600 151642 332652 151648
rect 331864 150476 331916 150482
rect 331864 150418 331916 150424
rect 331312 128308 331364 128314
rect 331312 128250 331364 128256
rect 330116 128240 330168 128246
rect 330116 128182 330168 128188
rect 328552 125588 328604 125594
rect 328552 125530 328604 125536
rect 324320 105868 324372 105874
rect 324320 105810 324372 105816
rect 327172 105868 327224 105874
rect 327172 105810 327224 105816
rect 324332 105505 324360 105810
rect 324318 105496 324374 105505
rect 324318 105431 324374 105440
rect 323030 104816 323086 104825
rect 323030 104751 323086 104760
rect 323044 96626 323072 104751
rect 330484 104168 330536 104174
rect 330484 104110 330536 104116
rect 326344 101448 326396 101454
rect 326344 101390 326396 101396
rect 324410 100872 324466 100881
rect 324410 100807 324466 100816
rect 323584 100020 323636 100026
rect 323584 99962 323636 99968
rect 323032 96620 323084 96626
rect 323032 96562 323084 96568
rect 322940 95056 322992 95062
rect 322940 94998 322992 95004
rect 321928 92404 321980 92410
rect 321928 92346 321980 92352
rect 322204 86284 322256 86290
rect 322204 86226 322256 86232
rect 322216 42770 322244 86226
rect 322204 42764 322256 42770
rect 322204 42706 322256 42712
rect 322216 41478 322244 42706
rect 321560 41472 321612 41478
rect 321560 41414 321612 41420
rect 322204 41472 322256 41478
rect 322204 41414 322256 41420
rect 321572 16574 321600 41414
rect 319456 16546 319760 16574
rect 320836 16546 320956 16574
rect 321572 16546 322152 16574
rect 319732 3942 319760 16546
rect 320928 4010 320956 16546
rect 320916 4004 320968 4010
rect 320916 3946 320968 3952
rect 319720 3936 319772 3942
rect 319720 3878 319772 3884
rect 318892 3460 318944 3466
rect 318892 3402 318944 3408
rect 319732 480 319760 3878
rect 320928 480 320956 3946
rect 322124 480 322152 16546
rect 323596 6914 323624 99962
rect 324320 95940 324372 95946
rect 324320 95882 324372 95888
rect 324332 16574 324360 95882
rect 324424 89622 324452 100807
rect 324412 89616 324464 89622
rect 324412 89558 324464 89564
rect 324964 87712 325016 87718
rect 324964 87654 325016 87660
rect 324976 76566 325004 87654
rect 326356 80034 326384 101390
rect 325700 80028 325752 80034
rect 325700 79970 325752 79976
rect 326344 80028 326396 80034
rect 326344 79970 326396 79976
rect 324964 76560 325016 76566
rect 324964 76502 325016 76508
rect 324332 16546 324452 16574
rect 323320 6886 323624 6914
rect 323320 4078 323348 6886
rect 323308 4072 323360 4078
rect 323308 4014 323360 4020
rect 323320 480 323348 4014
rect 324424 480 324452 16546
rect 324976 3534 325004 76502
rect 325712 16574 325740 79970
rect 330496 77246 330524 104110
rect 331220 83564 331272 83570
rect 331220 83506 331272 83512
rect 329840 77240 329892 77246
rect 329840 77182 329892 77188
rect 330484 77240 330536 77246
rect 330484 77182 330536 77188
rect 327080 32428 327132 32434
rect 327080 32370 327132 32376
rect 327092 16574 327120 32370
rect 329852 16574 329880 77182
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 324964 3528 325016 3534
rect 324964 3470 325016 3476
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 329196 3528 329248 3534
rect 329196 3470 329248 3476
rect 329208 480 329236 3470
rect 330404 480 330432 16546
rect 331232 3534 331260 83506
rect 331876 43450 331904 150418
rect 332704 137970 332732 177482
rect 332692 137964 332744 137970
rect 332692 137906 332744 137912
rect 331956 87644 332008 87650
rect 331956 87586 332008 87592
rect 331864 43444 331916 43450
rect 331864 43386 331916 43392
rect 331968 6914 331996 87586
rect 332598 66872 332654 66881
rect 332598 66807 332654 66816
rect 332612 66162 332640 66807
rect 332600 66156 332652 66162
rect 332600 66098 332652 66104
rect 331600 6886 331996 6914
rect 331600 4078 331628 6886
rect 331588 4072 331640 4078
rect 331588 4014 331640 4020
rect 331220 3528 331272 3534
rect 331220 3470 331272 3476
rect 331600 480 331628 4014
rect 332612 3534 332640 66098
rect 333256 4146 333284 180270
rect 333348 114510 333376 224198
rect 333992 173874 334020 295326
rect 335360 276072 335412 276078
rect 335360 276014 335412 276020
rect 334164 200796 334216 200802
rect 334164 200738 334216 200744
rect 334072 181688 334124 181694
rect 334072 181630 334124 181636
rect 333980 173868 334032 173874
rect 333980 173810 334032 173816
rect 333428 140820 333480 140826
rect 333428 140762 333480 140768
rect 333336 114504 333388 114510
rect 333336 114446 333388 114452
rect 333440 84862 333468 140762
rect 334084 139330 334112 181630
rect 334176 160070 334204 200738
rect 334256 176044 334308 176050
rect 334256 175986 334308 175992
rect 334268 171086 334296 175986
rect 334256 171080 334308 171086
rect 334256 171022 334308 171028
rect 334624 169788 334676 169794
rect 334624 169730 334676 169736
rect 334164 160064 334216 160070
rect 334164 160006 334216 160012
rect 334072 139324 334124 139330
rect 334072 139266 334124 139272
rect 333428 84856 333480 84862
rect 333428 84798 333480 84804
rect 334636 65618 334664 169730
rect 334716 146328 334768 146334
rect 334716 146270 334768 146276
rect 334728 83638 334756 146270
rect 335372 144906 335400 276014
rect 336096 211880 336148 211886
rect 336096 211822 336148 211828
rect 335452 184408 335504 184414
rect 335452 184350 335504 184356
rect 335464 162790 335492 184350
rect 335542 175944 335598 175953
rect 335542 175879 335598 175888
rect 335556 167006 335584 175879
rect 335544 167000 335596 167006
rect 335544 166942 335596 166948
rect 335452 162784 335504 162790
rect 335452 162726 335504 162732
rect 336004 158772 336056 158778
rect 336004 158714 336056 158720
rect 335360 144900 335412 144906
rect 335360 144842 335412 144848
rect 334716 83632 334768 83638
rect 334716 83574 334768 83580
rect 335360 73160 335412 73166
rect 335360 73102 335412 73108
rect 334624 65612 334676 65618
rect 334624 65554 334676 65560
rect 334072 46232 334124 46238
rect 334070 46200 334072 46209
rect 334124 46200 334126 46209
rect 334070 46135 334126 46144
rect 335372 16574 335400 73102
rect 336016 45558 336044 158714
rect 336108 135250 336136 211822
rect 336740 185768 336792 185774
rect 336740 185710 336792 185716
rect 336752 150414 336780 185710
rect 336832 177472 336884 177478
rect 336832 177414 336884 177420
rect 336844 157350 336872 177414
rect 336832 157344 336884 157350
rect 336832 157286 336884 157292
rect 336740 150408 336792 150414
rect 336740 150350 336792 150356
rect 336096 135244 336148 135250
rect 336096 135186 336148 135192
rect 337396 95198 337424 349687
rect 347044 347064 347096 347070
rect 347044 347006 347096 347012
rect 340144 324964 340196 324970
rect 340144 324906 340196 324912
rect 338120 267776 338172 267782
rect 338120 267718 338172 267724
rect 337476 200864 337528 200870
rect 337476 200806 337528 200812
rect 337488 113082 337516 200806
rect 338132 113150 338160 267718
rect 339592 238128 339644 238134
rect 339592 238070 339644 238076
rect 339500 228472 339552 228478
rect 339500 228414 339552 228420
rect 338212 211812 338264 211818
rect 338212 211754 338264 211760
rect 338224 164218 338252 211754
rect 338304 184204 338356 184210
rect 338304 184146 338356 184152
rect 338212 164212 338264 164218
rect 338212 164154 338264 164160
rect 338316 151774 338344 184146
rect 338764 177336 338816 177342
rect 338764 177278 338816 177284
rect 338304 151768 338356 151774
rect 338304 151710 338356 151716
rect 338120 113144 338172 113150
rect 338120 113086 338172 113092
rect 337476 113076 337528 113082
rect 337476 113018 337528 113024
rect 337384 95192 337436 95198
rect 337384 95134 337436 95140
rect 337396 94722 337424 95134
rect 336740 94716 336792 94722
rect 336740 94658 336792 94664
rect 337384 94716 337436 94722
rect 337384 94658 337436 94664
rect 336096 84856 336148 84862
rect 336096 84798 336148 84804
rect 336108 73166 336136 84798
rect 336096 73160 336148 73166
rect 336096 73102 336148 73108
rect 336004 45552 336056 45558
rect 336004 45494 336056 45500
rect 336752 16574 336780 94658
rect 338776 73098 338804 177278
rect 339512 139398 339540 228414
rect 339604 165578 339632 238070
rect 339684 182912 339736 182918
rect 339684 182854 339736 182860
rect 339592 165572 339644 165578
rect 339592 165514 339644 165520
rect 339696 155854 339724 182854
rect 339684 155848 339736 155854
rect 339684 155790 339736 155796
rect 339500 139392 339552 139398
rect 339500 139334 339552 139340
rect 340156 86970 340184 324906
rect 345664 323604 345716 323610
rect 345664 323546 345716 323552
rect 344284 300144 344336 300150
rect 344284 300086 344336 300092
rect 342258 296848 342314 296857
rect 342258 296783 342314 296792
rect 340878 295352 340934 295361
rect 340878 295287 340934 295296
rect 340236 164280 340288 164286
rect 340236 164222 340288 164228
rect 339500 86964 339552 86970
rect 339500 86906 339552 86912
rect 340144 86964 340196 86970
rect 340144 86906 340196 86912
rect 338764 73092 338816 73098
rect 338764 73034 338816 73040
rect 338776 71806 338804 73034
rect 338120 71800 338172 71806
rect 338120 71742 338172 71748
rect 338764 71800 338816 71806
rect 338764 71742 338816 71748
rect 338132 16574 338160 71742
rect 335372 16546 336320 16574
rect 336752 16546 337056 16574
rect 338132 16546 338712 16574
rect 335082 11792 335138 11801
rect 335082 11727 335138 11736
rect 332692 4140 332744 4146
rect 332692 4082 332744 4088
rect 333244 4140 333296 4146
rect 333244 4082 333296 4088
rect 332600 3528 332652 3534
rect 332600 3470 332652 3476
rect 332704 480 332732 4082
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 333900 480 333928 3470
rect 335096 480 335124 11727
rect 336292 480 336320 16546
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337028 354 337056 16546
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 86906
rect 340248 47598 340276 164222
rect 340892 161430 340920 295287
rect 340972 235272 341024 235278
rect 340972 235214 341024 235220
rect 340880 161424 340932 161430
rect 340880 161366 340932 161372
rect 340984 117298 341012 235214
rect 341156 180396 341208 180402
rect 341156 180338 341208 180344
rect 341064 177404 341116 177410
rect 341064 177346 341116 177352
rect 340972 117292 341024 117298
rect 340972 117234 341024 117240
rect 341076 110430 341104 177346
rect 341168 153202 341196 180338
rect 341524 157412 341576 157418
rect 341524 157354 341576 157360
rect 341156 153196 341208 153202
rect 341156 153138 341208 153144
rect 341064 110424 341116 110430
rect 341064 110366 341116 110372
rect 340880 49088 340932 49094
rect 340880 49030 340932 49036
rect 340236 47592 340288 47598
rect 340236 47534 340288 47540
rect 339868 8968 339920 8974
rect 339868 8910 339920 8916
rect 339880 4078 339908 8910
rect 339868 4072 339920 4078
rect 339868 4014 339920 4020
rect 340892 3534 340920 49030
rect 341536 49026 341564 157354
rect 342272 122806 342300 296783
rect 342352 282940 342404 282946
rect 342352 282882 342404 282888
rect 342364 132394 342392 282882
rect 342996 227044 343048 227050
rect 342996 226986 343048 226992
rect 342444 178764 342496 178770
rect 342444 178706 342496 178712
rect 342456 162858 342484 178706
rect 342444 162852 342496 162858
rect 342444 162794 342496 162800
rect 342904 161492 342956 161498
rect 342904 161434 342956 161440
rect 342352 132388 342404 132394
rect 342352 132330 342404 132336
rect 342260 122800 342312 122806
rect 342260 122742 342312 122748
rect 342350 87680 342406 87689
rect 342350 87615 342352 87624
rect 342404 87615 342406 87624
rect 342352 87586 342404 87592
rect 341524 49020 341576 49026
rect 341524 48962 341576 48968
rect 342916 42702 342944 161434
rect 343008 125594 343036 226986
rect 343640 191208 343692 191214
rect 343640 191150 343692 191156
rect 342996 125588 343048 125594
rect 342996 125530 343048 125536
rect 343652 115870 343680 191150
rect 343732 181552 343784 181558
rect 343732 181494 343784 181500
rect 343744 143478 343772 181494
rect 343824 180260 343876 180266
rect 343824 180202 343876 180208
rect 343836 158710 343864 180202
rect 343824 158704 343876 158710
rect 343824 158646 343876 158652
rect 343732 143472 343784 143478
rect 343732 143414 343784 143420
rect 343640 115864 343692 115870
rect 343640 115806 343692 115812
rect 344296 48278 344324 300086
rect 345112 291304 345164 291310
rect 345112 291246 345164 291252
rect 345020 184068 345072 184074
rect 345020 184010 345072 184016
rect 343640 48272 343692 48278
rect 343640 48214 343692 48220
rect 344284 48272 344336 48278
rect 344284 48214 344336 48220
rect 342996 43444 343048 43450
rect 342996 43386 343048 43392
rect 342904 42696 342956 42702
rect 342904 42638 342956 42644
rect 343008 4146 343036 43386
rect 343652 16574 343680 48214
rect 345032 16574 345060 184010
rect 345124 125526 345152 291246
rect 345204 248464 345256 248470
rect 345204 248406 345256 248412
rect 345112 125520 345164 125526
rect 345112 125462 345164 125468
rect 345216 109002 345244 248406
rect 345296 186992 345348 186998
rect 345296 186934 345348 186940
rect 345308 155922 345336 186934
rect 345676 184074 345704 323546
rect 346400 238808 346452 238814
rect 346400 238750 346452 238756
rect 345664 184068 345716 184074
rect 345664 184010 345716 184016
rect 345676 183598 345704 184010
rect 345664 183592 345716 183598
rect 345664 183534 345716 183540
rect 345296 155916 345348 155922
rect 345296 155858 345348 155864
rect 345664 142180 345716 142186
rect 345664 142122 345716 142128
rect 345204 108996 345256 109002
rect 345204 108938 345256 108944
rect 345676 89010 345704 142122
rect 346412 133890 346440 238750
rect 346492 192568 346544 192574
rect 346492 192510 346544 192516
rect 346504 146198 346532 192510
rect 346492 146192 346544 146198
rect 346492 146134 346544 146140
rect 346400 133884 346452 133890
rect 346400 133826 346452 133832
rect 345664 89004 345716 89010
rect 345664 88946 345716 88952
rect 343652 16546 344600 16574
rect 345032 16546 345336 16574
rect 343362 11792 343418 11801
rect 343362 11727 343418 11736
rect 342996 4140 343048 4146
rect 342996 4082 343048 4088
rect 340880 3528 340932 3534
rect 342168 3528 342220 3534
rect 340880 3470 340932 3476
rect 340970 3496 341026 3505
rect 340970 3431 341026 3440
rect 342074 3496 342130 3505
rect 342168 3470 342220 3476
rect 342074 3431 342076 3440
rect 340984 480 341012 3431
rect 342128 3431 342130 3440
rect 342076 3402 342128 3408
rect 342180 480 342208 3470
rect 343376 480 343404 11727
rect 344572 480 344600 16546
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 347056 6914 347084 347006
rect 349804 320884 349856 320890
rect 349804 320826 349856 320832
rect 347780 300960 347832 300966
rect 347780 300902 347832 300908
rect 347792 121378 347820 300902
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 349160 258120 349212 258126
rect 349160 258062 349212 258068
rect 347872 231192 347924 231198
rect 347872 231134 347924 231140
rect 347780 121372 347832 121378
rect 347780 121314 347832 121320
rect 347884 118590 347912 231134
rect 348422 174584 348478 174593
rect 348422 174519 348478 174528
rect 347872 118584 347924 118590
rect 347872 118526 347924 118532
rect 348436 89690 348464 174519
rect 349172 131102 349200 258062
rect 349264 149054 349292 266358
rect 349344 203652 349396 203658
rect 349344 203594 349396 203600
rect 349252 149048 349304 149054
rect 349252 148990 349304 148996
rect 349160 131096 349212 131102
rect 349160 131038 349212 131044
rect 349356 114442 349384 203594
rect 349344 114436 349396 114442
rect 349344 114378 349396 114384
rect 348424 89684 348476 89690
rect 348424 89626 348476 89632
rect 348436 89282 348464 89626
rect 347780 89276 347832 89282
rect 347780 89218 347832 89224
rect 348424 89276 348476 89282
rect 348424 89218 348476 89224
rect 347792 16574 347820 89218
rect 349816 52426 349844 320826
rect 351920 318096 351972 318102
rect 351920 318038 351972 318044
rect 350540 300892 350592 300898
rect 350540 300834 350592 300840
rect 350552 147626 350580 300834
rect 351184 267028 351236 267034
rect 351184 266970 351236 266976
rect 350632 189848 350684 189854
rect 350632 189790 350684 189796
rect 350540 147620 350592 147626
rect 350540 147562 350592 147568
rect 350644 115938 350672 189790
rect 350632 115932 350684 115938
rect 350632 115874 350684 115880
rect 349804 52420 349856 52426
rect 349804 52362 349856 52368
rect 349816 51134 349844 52362
rect 349160 51128 349212 51134
rect 349160 51070 349212 51076
rect 349804 51128 349856 51134
rect 349804 51070 349856 51076
rect 349172 16574 349200 51070
rect 347792 16546 348096 16574
rect 349172 16546 349292 16574
rect 346964 6886 347084 6914
rect 346964 4078 346992 6886
rect 346952 4072 347004 4078
rect 346952 4014 347004 4020
rect 346964 480 346992 4014
rect 348068 480 348096 16546
rect 349264 480 349292 16546
rect 351196 4146 351224 266970
rect 351932 96558 351960 318038
rect 356060 311908 356112 311914
rect 356060 311850 356112 311856
rect 353392 291236 353444 291242
rect 353392 291178 353444 291184
rect 353300 280220 353352 280226
rect 353300 280162 353352 280168
rect 352012 232620 352064 232626
rect 352012 232562 352064 232568
rect 352024 129742 352052 232562
rect 352104 193860 352156 193866
rect 352104 193802 352156 193808
rect 352012 129736 352064 129742
rect 352012 129678 352064 129684
rect 352116 121446 352144 193802
rect 352564 155984 352616 155990
rect 352564 155926 352616 155932
rect 352104 121440 352156 121446
rect 352104 121382 352156 121388
rect 351920 96552 351972 96558
rect 351920 96494 351972 96500
rect 351932 95946 351960 96494
rect 351920 95940 351972 95946
rect 351920 95882 351972 95888
rect 352576 46306 352604 155926
rect 353312 124166 353340 280162
rect 353404 146266 353432 291178
rect 354036 207664 354088 207670
rect 354036 207606 354088 207612
rect 353944 171148 353996 171154
rect 353944 171090 353996 171096
rect 353392 146260 353444 146266
rect 353392 146202 353444 146208
rect 353300 124160 353352 124166
rect 353300 124102 353352 124108
rect 352656 90364 352708 90370
rect 352656 90306 352708 90312
rect 352564 46300 352616 46306
rect 352564 46242 352616 46248
rect 351184 4140 351236 4146
rect 351184 4082 351236 4088
rect 351644 4140 351696 4146
rect 351644 4082 351696 4088
rect 350448 3528 350500 3534
rect 350448 3470 350500 3476
rect 350460 480 350488 3470
rect 351656 480 351684 4082
rect 352668 4078 352696 90306
rect 353956 13734 353984 171090
rect 354048 103494 354076 207606
rect 354680 187060 354732 187066
rect 354680 187002 354732 187008
rect 354692 118658 354720 187002
rect 355324 173936 355376 173942
rect 355324 173878 355376 173884
rect 354680 118652 354732 118658
rect 354680 118594 354732 118600
rect 354036 103488 354088 103494
rect 354036 103430 354088 103436
rect 355336 78062 355364 173878
rect 356072 142118 356100 311850
rect 356704 176724 356756 176730
rect 356704 176666 356756 176672
rect 356060 142112 356112 142118
rect 356060 142054 356112 142060
rect 355324 78056 355376 78062
rect 355324 77998 355376 78004
rect 356716 50590 356744 176666
rect 356796 154624 356848 154630
rect 356796 154566 356848 154572
rect 356704 50584 356756 50590
rect 356704 50526 356756 50532
rect 356808 33046 356836 154566
rect 357452 33114 357480 400182
rect 357532 294024 357584 294030
rect 357532 293966 357584 293972
rect 357544 132462 357572 293966
rect 358084 143608 358136 143614
rect 358084 143550 358136 143556
rect 357532 132456 357584 132462
rect 357532 132398 357584 132404
rect 358096 90438 358124 143550
rect 358084 90432 358136 90438
rect 358084 90374 358136 90380
rect 358832 49706 358860 401610
rect 360844 383716 360896 383722
rect 360844 383658 360896 383664
rect 359464 153264 359516 153270
rect 359464 153206 359516 153212
rect 358820 49700 358872 49706
rect 358820 49642 358872 49648
rect 359280 49700 359332 49706
rect 359280 49642 359332 49648
rect 359292 49094 359320 49642
rect 359280 49088 359332 49094
rect 359280 49030 359332 49036
rect 357440 33108 357492 33114
rect 357440 33050 357492 33056
rect 356796 33040 356848 33046
rect 356796 32982 356848 32988
rect 357452 32434 357480 33050
rect 357440 32428 357492 32434
rect 357440 32370 357492 32376
rect 353944 13728 353996 13734
rect 353944 13670 353996 13676
rect 359476 4826 359504 153206
rect 360856 11014 360884 383658
rect 377404 340196 377456 340202
rect 377404 340138 377456 340144
rect 367744 305040 367796 305046
rect 367744 304982 367796 304988
rect 360936 178084 360988 178090
rect 360936 178026 360988 178032
rect 360948 51882 360976 178026
rect 363604 149116 363656 149122
rect 363604 149058 363656 149064
rect 360936 51876 360988 51882
rect 360936 51818 360988 51824
rect 363616 16590 363644 149058
rect 367756 111790 367784 304982
rect 370504 243636 370556 243642
rect 370504 243578 370556 243584
rect 367744 111784 367796 111790
rect 367744 111726 367796 111732
rect 370516 97986 370544 243578
rect 371884 221536 371936 221542
rect 371884 221478 371936 221484
rect 371896 106282 371924 221478
rect 374644 147688 374696 147694
rect 374644 147630 374696 147636
rect 371884 106276 371936 106282
rect 371884 106218 371936 106224
rect 370504 97980 370556 97986
rect 370504 97922 370556 97928
rect 363604 16584 363656 16590
rect 363604 16526 363656 16532
rect 360844 11008 360896 11014
rect 360844 10950 360896 10956
rect 359464 4820 359516 4826
rect 359464 4762 359516 4768
rect 352656 4072 352708 4078
rect 352656 4014 352708 4020
rect 360856 3534 360884 10950
rect 374656 9654 374684 147630
rect 376024 136672 376076 136678
rect 376024 136614 376076 136620
rect 376036 101454 376064 136614
rect 377416 128314 377444 340138
rect 395344 313336 395396 313342
rect 395344 313278 395396 313284
rect 378784 296744 378836 296750
rect 378784 296686 378836 296692
rect 378796 133890 378824 296686
rect 382924 286340 382976 286346
rect 382924 286282 382976 286288
rect 381544 238264 381596 238270
rect 381544 238206 381596 238212
rect 378784 133884 378836 133890
rect 378784 133826 378836 133832
rect 377404 128308 377456 128314
rect 377404 128250 377456 128256
rect 376024 101448 376076 101454
rect 376024 101390 376076 101396
rect 381556 96626 381584 238206
rect 382936 102134 382964 286282
rect 388444 263628 388496 263634
rect 388444 263570 388496 263576
rect 385684 180872 385736 180878
rect 385684 180814 385736 180820
rect 382924 102128 382976 102134
rect 382924 102070 382976 102076
rect 381544 96620 381596 96626
rect 381544 96562 381596 96568
rect 385696 66162 385724 180814
rect 388456 99346 388484 263570
rect 393964 231124 394016 231130
rect 393964 231066 394016 231072
rect 392584 205012 392636 205018
rect 392584 204954 392636 204960
rect 389824 180192 389876 180198
rect 389824 180134 389876 180140
rect 389836 100638 389864 180134
rect 389824 100632 389876 100638
rect 389824 100574 389876 100580
rect 388444 99340 388496 99346
rect 388444 99282 388496 99288
rect 392596 97918 392624 204954
rect 393976 99278 394004 231066
rect 395356 104854 395384 313278
rect 410524 312588 410576 312594
rect 410524 312530 410576 312536
rect 407764 280832 407816 280838
rect 407764 280774 407816 280780
rect 406384 275392 406436 275398
rect 406384 275334 406436 275340
rect 399484 256080 399536 256086
rect 399484 256022 399536 256028
rect 396724 214600 396776 214606
rect 396724 214542 396776 214548
rect 395344 104848 395396 104854
rect 395344 104790 395396 104796
rect 393964 99272 394016 99278
rect 393964 99214 394016 99220
rect 396736 99210 396764 214542
rect 399496 122806 399524 256022
rect 400864 253224 400916 253230
rect 400864 253166 400916 253172
rect 399484 122800 399536 122806
rect 399484 122742 399536 122748
rect 400876 120086 400904 253166
rect 403624 232552 403676 232558
rect 403624 232494 403676 232500
rect 403636 199510 403664 232494
rect 403624 199504 403676 199510
rect 403624 199446 403676 199452
rect 403624 135312 403676 135318
rect 403624 135254 403676 135260
rect 400864 120080 400916 120086
rect 400864 120022 400916 120028
rect 403636 104174 403664 135254
rect 406396 126954 406424 275334
rect 407776 180062 407804 280774
rect 407764 180056 407816 180062
rect 407764 179998 407816 180004
rect 408408 180056 408460 180062
rect 408408 179998 408460 180004
rect 408420 179450 408448 179998
rect 408408 179444 408460 179450
rect 408408 179386 408460 179392
rect 408420 129742 408448 179386
rect 410536 132462 410564 312530
rect 419540 298784 419592 298790
rect 419540 298726 419592 298732
rect 417424 272536 417476 272542
rect 417424 272478 417476 272484
rect 414664 262948 414716 262954
rect 414664 262890 414716 262896
rect 413284 242208 413336 242214
rect 413284 242150 413336 242156
rect 411904 139460 411956 139466
rect 411904 139402 411956 139408
rect 410524 132456 410576 132462
rect 410524 132398 410576 132404
rect 408408 129736 408460 129742
rect 408408 129678 408460 129684
rect 406384 126948 406436 126954
rect 406384 126890 406436 126896
rect 403624 104168 403676 104174
rect 403624 104110 403676 104116
rect 411916 100026 411944 139402
rect 413296 107642 413324 242150
rect 414676 118658 414704 262890
rect 416778 178664 416834 178673
rect 416778 178599 416834 178608
rect 416792 178090 416820 178599
rect 416780 178084 416832 178090
rect 416780 178026 416832 178032
rect 416778 177032 416834 177041
rect 416778 176967 416834 176976
rect 416792 176730 416820 176967
rect 416780 176724 416832 176730
rect 416780 176666 416832 176672
rect 416778 175264 416834 175273
rect 416778 175199 416834 175208
rect 416792 173942 416820 175199
rect 416780 173936 416832 173942
rect 416780 173878 416832 173884
rect 416778 171864 416834 171873
rect 416778 171799 416834 171808
rect 416792 171154 416820 171799
rect 416780 171148 416832 171154
rect 416780 171090 416832 171096
rect 416778 170232 416834 170241
rect 416778 170167 416834 170176
rect 416792 169794 416820 170167
rect 416780 169788 416832 169794
rect 416780 169730 416832 169736
rect 416778 165064 416834 165073
rect 416778 164999 416834 165008
rect 416792 164286 416820 164999
rect 416780 164280 416832 164286
rect 416780 164222 416832 164228
rect 416778 161800 416834 161809
rect 416778 161735 416834 161744
rect 416792 161498 416820 161735
rect 416780 161492 416832 161498
rect 416780 161434 416832 161440
rect 416778 160032 416834 160041
rect 416778 159967 416834 159976
rect 416792 158778 416820 159967
rect 416780 158772 416832 158778
rect 416780 158714 416832 158720
rect 416778 158400 416834 158409
rect 416778 158335 416834 158344
rect 416792 157418 416820 158335
rect 416780 157412 416832 157418
rect 416780 157354 416832 157360
rect 416778 156632 416834 156641
rect 416778 156567 416834 156576
rect 416792 155990 416820 156567
rect 416780 155984 416832 155990
rect 416780 155926 416832 155932
rect 416778 155000 416834 155009
rect 416778 154935 416834 154944
rect 416792 154630 416820 154935
rect 416780 154624 416832 154630
rect 416780 154566 416832 154572
rect 416780 153264 416832 153270
rect 416778 153232 416780 153241
rect 416832 153232 416834 153241
rect 416778 153167 416834 153176
rect 416778 151600 416834 151609
rect 416778 151535 416834 151544
rect 416792 150482 416820 151535
rect 416780 150476 416832 150482
rect 416780 150418 416832 150424
rect 416778 149832 416834 149841
rect 416778 149767 416834 149776
rect 416792 149122 416820 149767
rect 416780 149116 416832 149122
rect 416780 149058 416832 149064
rect 416778 148200 416834 148209
rect 416778 148135 416834 148144
rect 416792 147694 416820 148135
rect 416780 147688 416832 147694
rect 416780 147630 416832 147636
rect 416778 146568 416834 146577
rect 416778 146503 416834 146512
rect 416792 146334 416820 146503
rect 416780 146328 416832 146334
rect 416780 146270 416832 146276
rect 416778 144800 416834 144809
rect 416778 144735 416834 144744
rect 416792 143614 416820 144735
rect 416780 143608 416832 143614
rect 416780 143550 416832 143556
rect 416778 143168 416834 143177
rect 416778 143103 416834 143112
rect 416792 142186 416820 143103
rect 416780 142180 416832 142186
rect 416780 142122 416832 142128
rect 416778 141400 416834 141409
rect 416778 141335 416834 141344
rect 416792 140826 416820 141335
rect 416780 140820 416832 140826
rect 416780 140762 416832 140768
rect 416778 139768 416834 139777
rect 416778 139703 416834 139712
rect 416792 139466 416820 139703
rect 416780 139460 416832 139466
rect 416780 139402 416832 139408
rect 416778 138000 416834 138009
rect 416778 137935 416834 137944
rect 416792 136678 416820 137935
rect 416780 136672 416832 136678
rect 416780 136614 416832 136620
rect 416778 136368 416834 136377
rect 416778 136303 416834 136312
rect 416792 135318 416820 136303
rect 416780 135312 416832 135318
rect 416780 135254 416832 135260
rect 417332 135244 417384 135250
rect 417332 135186 417384 135192
rect 417344 134609 417372 135186
rect 417330 134600 417386 134609
rect 417330 134535 417386 134544
rect 416780 129736 416832 129742
rect 416780 129678 416832 129684
rect 416792 129577 416820 129678
rect 416778 129568 416834 129577
rect 416778 129503 416834 129512
rect 416780 120080 416832 120086
rect 416780 120022 416832 120028
rect 416792 119377 416820 120022
rect 416778 119368 416834 119377
rect 416778 119303 416834 119312
rect 414664 118652 414716 118658
rect 414664 118594 414716 118600
rect 416964 118652 417016 118658
rect 416964 118594 417016 118600
rect 416976 117745 417004 118594
rect 416962 117736 417018 117745
rect 416962 117671 417018 117680
rect 416780 114504 416832 114510
rect 416780 114446 416832 114452
rect 416792 114345 416820 114446
rect 416778 114336 416834 114345
rect 416778 114271 416834 114280
rect 416780 113076 416832 113082
rect 416780 113018 416832 113024
rect 416792 112713 416820 113018
rect 416778 112704 416834 112713
rect 416778 112639 416834 112648
rect 416780 111784 416832 111790
rect 416780 111726 416832 111732
rect 416792 110945 416820 111726
rect 416778 110936 416834 110945
rect 416778 110871 416834 110880
rect 417436 109313 417464 272478
rect 419448 271924 419500 271930
rect 419448 271866 419500 271872
rect 419264 186992 419316 186998
rect 419264 186934 419316 186940
rect 417514 177304 417570 177313
rect 417514 177239 417570 177248
rect 417528 121145 417556 177239
rect 419170 134600 419226 134609
rect 419170 134535 419226 134544
rect 417608 132456 417660 132462
rect 417608 132398 417660 132404
rect 417620 131345 417648 132398
rect 417606 131336 417662 131345
rect 417606 131271 417662 131280
rect 418528 126948 418580 126954
rect 418528 126890 418580 126896
rect 418540 126177 418568 126890
rect 418526 126168 418582 126177
rect 418526 126103 418582 126112
rect 418528 125588 418580 125594
rect 418528 125530 418580 125536
rect 418540 124545 418568 125530
rect 418526 124536 418582 124545
rect 418526 124471 418582 124480
rect 417514 121136 417570 121145
rect 417514 121071 417570 121080
rect 417422 109304 417478 109313
rect 417422 109239 417478 109248
rect 413284 107636 413336 107642
rect 413284 107578 413336 107584
rect 416780 107636 416832 107642
rect 416780 107578 416832 107584
rect 416792 107545 416820 107578
rect 416778 107536 416834 107545
rect 416778 107471 416834 107480
rect 416780 106276 416832 106282
rect 416780 106218 416832 106224
rect 416792 105913 416820 106218
rect 416778 105904 416834 105913
rect 416778 105839 416834 105848
rect 416780 104848 416832 104854
rect 416780 104790 416832 104796
rect 416792 104145 416820 104790
rect 416778 104136 416834 104145
rect 416778 104071 416834 104080
rect 416780 103488 416832 103494
rect 416780 103430 416832 103436
rect 416792 102513 416820 103430
rect 416778 102504 416834 102513
rect 416778 102439 416834 102448
rect 416780 102128 416832 102134
rect 416780 102070 416832 102076
rect 416792 100881 416820 102070
rect 416778 100872 416834 100881
rect 416778 100807 416834 100816
rect 411904 100020 411956 100026
rect 411904 99962 411956 99968
rect 396724 99204 396776 99210
rect 396724 99146 396776 99152
rect 392584 97912 392636 97918
rect 392584 97854 392636 97860
rect 414664 96960 414716 96966
rect 414664 96902 414716 96908
rect 385684 66156 385736 66162
rect 385684 66098 385736 66104
rect 414676 14482 414704 96902
rect 419184 95946 419212 134535
rect 419276 126954 419304 186934
rect 419356 133884 419408 133890
rect 419356 133826 419408 133832
rect 419368 132977 419396 133826
rect 419354 132968 419410 132977
rect 419354 132903 419410 132912
rect 419264 126948 419316 126954
rect 419264 126890 419316 126896
rect 419172 95940 419224 95946
rect 419172 95882 419224 95888
rect 419368 73166 419396 132903
rect 419460 125594 419488 271866
rect 419448 125588 419500 125594
rect 419448 125530 419500 125536
rect 419552 122806 419580 298726
rect 419632 191208 419684 191214
rect 419632 191150 419684 191156
rect 419644 128314 419672 191150
rect 420932 179466 420960 534686
rect 425072 190454 425100 538222
rect 429212 534750 429240 702782
rect 478524 702778 478552 703520
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 494808 702710 494836 703520
rect 453948 702704 454000 702710
rect 453948 702646 454000 702652
rect 492588 702704 492640 702710
rect 492588 702646 492640 702652
rect 494796 702704 494848 702710
rect 494796 702646 494848 702652
rect 453960 700330 453988 702646
rect 483664 701752 483716 701758
rect 483664 701694 483716 701700
rect 450544 700324 450596 700330
rect 450544 700266 450596 700272
rect 453948 700324 454000 700330
rect 453948 700266 454000 700272
rect 431224 575544 431276 575550
rect 431224 575486 431276 575492
rect 431236 565146 431264 575486
rect 431224 565140 431276 565146
rect 431224 565082 431276 565088
rect 429200 534744 429252 534750
rect 429200 534686 429252 534692
rect 431224 510672 431276 510678
rect 431224 510614 431276 510620
rect 430580 496800 430632 496806
rect 430580 496742 430632 496748
rect 430592 496262 430620 496742
rect 431236 496262 431264 510614
rect 430580 496256 430632 496262
rect 430580 496198 430632 496204
rect 431224 496256 431276 496262
rect 431224 496198 431276 496204
rect 427820 464364 427872 464370
rect 427820 464306 427872 464312
rect 425072 190426 425376 190454
rect 422944 185632 422996 185638
rect 422944 185574 422996 185580
rect 422956 179466 422984 185574
rect 425348 179466 425376 190426
rect 427832 179466 427860 464306
rect 430592 184890 430620 496198
rect 431960 457496 432012 457502
rect 431960 457438 432012 457444
rect 431972 190454 432000 457438
rect 441620 377460 441672 377466
rect 441620 377402 441672 377408
rect 436098 292632 436154 292641
rect 436098 292567 436154 292576
rect 434720 268388 434772 268394
rect 434720 268330 434772 268336
rect 431972 190426 432368 190454
rect 429936 184884 429988 184890
rect 429936 184826 429988 184832
rect 430580 184884 430632 184890
rect 430580 184826 430632 184832
rect 429948 179466 429976 184826
rect 432340 179466 432368 190426
rect 434732 179466 434760 268330
rect 436112 190454 436140 292567
rect 436112 190426 436968 190454
rect 436940 179466 436968 190426
rect 439412 181620 439464 181626
rect 439412 181562 439464 181568
rect 439424 179466 439452 181562
rect 441632 179466 441660 377402
rect 448520 282192 448572 282198
rect 448520 282134 448572 282140
rect 447784 271176 447836 271182
rect 447784 271118 447836 271124
rect 443000 246424 443052 246430
rect 443000 246366 443052 246372
rect 443012 190454 443040 246366
rect 445760 233980 445812 233986
rect 445760 233922 445812 233928
rect 445772 190454 445800 233922
rect 443012 190426 443960 190454
rect 445772 190426 446352 190454
rect 443932 179466 443960 190426
rect 446324 179466 446352 190426
rect 447796 181354 447824 271118
rect 447784 181348 447836 181354
rect 447784 181290 447836 181296
rect 448532 179466 448560 282134
rect 450556 185638 450584 700266
rect 464344 311160 464396 311166
rect 464344 311102 464396 311108
rect 452660 236700 452712 236706
rect 452660 236642 452712 236648
rect 452672 190454 452700 236642
rect 455418 232520 455474 232529
rect 455418 232455 455474 232464
rect 455432 190454 455460 232455
rect 462318 225584 462374 225593
rect 462318 225519 462374 225528
rect 457444 223644 457496 223650
rect 457444 223586 457496 223592
rect 452672 190426 453160 190454
rect 455432 190426 455552 190454
rect 450544 185632 450596 185638
rect 450544 185574 450596 185580
rect 451372 181348 451424 181354
rect 451372 181290 451424 181296
rect 451384 179466 451412 181290
rect 420932 179438 421130 179466
rect 422956 179438 423430 179466
rect 425348 179438 425730 179466
rect 427832 179438 428030 179466
rect 429948 179438 430422 179466
rect 432340 179438 432722 179466
rect 434732 179438 435022 179466
rect 436940 179438 437322 179466
rect 439424 179438 439714 179466
rect 441632 179438 442014 179466
rect 443932 179438 444314 179466
rect 446324 179438 446706 179466
rect 448532 179438 449006 179466
rect 451306 179438 451412 179466
rect 453132 179466 453160 190426
rect 455524 179466 455552 190426
rect 457456 182170 457484 223586
rect 459560 199504 459612 199510
rect 459560 199446 459612 199452
rect 459572 190454 459600 199446
rect 462332 190454 462360 225519
rect 459572 190426 460152 190454
rect 462332 190426 462544 190454
rect 457444 182164 457496 182170
rect 457444 182106 457496 182112
rect 458180 182164 458232 182170
rect 458180 182106 458232 182112
rect 458192 179466 458220 182106
rect 460124 179466 460152 190426
rect 462516 179466 462544 190426
rect 464356 184210 464384 311102
rect 475384 308440 475436 308446
rect 475384 308382 475436 308388
rect 467104 307828 467156 307834
rect 467104 307770 467156 307776
rect 466460 221468 466512 221474
rect 466460 221410 466512 221416
rect 465080 202156 465132 202162
rect 465080 202098 465132 202104
rect 464344 184204 464396 184210
rect 464344 184146 464396 184152
rect 465092 179466 465120 202098
rect 466472 180794 466500 221410
rect 467116 184346 467144 307770
rect 471244 262880 471296 262886
rect 471244 262822 471296 262828
rect 468484 229764 468536 229770
rect 468484 229706 468536 229712
rect 467104 184340 467156 184346
rect 467104 184282 467156 184288
rect 466472 180766 467144 180794
rect 467116 179466 467144 180766
rect 468496 180198 468524 229706
rect 469220 192500 469272 192506
rect 469220 192442 469272 192448
rect 469232 190454 469260 192442
rect 469232 190426 469536 190454
rect 468484 180192 468536 180198
rect 468484 180134 468536 180140
rect 469508 179466 469536 190426
rect 471256 181558 471284 262822
rect 472624 251864 472676 251870
rect 472624 251806 472676 251812
rect 471980 192636 472032 192642
rect 471980 192578 472032 192584
rect 471244 181552 471296 181558
rect 471244 181494 471296 181500
rect 471992 179466 472020 192578
rect 472636 184278 472664 251806
rect 473360 215960 473412 215966
rect 473360 215902 473412 215908
rect 473372 190454 473400 215902
rect 473372 190426 474136 190454
rect 472624 184272 472676 184278
rect 472624 184214 472676 184220
rect 474108 179466 474136 190426
rect 475396 182170 475424 308382
rect 482284 303680 482336 303686
rect 482284 303622 482336 303628
rect 478880 250504 478932 250510
rect 478880 250446 478932 250452
rect 475384 182164 475436 182170
rect 475384 182106 475436 182112
rect 476580 182164 476632 182170
rect 476580 182106 476632 182112
rect 476592 179466 476620 182106
rect 478892 179466 478920 250446
rect 480260 209092 480312 209098
rect 480260 209034 480312 209040
rect 480272 190454 480300 209034
rect 480272 190426 481128 190454
rect 481100 179466 481128 190426
rect 482296 181626 482324 303622
rect 483676 181694 483704 701694
rect 492600 700330 492628 702646
rect 527192 702642 527220 703520
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 511908 702568 511960 702574
rect 511908 702510 511960 702516
rect 511920 700330 511948 702510
rect 543476 702506 543504 703520
rect 559668 702574 559696 703520
rect 550548 702568 550600 702574
rect 550548 702510 550600 702516
rect 559656 702568 559708 702574
rect 559656 702510 559708 702516
rect 543464 702500 543516 702506
rect 543464 702442 543516 702448
rect 550560 700330 550588 702510
rect 492588 700324 492640 700330
rect 492588 700266 492640 700272
rect 511908 700324 511960 700330
rect 511908 700266 511960 700272
rect 550548 700324 550600 700330
rect 550548 700266 550600 700272
rect 511920 699718 511948 700266
rect 511264 699712 511316 699718
rect 511264 699654 511316 699660
rect 511908 699712 511960 699718
rect 511908 699654 511960 699660
rect 497464 565140 497516 565146
rect 497464 565082 497516 565088
rect 504364 565140 504416 565146
rect 504364 565082 504416 565088
rect 497476 464370 497504 565082
rect 504376 563718 504404 565082
rect 504364 563712 504416 563718
rect 504364 563654 504416 563660
rect 497464 464364 497516 464370
rect 497464 464306 497516 464312
rect 504364 352572 504416 352578
rect 504364 352514 504416 352520
rect 485044 341556 485096 341562
rect 485044 341498 485096 341504
rect 483664 181688 483716 181694
rect 483664 181630 483716 181636
rect 482284 181620 482336 181626
rect 482284 181562 482336 181568
rect 485056 181490 485084 341498
rect 499580 331900 499632 331906
rect 499580 331842 499632 331848
rect 495440 284368 495492 284374
rect 495440 284310 495492 284316
rect 493324 275324 493376 275330
rect 493324 275266 493376 275272
rect 489920 265668 489972 265674
rect 489920 265610 489972 265616
rect 485780 257372 485832 257378
rect 485780 257314 485832 257320
rect 483572 181484 483624 181490
rect 483572 181426 483624 181432
rect 485044 181484 485096 181490
rect 485044 181426 485096 181432
rect 483584 179466 483612 181426
rect 485792 179466 485820 257314
rect 489184 218816 489236 218822
rect 489184 218758 489236 218764
rect 488540 217320 488592 217326
rect 488540 217262 488592 217268
rect 488552 190454 488580 217262
rect 488552 190426 488672 190454
rect 488644 179466 488672 190426
rect 489196 181762 489224 218758
rect 489932 190454 489960 265610
rect 489932 190426 490512 190454
rect 489184 181756 489236 181762
rect 489184 181698 489236 181704
rect 453132 179438 453606 179466
rect 455524 179438 455998 179466
rect 458192 179438 458298 179466
rect 460124 179438 460598 179466
rect 462516 179438 462990 179466
rect 465092 179438 465290 179466
rect 467116 179438 467590 179466
rect 469508 179438 469890 179466
rect 471992 179438 472282 179466
rect 474108 179438 474582 179466
rect 476592 179438 476882 179466
rect 478892 179438 479274 179466
rect 481100 179438 481574 179466
rect 483584 179438 483874 179466
rect 485792 179438 486174 179466
rect 488566 179438 488672 179466
rect 490484 179466 490512 190426
rect 492864 181756 492916 181762
rect 492864 181698 492916 181704
rect 491300 180872 491352 180878
rect 491300 180814 491352 180820
rect 490484 179438 490866 179466
rect 491312 179353 491340 180814
rect 492876 179466 492904 181698
rect 493336 180266 493364 275266
rect 494244 247104 494296 247110
rect 494244 247046 494296 247052
rect 493324 180260 493376 180266
rect 493324 180202 493376 180208
rect 492876 179438 493166 179466
rect 491298 179344 491354 179353
rect 491298 179279 491354 179288
rect 494150 171048 494206 171057
rect 494150 170983 494206 170992
rect 419722 131336 419778 131345
rect 419722 131271 419778 131280
rect 419632 128308 419684 128314
rect 419632 128250 419684 128256
rect 419540 122800 419592 122806
rect 419538 122768 419540 122777
rect 419592 122768 419594 122777
rect 419538 122703 419594 122712
rect 419736 100706 419764 131271
rect 419816 128308 419868 128314
rect 419816 128250 419868 128256
rect 419828 127945 419856 128250
rect 419814 127936 419870 127945
rect 419814 127871 419870 127880
rect 419724 100700 419776 100706
rect 419724 100642 419776 100648
rect 494058 100056 494114 100065
rect 420564 96966 420592 100028
rect 420932 100014 421774 100042
rect 422312 100014 422970 100042
rect 423692 100014 424166 100042
rect 425072 100014 425362 100042
rect 420552 96960 420604 96966
rect 420552 96902 420604 96908
rect 420932 91050 420960 100014
rect 421012 97368 421064 97374
rect 421012 97310 421064 97316
rect 421024 96558 421052 97310
rect 421564 97300 421616 97306
rect 421564 97242 421616 97248
rect 421012 96552 421064 96558
rect 421012 96494 421064 96500
rect 420920 91044 420972 91050
rect 420920 90986 420972 90992
rect 419356 73160 419408 73166
rect 419356 73102 419408 73108
rect 414664 14476 414716 14482
rect 414664 14418 414716 14424
rect 421576 11014 421604 97242
rect 422312 73098 422340 100014
rect 422300 73092 422352 73098
rect 422300 73034 422352 73040
rect 421564 11008 421616 11014
rect 421564 10950 421616 10956
rect 374644 9648 374696 9654
rect 374644 9590 374696 9596
rect 423692 8974 423720 100014
rect 425072 33114 425100 100014
rect 426544 97374 426572 100028
rect 426532 97368 426584 97374
rect 426532 97310 426584 97316
rect 427740 94518 427768 100028
rect 427832 100014 428950 100042
rect 429212 100014 430146 100042
rect 430592 100014 431342 100042
rect 431972 100014 432538 100042
rect 433352 100014 433734 100042
rect 434732 100014 434930 100042
rect 436126 100014 436232 100042
rect 427728 94512 427780 94518
rect 427728 94454 427780 94460
rect 427832 44878 427860 100014
rect 427820 44872 427872 44878
rect 427820 44814 427872 44820
rect 429212 43518 429240 100014
rect 429200 43512 429252 43518
rect 429200 43454 429252 43460
rect 425060 33108 425112 33114
rect 425060 33050 425112 33056
rect 423680 8968 423732 8974
rect 373998 8936 374054 8945
rect 423680 8910 423732 8916
rect 373998 8871 374054 8880
rect 374012 4146 374040 8871
rect 430592 6798 430620 100014
rect 431972 7614 432000 100014
rect 433352 40730 433380 100014
rect 433340 40724 433392 40730
rect 433340 40666 433392 40672
rect 434732 39370 434760 100014
rect 434720 39364 434772 39370
rect 434720 39306 434772 39312
rect 436204 38010 436232 100014
rect 436296 100014 437322 100042
rect 437492 100014 438518 100042
rect 438872 100014 439714 100042
rect 436192 38004 436244 38010
rect 436192 37946 436244 37952
rect 436296 36650 436324 100014
rect 436284 36644 436336 36650
rect 436284 36586 436336 36592
rect 437492 35222 437520 100014
rect 437480 35216 437532 35222
rect 437480 35158 437532 35164
rect 438872 31142 438900 100014
rect 440896 96966 440924 100028
rect 441632 100014 442106 100042
rect 443012 100014 443302 100042
rect 444392 100014 444498 100042
rect 445786 100014 445892 100042
rect 439504 96960 439556 96966
rect 439504 96902 439556 96908
rect 440884 96960 440936 96966
rect 440884 96902 440936 96908
rect 438860 31136 438912 31142
rect 438860 31078 438912 31084
rect 431960 7608 432012 7614
rect 431960 7550 432012 7556
rect 439516 6866 439544 96902
rect 441632 30326 441660 100014
rect 441620 30320 441672 30326
rect 441620 30262 441672 30268
rect 443012 28286 443040 100014
rect 443000 28280 443052 28286
rect 443000 28222 443052 28228
rect 444392 26926 444420 100014
rect 444380 26920 444432 26926
rect 444380 26862 444432 26868
rect 445864 25702 445892 100014
rect 445956 100014 446982 100042
rect 447152 100014 448178 100042
rect 448532 100014 449374 100042
rect 449912 100014 450570 100042
rect 451292 100014 451766 100042
rect 452672 100014 452962 100042
rect 445852 25696 445904 25702
rect 445852 25638 445904 25644
rect 445956 24206 445984 100014
rect 445944 24200 445996 24206
rect 445944 24142 445996 24148
rect 447152 22846 447180 100014
rect 447140 22840 447192 22846
rect 447140 22782 447192 22788
rect 439504 6860 439556 6866
rect 439504 6802 439556 6808
rect 430580 6792 430632 6798
rect 430580 6734 430632 6740
rect 448532 5506 448560 100014
rect 449912 22098 449940 100014
rect 449900 22092 449952 22098
rect 449900 22034 449952 22040
rect 451292 20058 451320 100014
rect 451280 20052 451332 20058
rect 451280 19994 451332 20000
rect 452672 18698 452700 100014
rect 454040 96960 454092 96966
rect 454040 96902 454092 96908
rect 452660 18692 452712 18698
rect 452660 18634 452712 18640
rect 454052 15978 454080 96902
rect 454144 17270 454172 100028
rect 455064 100014 455354 100042
rect 455064 96966 455092 100014
rect 456536 97306 456564 100028
rect 456812 100014 457746 100042
rect 458192 100014 458942 100042
rect 456524 97300 456576 97306
rect 456524 97242 456576 97248
rect 455052 96960 455104 96966
rect 455052 96902 455104 96908
rect 456812 90370 456840 100014
rect 457444 96824 457496 96830
rect 457444 96766 457496 96772
rect 456800 90364 456852 90370
rect 456800 90306 456852 90312
rect 457456 86970 457484 96766
rect 458192 87650 458220 100014
rect 460124 96830 460152 100028
rect 460952 100014 461334 100042
rect 462332 100014 462530 100042
rect 463726 100014 463832 100042
rect 460112 96824 460164 96830
rect 460112 96766 460164 96772
rect 458180 87644 458232 87650
rect 458180 87586 458232 87592
rect 457444 86964 457496 86970
rect 457444 86906 457496 86912
rect 460952 84862 460980 100014
rect 461584 97300 461636 97306
rect 461584 97242 461636 97248
rect 460940 84856 460992 84862
rect 460940 84798 460992 84804
rect 461596 71194 461624 97242
rect 461584 71188 461636 71194
rect 461584 71130 461636 71136
rect 462332 43450 462360 100014
rect 463804 83502 463832 100014
rect 463896 100014 464922 100042
rect 465092 100014 466118 100042
rect 466472 100014 467314 100042
rect 467852 100014 468510 100042
rect 469232 100014 469706 100042
rect 470612 100014 470994 100042
rect 471992 100014 472190 100042
rect 463792 83496 463844 83502
rect 463792 83438 463844 83444
rect 463896 76566 463924 100014
rect 463884 76560 463936 76566
rect 463884 76502 463936 76508
rect 462320 43444 462372 43450
rect 462320 43386 462372 43392
rect 465092 42770 465120 100014
rect 466472 82142 466500 100014
rect 466460 82136 466512 82142
rect 466460 82078 466512 82084
rect 465080 42764 465132 42770
rect 465080 42706 465132 42712
rect 454132 17264 454184 17270
rect 454132 17206 454184 17212
rect 454040 15972 454092 15978
rect 454040 15914 454092 15920
rect 467852 13802 467880 100014
rect 469232 77994 469260 100014
rect 470612 80714 470640 100014
rect 470600 80708 470652 80714
rect 470600 80650 470652 80656
rect 471992 79354 472020 100014
rect 471980 79348 472032 79354
rect 471980 79290 472032 79296
rect 469220 77988 469272 77994
rect 469220 77930 469272 77936
rect 473372 75206 473400 100028
rect 474568 97306 474596 100028
rect 474752 100014 475778 100042
rect 476132 100014 476974 100042
rect 477512 100014 478170 100042
rect 478892 100014 479366 100042
rect 480272 100014 480562 100042
rect 474556 97300 474608 97306
rect 474556 97242 474608 97248
rect 473360 75200 473412 75206
rect 473360 75142 473412 75148
rect 474752 69766 474780 100014
rect 475384 97300 475436 97306
rect 475384 97242 475436 97248
rect 474740 69760 474792 69766
rect 474740 69702 474792 69708
rect 475396 54602 475424 97242
rect 476132 68406 476160 100014
rect 476120 68400 476172 68406
rect 476120 68342 476172 68348
rect 477512 67561 477540 100014
rect 477498 67552 477554 67561
rect 477498 67487 477554 67496
rect 475384 54596 475436 54602
rect 475384 54538 475436 54544
rect 467840 13796 467892 13802
rect 467840 13738 467892 13744
rect 478892 12442 478920 100014
rect 480272 66230 480300 100014
rect 481640 96960 481692 96966
rect 481640 96902 481692 96908
rect 480260 66224 480312 66230
rect 480260 66166 480312 66172
rect 481652 64870 481680 96902
rect 481744 91798 481772 100028
rect 482664 100014 482954 100042
rect 483032 100014 484150 100042
rect 484412 100014 485346 100042
rect 485792 100014 486542 100042
rect 482664 96966 482692 100014
rect 482652 96960 482704 96966
rect 482652 96902 482704 96908
rect 481732 91792 481784 91798
rect 481732 91734 481784 91740
rect 481640 64864 481692 64870
rect 481640 64806 481692 64812
rect 483032 62898 483060 100014
rect 483020 62892 483072 62898
rect 483020 62834 483072 62840
rect 484412 62082 484440 100014
rect 484400 62076 484452 62082
rect 484400 62018 484452 62024
rect 485792 60722 485820 100014
rect 487724 96966 487752 100028
rect 488552 100014 488934 100042
rect 489932 100014 490130 100042
rect 486424 96960 486476 96966
rect 486424 96902 486476 96908
rect 487712 96960 487764 96966
rect 487712 96902 487764 96908
rect 485780 60716 485832 60722
rect 485780 60658 485832 60664
rect 478880 12436 478932 12442
rect 478880 12378 478932 12384
rect 486436 10334 486464 96902
rect 488552 58750 488580 100014
rect 488540 58744 488592 58750
rect 488540 58686 488592 58692
rect 489932 57254 489960 100014
rect 489920 57248 489972 57254
rect 489920 57190 489972 57196
rect 491312 55962 491340 100028
rect 492508 97306 492536 100028
rect 492692 100014 493718 100042
rect 492496 97300 492548 97306
rect 492496 97242 492548 97248
rect 491300 55956 491352 55962
rect 491300 55898 491352 55904
rect 492692 53174 492720 100014
rect 494058 99991 494114 100000
rect 494072 99210 494100 99991
rect 494060 99204 494112 99210
rect 494060 99146 494112 99152
rect 492680 53168 492732 53174
rect 492680 53110 492732 53116
rect 494164 49706 494192 170983
rect 494256 132161 494284 247046
rect 494336 191140 494388 191146
rect 494336 191082 494388 191088
rect 494242 132152 494298 132161
rect 494242 132087 494298 132096
rect 494348 131073 494376 191082
rect 494426 171728 494482 171737
rect 494426 171663 494482 171672
rect 494334 131064 494390 131073
rect 494334 130999 494390 131008
rect 494152 49700 494204 49706
rect 494152 49642 494204 49648
rect 494440 46238 494468 171663
rect 495452 132977 495480 284310
rect 496820 278044 496872 278050
rect 496820 277986 496872 277992
rect 495624 180124 495676 180130
rect 495624 180066 495676 180072
rect 495530 168872 495586 168881
rect 495530 168807 495586 168816
rect 495438 132968 495494 132977
rect 495438 132903 495494 132912
rect 495438 104952 495494 104961
rect 495438 104887 495494 104896
rect 495452 102882 495480 104887
rect 495440 102876 495492 102882
rect 495440 102818 495492 102824
rect 495438 102776 495494 102785
rect 495438 102711 495494 102720
rect 495452 97986 495480 102711
rect 495440 97980 495492 97986
rect 495440 97922 495492 97928
rect 495544 52426 495572 168807
rect 495636 121825 495664 180066
rect 495714 147656 495770 147665
rect 495714 147591 495770 147600
rect 495622 121816 495678 121825
rect 495622 121751 495678 121760
rect 495624 102876 495676 102882
rect 495624 102818 495676 102824
rect 495636 96626 495664 102818
rect 495624 96620 495676 96626
rect 495624 96562 495676 96568
rect 495728 93809 495756 147591
rect 496832 141438 496860 277986
rect 498292 243568 498344 243574
rect 498292 243510 498344 243516
rect 496912 196648 496964 196654
rect 496912 196590 496964 196596
rect 496820 141432 496872 141438
rect 496820 141374 496872 141380
rect 496832 140865 496860 141374
rect 496818 140856 496874 140865
rect 496818 140791 496874 140800
rect 496820 140752 496872 140758
rect 496820 140694 496872 140700
rect 496832 139777 496860 140694
rect 496818 139768 496874 139777
rect 496818 139703 496874 139712
rect 496820 139392 496872 139398
rect 496820 139334 496872 139340
rect 496832 138689 496860 139334
rect 496818 138680 496874 138689
rect 496818 138615 496874 138624
rect 496820 137964 496872 137970
rect 496820 137906 496872 137912
rect 496832 137465 496860 137906
rect 496818 137456 496874 137465
rect 496818 137391 496874 137400
rect 496820 136604 496872 136610
rect 496820 136546 496872 136552
rect 496832 136377 496860 136546
rect 496818 136368 496874 136377
rect 496818 136303 496874 136312
rect 496820 135244 496872 135250
rect 496820 135186 496872 135192
rect 496832 134201 496860 135186
rect 496818 134192 496874 134201
rect 496818 134127 496874 134136
rect 496924 132494 496952 196590
rect 497002 177848 497058 177857
rect 497002 177783 497058 177792
rect 497016 177002 497044 177783
rect 497004 176996 497056 177002
rect 497004 176938 497056 176944
rect 497002 176760 497058 176769
rect 497002 176695 497004 176704
rect 497056 176695 497058 176704
rect 497004 176666 497056 176672
rect 498106 175672 498162 175681
rect 498162 175630 498240 175658
rect 498106 175607 498162 175616
rect 497002 174448 497058 174457
rect 497002 174383 497058 174392
rect 497016 174282 497044 174383
rect 497004 174276 497056 174282
rect 497004 174218 497056 174224
rect 497004 170808 497056 170814
rect 497004 170750 497056 170756
rect 497016 169969 497044 170750
rect 497002 169960 497058 169969
rect 497002 169895 497058 169904
rect 497004 168360 497056 168366
rect 497004 168302 497056 168308
rect 497016 167793 497044 168302
rect 497002 167784 497058 167793
rect 497002 167719 497058 167728
rect 497004 167000 497056 167006
rect 497004 166942 497056 166948
rect 497016 166705 497044 166942
rect 497002 166696 497058 166705
rect 497002 166631 497058 166640
rect 497096 165572 497148 165578
rect 497096 165514 497148 165520
rect 497002 165472 497058 165481
rect 497002 165407 497058 165416
rect 497016 164898 497044 165407
rect 497004 164892 497056 164898
rect 497004 164834 497056 164840
rect 497108 164393 497136 165514
rect 497094 164384 497150 164393
rect 497094 164319 497150 164328
rect 497004 164212 497056 164218
rect 497004 164154 497056 164160
rect 497016 163305 497044 164154
rect 497002 163296 497058 163305
rect 497002 163231 497058 163240
rect 497004 162852 497056 162858
rect 497004 162794 497056 162800
rect 497016 162217 497044 162794
rect 497002 162208 497058 162217
rect 497002 162143 497058 162152
rect 497004 161424 497056 161430
rect 497004 161366 497056 161372
rect 497016 160993 497044 161366
rect 497002 160984 497058 160993
rect 497002 160919 497058 160928
rect 497004 160064 497056 160070
rect 497004 160006 497056 160012
rect 497016 159905 497044 160006
rect 497096 159996 497148 160002
rect 497096 159938 497148 159944
rect 497002 159896 497058 159905
rect 497002 159831 497058 159840
rect 497108 158817 497136 159938
rect 497094 158808 497150 158817
rect 497094 158743 497150 158752
rect 497004 158704 497056 158710
rect 497004 158646 497056 158652
rect 497016 157729 497044 158646
rect 497002 157720 497058 157729
rect 497002 157655 497058 157664
rect 497004 157344 497056 157350
rect 497004 157286 497056 157292
rect 497016 156505 497044 157286
rect 497002 156496 497058 156505
rect 497002 156431 497058 156440
rect 497004 155916 497056 155922
rect 497004 155858 497056 155864
rect 497016 155417 497044 155858
rect 497002 155408 497058 155417
rect 497002 155343 497058 155352
rect 497004 154556 497056 154562
rect 497004 154498 497056 154504
rect 497016 154329 497044 154498
rect 497096 154488 497148 154494
rect 497096 154430 497148 154436
rect 497002 154320 497058 154329
rect 497002 154255 497058 154264
rect 497108 153241 497136 154430
rect 497094 153232 497150 153241
rect 497004 153196 497056 153202
rect 497094 153167 497150 153176
rect 497004 153138 497056 153144
rect 497016 152153 497044 153138
rect 497002 152144 497058 152153
rect 497002 152079 497058 152088
rect 497004 151768 497056 151774
rect 497004 151710 497056 151716
rect 497016 150929 497044 151710
rect 497002 150920 497058 150929
rect 497002 150855 497058 150864
rect 497004 150408 497056 150414
rect 497004 150350 497056 150356
rect 497016 149841 497044 150350
rect 497002 149832 497058 149841
rect 497002 149767 497058 149776
rect 497004 149048 497056 149054
rect 497004 148990 497056 148996
rect 497016 148753 497044 148990
rect 497002 148744 497058 148753
rect 497002 148679 497058 148688
rect 497004 147620 497056 147626
rect 497004 147562 497056 147568
rect 497016 146441 497044 147562
rect 497002 146432 497058 146441
rect 497002 146367 497058 146376
rect 497002 145344 497058 145353
rect 497002 145279 497058 145288
rect 497016 144974 497044 145279
rect 497004 144968 497056 144974
rect 497004 144910 497056 144916
rect 497094 144256 497150 144265
rect 497094 144191 497150 144200
rect 497108 143614 497136 144191
rect 497096 143608 497148 143614
rect 497096 143550 497148 143556
rect 497004 143540 497056 143546
rect 497004 143482 497056 143488
rect 497016 143177 497044 143482
rect 497002 143168 497058 143177
rect 497002 143103 497058 143112
rect 497004 142112 497056 142118
rect 497004 142054 497056 142060
rect 497016 141953 497044 142054
rect 497002 141944 497058 141953
rect 497002 141879 497058 141888
rect 497004 136536 497056 136542
rect 497004 136478 497056 136484
rect 497016 135289 497044 136478
rect 497002 135280 497058 135289
rect 497002 135215 497058 135224
rect 496924 132466 497044 132494
rect 496820 129736 496872 129742
rect 496818 129704 496820 129713
rect 496872 129704 496874 129713
rect 496818 129639 496874 129648
rect 496912 129668 496964 129674
rect 496912 129610 496964 129616
rect 496924 128489 496952 129610
rect 496910 128480 496966 128489
rect 496910 128415 496966 128424
rect 496912 127016 496964 127022
rect 496912 126958 496964 126964
rect 496820 126948 496872 126954
rect 496820 126890 496872 126896
rect 496832 126313 496860 126890
rect 496818 126304 496874 126313
rect 496818 126239 496874 126248
rect 496820 125588 496872 125594
rect 496820 125530 496872 125536
rect 496832 125225 496860 125530
rect 496818 125216 496874 125225
rect 496818 125151 496874 125160
rect 496820 124160 496872 124166
rect 496818 124128 496820 124137
rect 496872 124128 496874 124137
rect 496818 124063 496874 124072
rect 496924 122913 496952 126958
rect 496910 122904 496966 122913
rect 496910 122839 496966 122848
rect 496820 121440 496872 121446
rect 496820 121382 496872 121388
rect 496832 120737 496860 121382
rect 496818 120728 496874 120737
rect 496818 120663 496874 120672
rect 496820 119808 496872 119814
rect 496820 119750 496872 119756
rect 496832 119649 496860 119750
rect 496818 119640 496874 119649
rect 496818 119575 496874 119584
rect 496820 118652 496872 118658
rect 496820 118594 496872 118600
rect 496832 118425 496860 118594
rect 496912 118584 496964 118590
rect 496912 118526 496964 118532
rect 496818 118416 496874 118425
rect 496818 118351 496874 118360
rect 496924 117337 496952 118526
rect 496910 117328 496966 117337
rect 496910 117263 496966 117272
rect 497016 116249 497044 132466
rect 497002 116240 497058 116249
rect 497002 116175 497058 116184
rect 496820 115932 496872 115938
rect 496820 115874 496872 115880
rect 496832 115161 496860 115874
rect 496818 115152 496874 115161
rect 496818 115087 496874 115096
rect 496820 114504 496872 114510
rect 496820 114446 496872 114452
rect 496832 113937 496860 114446
rect 496818 113928 496874 113937
rect 496818 113863 496874 113872
rect 496820 113144 496872 113150
rect 496820 113086 496872 113092
rect 496832 112849 496860 113086
rect 496818 112840 496874 112849
rect 496818 112775 496874 112784
rect 496912 111784 496964 111790
rect 496818 111752 496874 111761
rect 496912 111726 496964 111732
rect 496818 111687 496820 111696
rect 496872 111687 496874 111696
rect 496820 111658 496872 111664
rect 496924 110673 496952 111726
rect 496910 110664 496966 110673
rect 496910 110599 496966 110608
rect 496820 110424 496872 110430
rect 496820 110366 496872 110372
rect 496832 109449 496860 110366
rect 496818 109440 496874 109449
rect 496818 109375 496874 109384
rect 497002 108352 497058 108361
rect 497002 108287 497058 108296
rect 496818 106176 496874 106185
rect 496818 106111 496874 106120
rect 496832 100638 496860 106111
rect 496910 103864 496966 103873
rect 496910 103799 496966 103808
rect 496820 100632 496872 100638
rect 496820 100574 496872 100580
rect 496924 97918 496952 103799
rect 497016 99278 497044 108287
rect 497094 107264 497150 107273
rect 497094 107199 497150 107208
rect 497108 99346 497136 107199
rect 497096 99340 497148 99346
rect 497096 99282 497148 99288
rect 497004 99272 497056 99278
rect 497004 99214 497056 99220
rect 496912 97912 496964 97918
rect 496912 97854 496964 97860
rect 495714 93800 495770 93809
rect 495714 93735 495770 93744
rect 495532 52420 495584 52426
rect 495532 52362 495584 52368
rect 498212 48278 498240 175630
rect 498304 127022 498332 243510
rect 498384 206304 498436 206310
rect 498384 206246 498436 206252
rect 498292 127016 498344 127022
rect 498292 126958 498344 126964
rect 498396 101697 498424 206246
rect 498476 176996 498528 177002
rect 498476 176938 498528 176944
rect 498382 101688 498438 101697
rect 498382 101623 498438 101632
rect 498488 95198 498516 176938
rect 499592 124166 499620 331842
rect 499672 246356 499724 246362
rect 499672 246298 499724 246304
rect 499580 124160 499632 124166
rect 499580 124102 499632 124108
rect 499684 114510 499712 246298
rect 502340 233912 502392 233918
rect 502340 233854 502392 233860
rect 501052 214668 501104 214674
rect 501052 214610 501104 214616
rect 499764 184340 499816 184346
rect 499764 184282 499816 184288
rect 499776 119814 499804 184282
rect 499856 183592 499908 183598
rect 499856 183534 499908 183540
rect 499868 170814 499896 183534
rect 500960 176724 501012 176730
rect 500960 176666 501012 176672
rect 499856 170808 499908 170814
rect 499856 170750 499908 170756
rect 499764 119808 499816 119814
rect 499764 119750 499816 119756
rect 499672 114504 499724 114510
rect 499672 114446 499724 114452
rect 498476 95192 498528 95198
rect 498476 95134 498528 95140
rect 498200 48272 498252 48278
rect 498200 48214 498252 48220
rect 494428 46232 494480 46238
rect 494428 46174 494480 46180
rect 486424 10328 486476 10334
rect 486424 10270 486476 10276
rect 448520 5500 448572 5506
rect 448520 5442 448572 5448
rect 374000 4140 374052 4146
rect 374000 4082 374052 4088
rect 360844 3528 360896 3534
rect 360844 3470 360896 3476
rect 500972 3466 501000 176666
rect 501064 113150 501092 214610
rect 501236 203584 501288 203590
rect 501236 203526 501288 203532
rect 501144 174276 501196 174282
rect 501144 174218 501196 174224
rect 501052 113144 501104 113150
rect 501052 113086 501104 113092
rect 501156 89690 501184 174218
rect 501248 150414 501276 203526
rect 502352 168366 502380 233854
rect 503720 218748 503772 218754
rect 503720 218690 503772 218696
rect 502524 182844 502576 182850
rect 502524 182786 502576 182792
rect 502432 181688 502484 181694
rect 502432 181630 502484 181636
rect 502340 168360 502392 168366
rect 502340 168302 502392 168308
rect 501236 150408 501288 150414
rect 501236 150350 501288 150356
rect 502340 144968 502392 144974
rect 502340 144910 502392 144916
rect 501144 89684 501196 89690
rect 501144 89626 501196 89632
rect 502352 74526 502380 144910
rect 502444 111722 502472 181630
rect 502536 154562 502564 182786
rect 502616 181620 502668 181626
rect 502616 181562 502668 181568
rect 502524 154556 502576 154562
rect 502524 154498 502576 154504
rect 502628 154494 502656 181562
rect 503628 168360 503680 168366
rect 503628 168302 503680 168308
rect 503640 167686 503668 168302
rect 503628 167680 503680 167686
rect 503628 167622 503680 167628
rect 502616 154488 502668 154494
rect 502616 154430 502668 154436
rect 502984 145580 503036 145586
rect 502984 145522 503036 145528
rect 502996 140758 503024 145522
rect 503260 141432 503312 141438
rect 503260 141374 503312 141380
rect 502984 140752 503036 140758
rect 502984 140694 503036 140700
rect 503272 140078 503300 141374
rect 503260 140072 503312 140078
rect 503260 140014 503312 140020
rect 503732 115938 503760 218690
rect 503810 188320 503866 188329
rect 503810 188255 503866 188264
rect 503720 115932 503772 115938
rect 503720 115874 503772 115880
rect 503824 111790 503852 188255
rect 503904 180192 503956 180198
rect 503904 180134 503956 180140
rect 503916 164898 503944 180134
rect 503904 164892 503956 164898
rect 503904 164834 503956 164840
rect 503916 164490 503944 164834
rect 503904 164484 503956 164490
rect 503904 164426 503956 164432
rect 504376 160002 504404 352514
rect 506480 338768 506532 338774
rect 506480 338710 506532 338716
rect 505284 189780 505336 189786
rect 505284 189722 505336 189728
rect 505192 181484 505244 181490
rect 505192 181426 505244 181432
rect 505100 178696 505152 178702
rect 505100 178638 505152 178644
rect 504456 164484 504508 164490
rect 504456 164426 504508 164432
rect 504364 159996 504416 160002
rect 504364 159938 504416 159944
rect 503812 111784 503864 111790
rect 503812 111726 503864 111732
rect 502432 111716 502484 111722
rect 502432 111658 502484 111664
rect 504468 86970 504496 164426
rect 505112 147626 505140 178638
rect 505204 153202 505232 181426
rect 505296 167006 505324 189722
rect 505284 167000 505336 167006
rect 505284 166942 505336 166948
rect 505296 166326 505324 166942
rect 505284 166320 505336 166326
rect 505284 166262 505336 166268
rect 505192 153196 505244 153202
rect 505192 153138 505244 153144
rect 505100 147620 505152 147626
rect 505100 147562 505152 147568
rect 506492 136542 506520 338710
rect 507860 287700 507912 287706
rect 507860 287642 507912 287648
rect 506572 195288 506624 195294
rect 506572 195230 506624 195236
rect 506480 136536 506532 136542
rect 506480 136478 506532 136484
rect 506584 110430 506612 195230
rect 506664 184272 506716 184278
rect 506664 184214 506716 184220
rect 506676 129674 506704 184214
rect 507872 165578 507900 287642
rect 508504 254584 508556 254590
rect 508504 254526 508556 254532
rect 508516 206310 508544 254526
rect 508504 206304 508556 206310
rect 508504 206246 508556 206252
rect 508044 181552 508096 181558
rect 508044 181494 508096 181500
rect 507952 180260 508004 180266
rect 507952 180202 508004 180208
rect 507860 165572 507912 165578
rect 507860 165514 507912 165520
rect 507872 164898 507900 165514
rect 507860 164892 507912 164898
rect 507860 164834 507912 164840
rect 507964 142118 507992 180202
rect 508056 151774 508084 181494
rect 508516 162858 508544 206246
rect 509240 199436 509292 199442
rect 509240 199378 509292 199384
rect 508504 162852 508556 162858
rect 508504 162794 508556 162800
rect 508044 151768 508096 151774
rect 508044 151710 508096 151716
rect 508044 144220 508096 144226
rect 508044 144162 508096 144168
rect 509148 144220 509200 144226
rect 509148 144162 509200 144168
rect 508056 143614 508084 144162
rect 508044 143608 508096 143614
rect 508044 143550 508096 143556
rect 507952 142112 508004 142118
rect 507952 142054 508004 142060
rect 507964 140826 507992 142054
rect 507952 140820 508004 140826
rect 507952 140762 508004 140768
rect 506664 129668 506716 129674
rect 506664 129610 506716 129616
rect 506572 110424 506624 110430
rect 506572 110366 506624 110372
rect 504456 86964 504508 86970
rect 504456 86906 504508 86912
rect 502340 74520 502392 74526
rect 502340 74462 502392 74468
rect 509160 20670 509188 144162
rect 509252 118590 509280 199378
rect 510620 198008 510672 198014
rect 510620 197950 510672 197956
rect 509332 193248 509384 193254
rect 509332 193190 509384 193196
rect 509344 149054 509372 193190
rect 509332 149048 509384 149054
rect 509332 148990 509384 148996
rect 510632 129742 510660 197950
rect 511276 155922 511304 699654
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580908 670744 580960 670750
rect 580906 670712 580908 670721
rect 580960 670712 580962 670721
rect 580906 670647 580962 670656
rect 582378 670712 582434 670721
rect 582378 670647 582434 670656
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616146 580212 617471
rect 580172 616140 580224 616146
rect 580172 616082 580224 616088
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 556804 590708 556856 590714
rect 556804 590650 556856 590656
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 556816 554062 556844 590650
rect 580170 582448 580226 582457
rect 580170 582383 580226 582392
rect 580184 577697 580212 582383
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563718 580212 564295
rect 580172 563712 580224 563718
rect 580172 563654 580224 563660
rect 556804 554056 556856 554062
rect 556804 553998 556856 554004
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 579804 525768 579856 525774
rect 579804 525710 579856 525716
rect 579816 524521 579844 525710
rect 579802 524512 579858 524521
rect 579802 524447 579858 524456
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580354 490512 580410 490521
rect 580354 490447 580410 490456
rect 579620 489184 579672 489190
rect 579620 489126 579672 489132
rect 579632 458153 579660 489126
rect 580368 484673 580396 490447
rect 580354 484664 580410 484673
rect 580354 484599 580410 484608
rect 579894 471472 579950 471481
rect 579894 471407 579950 471416
rect 579908 470626 579936 471407
rect 579896 470620 579948 470626
rect 579896 470562 579948 470568
rect 579618 458144 579674 458153
rect 579618 458079 579674 458088
rect 579632 457502 579660 458079
rect 579620 457496 579672 457502
rect 579620 457438 579672 457444
rect 579804 431928 579856 431934
rect 579804 431870 579856 431876
rect 579816 431633 579844 431870
rect 579802 431624 579858 431633
rect 579802 431559 579858 431568
rect 579620 428460 579672 428466
rect 579620 428402 579672 428408
rect 579632 418810 579660 428402
rect 525064 418804 525116 418810
rect 525064 418746 525116 418752
rect 579620 418804 579672 418810
rect 579620 418746 579672 418752
rect 579988 418804 580040 418810
rect 579988 418746 580040 418752
rect 519544 378820 519596 378826
rect 519544 378762 519596 378768
rect 514760 306400 514812 306406
rect 514760 306342 514812 306348
rect 512000 294704 512052 294710
rect 512000 294646 512052 294652
rect 512012 289134 512040 294646
rect 512000 289128 512052 289134
rect 512000 289070 512052 289076
rect 512012 160070 512040 289070
rect 513380 228404 513432 228410
rect 513380 228346 513432 228352
rect 512092 213240 512144 213246
rect 512092 213182 512144 213188
rect 512000 160064 512052 160070
rect 512000 160006 512052 160012
rect 511264 155916 511316 155922
rect 511264 155858 511316 155864
rect 512104 144226 512132 213182
rect 512184 184204 512236 184210
rect 512184 184146 512236 184152
rect 512092 144220 512144 144226
rect 512092 144162 512144 144168
rect 511264 140820 511316 140826
rect 511264 140762 511316 140768
rect 510620 129736 510672 129742
rect 510620 129678 510672 129684
rect 509240 118584 509292 118590
rect 509240 118526 509292 118532
rect 511276 101454 511304 140762
rect 512196 118658 512224 184146
rect 513392 143546 513420 228346
rect 513380 143540 513432 143546
rect 513380 143482 513432 143488
rect 513392 143410 513420 143482
rect 513380 143404 513432 143410
rect 513380 143346 513432 143352
rect 514772 126954 514800 306342
rect 517612 260160 517664 260166
rect 517612 260102 517664 260108
rect 517520 249076 517572 249082
rect 517520 249018 517572 249024
rect 515404 232552 515456 232558
rect 515404 232494 515456 232500
rect 515416 161430 515444 232494
rect 515404 161424 515456 161430
rect 515404 161366 515456 161372
rect 515404 143404 515456 143410
rect 515404 143346 515456 143352
rect 514760 126948 514812 126954
rect 514760 126890 514812 126896
rect 512184 118652 512236 118658
rect 512184 118594 512236 118600
rect 511264 101448 511316 101454
rect 511264 101390 511316 101396
rect 515416 60722 515444 143346
rect 517532 121446 517560 249018
rect 517624 164218 517652 260102
rect 517612 164212 517664 164218
rect 517612 164154 517664 164160
rect 519556 158710 519584 378762
rect 521660 309800 521712 309806
rect 521660 309742 521712 309748
rect 520924 256012 520976 256018
rect 520924 255954 520976 255960
rect 520936 218754 520964 255954
rect 520924 218748 520976 218754
rect 520924 218690 520976 218696
rect 519544 158704 519596 158710
rect 519544 158646 519596 158652
rect 520936 139398 520964 218690
rect 520924 139392 520976 139398
rect 520924 139334 520976 139340
rect 521672 125594 521700 309742
rect 525076 135250 525104 418746
rect 580000 418305 580028 418746
rect 579986 418296 580042 418305
rect 579986 418231 580042 418240
rect 579618 404968 579674 404977
rect 579618 404903 579674 404912
rect 579632 404394 579660 404903
rect 579620 404388 579672 404394
rect 579620 404330 579672 404336
rect 579632 378826 579660 404330
rect 579620 378820 579672 378826
rect 579620 378762 579672 378768
rect 580354 378448 580410 378457
rect 580354 378383 580410 378392
rect 579620 366376 579672 366382
rect 579620 366318 579672 366324
rect 579632 352578 579660 366318
rect 580262 365120 580318 365129
rect 580262 365055 580318 365064
rect 579620 352572 579672 352578
rect 579620 352514 579672 352520
rect 579632 351937 579660 352514
rect 579618 351928 579674 351937
rect 579618 351863 579674 351872
rect 580276 338774 580304 365055
rect 580368 354006 580396 378383
rect 580356 354000 580408 354006
rect 580356 353942 580408 353948
rect 580264 338768 580316 338774
rect 580264 338710 580316 338716
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311166 580212 312015
rect 539508 311160 539560 311166
rect 539508 311102 539560 311108
rect 580172 311160 580224 311166
rect 580172 311102 580224 311108
rect 539520 310554 539548 311102
rect 538220 310548 538272 310554
rect 538220 310490 538272 310496
rect 539508 310548 539560 310554
rect 539508 310490 539560 310496
rect 525800 294636 525852 294642
rect 525800 294578 525852 294584
rect 525812 146266 525840 294578
rect 536104 164892 536156 164898
rect 536104 164834 536156 164840
rect 525800 146260 525852 146266
rect 525800 146202 525852 146208
rect 525812 145586 525840 146202
rect 525800 145580 525852 145586
rect 525800 145522 525852 145528
rect 525064 135244 525116 135250
rect 525064 135186 525116 135192
rect 536116 127634 536144 164834
rect 538232 136610 538260 310490
rect 580276 298790 580304 325207
rect 580264 298784 580316 298790
rect 580264 298726 580316 298732
rect 580906 298752 580962 298761
rect 580906 298687 580962 298696
rect 580920 294710 580948 298687
rect 580908 294704 580960 294710
rect 580908 294646 580960 294652
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 547880 258732 547932 258738
rect 547880 258674 547932 258680
rect 547892 258126 547920 258674
rect 580184 258126 580212 258839
rect 547880 258120 547932 258126
rect 547880 258062 547932 258068
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 543004 167680 543056 167686
rect 543004 167622 543056 167628
rect 538220 136604 538272 136610
rect 538220 136546 538272 136552
rect 536104 127628 536156 127634
rect 536104 127570 536156 127576
rect 521660 125588 521712 125594
rect 521660 125530 521712 125536
rect 517520 121440 517572 121446
rect 517520 121382 517572 121388
rect 515404 60716 515456 60722
rect 515404 60658 515456 60664
rect 509148 20664 509200 20670
rect 509148 20606 509200 20612
rect 543016 6866 543044 167622
rect 544384 166320 544436 166326
rect 544384 166262 544436 166268
rect 544396 46918 544424 166262
rect 546500 165640 546552 165646
rect 546500 165582 546552 165588
rect 546512 164218 546540 165582
rect 546500 164212 546552 164218
rect 546500 164154 546552 164160
rect 547892 137970 547920 258062
rect 579986 245576 580042 245585
rect 579986 245511 580042 245520
rect 580000 244322 580028 245511
rect 579620 244316 579672 244322
rect 579620 244258 579672 244264
rect 579988 244316 580040 244322
rect 579988 244258 580040 244264
rect 579632 232558 579660 244258
rect 579620 232552 579672 232558
rect 579620 232494 579672 232500
rect 580262 232384 580318 232393
rect 580262 232319 580318 232328
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580184 218754 580212 218991
rect 580172 218748 580224 218754
rect 580172 218690 580224 218696
rect 580172 206304 580224 206310
rect 580172 206246 580224 206252
rect 580184 205737 580212 206246
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580184 191214 580212 192471
rect 580172 191208 580224 191214
rect 580172 191150 580224 191156
rect 580276 186998 580304 232319
rect 580264 186992 580316 186998
rect 580264 186934 580316 186940
rect 574744 179444 574796 179450
rect 574744 179386 574796 179392
rect 574756 153202 574784 179386
rect 580262 179208 580318 179217
rect 580262 179143 580318 179152
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 574744 153196 574796 153202
rect 574744 153138 574796 153144
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 580276 146266 580304 179143
rect 582392 157350 582420 670647
rect 582380 157344 582432 157350
rect 582380 157286 582432 157292
rect 580264 146260 580316 146266
rect 580264 146202 580316 146208
rect 580172 140072 580224 140078
rect 580172 140014 580224 140020
rect 580184 139369 580212 140014
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 547880 137964 547932 137970
rect 547880 137906 547932 137912
rect 580172 127628 580224 127634
rect 580172 127570 580224 127576
rect 580184 126041 580212 127570
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580262 112840 580318 112849
rect 580262 112775 580318 112784
rect 580172 101448 580224 101454
rect 580172 101390 580224 101396
rect 580184 99521 580212 101390
rect 580276 100706 580304 112775
rect 580264 100700 580316 100706
rect 580264 100642 580316 100648
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580264 95940 580316 95946
rect 580264 95882 580316 95888
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 544384 46912 544436 46918
rect 544384 46854 544436 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580276 33153 580304 95882
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 543004 6860 543056 6866
rect 543004 6802 543056 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 500960 3460 501012 3466
rect 500960 3402 501012 3408
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3514 658144 3570 658200
rect 3514 632068 3516 632088
rect 3516 632068 3568 632088
rect 3568 632068 3570 632088
rect 3514 632032 3570 632068
rect 3514 619112 3570 619168
rect 3514 606056 3570 606112
rect 3422 579944 3478 580000
rect 3238 566888 3294 566944
rect 3514 553832 3570 553888
rect 3146 527856 3202 527912
rect 2778 514820 2834 514856
rect 2778 514800 2780 514820
rect 2780 514800 2832 514820
rect 2832 514800 2834 514820
rect 3422 501744 3478 501800
rect 3422 475632 3478 475688
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3146 449520 3202 449576
rect 3514 423544 3570 423600
rect 3422 410488 3478 410544
rect 3146 397432 3202 397488
rect 3238 371320 3294 371376
rect 3146 358400 3202 358456
rect 2778 345344 2834 345400
rect 3422 319232 3478 319288
rect 33782 360032 33838 360088
rect 33046 347656 33102 347712
rect 3422 306212 3424 306232
rect 3424 306212 3476 306232
rect 3476 306212 3478 306232
rect 3422 306176 3478 306212
rect 3054 293120 3110 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 3146 241032 3202 241088
rect 3422 214920 3478 214976
rect 3238 201864 3294 201920
rect 1306 181328 1362 181384
rect 3514 188844 3516 188864
rect 3516 188844 3568 188864
rect 3568 188844 3570 188864
rect 3514 188808 3570 188844
rect 3422 162832 3478 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3698 110608 3754 110664
rect 2778 97552 2834 97608
rect 4066 93744 4122 93800
rect 3146 84632 3202 84688
rect 12438 76472 12494 76528
rect 3422 71612 3424 71632
rect 3424 71612 3476 71632
rect 3476 71612 3478 71632
rect 3422 71576 3478 71612
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 2870 28192 2926 28248
rect 3422 19352 3478 19408
rect 9678 26832 9734 26888
rect 3422 6432 3478 6488
rect 31758 46144 31814 46200
rect 38566 525816 38622 525872
rect 39946 77152 40002 77208
rect 42706 433200 42762 433256
rect 42614 302096 42670 302152
rect 45374 357448 45430 357504
rect 50710 492632 50766 492688
rect 49606 474680 49662 474736
rect 49606 380160 49662 380216
rect 54942 583752 54998 583808
rect 50894 387640 50950 387696
rect 54114 493348 54116 493368
rect 54116 493348 54168 493368
rect 54168 493348 54170 493368
rect 54114 493312 54170 493348
rect 54942 480256 54998 480312
rect 53746 377712 53802 377768
rect 55954 474680 56010 474736
rect 55034 339632 55090 339688
rect 55034 332036 55090 332072
rect 55034 332016 55036 332036
rect 55036 332016 55088 332036
rect 55088 332016 55090 332036
rect 56322 370504 56378 370560
rect 57242 390496 57298 390552
rect 57242 292848 57298 292904
rect 49698 57160 49754 57216
rect 58070 481480 58126 481536
rect 59174 481480 59230 481536
rect 59174 480256 59230 480312
rect 58530 388320 58586 388376
rect 59082 377984 59138 378040
rect 57886 347656 57942 347712
rect 58990 338000 59046 338056
rect 63222 477436 63224 477456
rect 63224 477436 63276 477456
rect 63276 477436 63278 477456
rect 63222 477400 63278 477436
rect 60554 236544 60610 236600
rect 59266 93608 59322 93664
rect 63314 448568 63370 448624
rect 64510 480120 64566 480176
rect 65982 490456 66038 490512
rect 64970 477536 65026 477592
rect 64142 368328 64198 368384
rect 64786 380160 64842 380216
rect 64786 378120 64842 378176
rect 63314 330520 63370 330576
rect 67638 581304 67694 581360
rect 67730 579128 67786 579184
rect 67638 578448 67694 578504
rect 67638 577768 67694 577824
rect 67546 577088 67602 577144
rect 67454 572736 67510 572792
rect 66074 470464 66130 470520
rect 67362 564440 67418 564496
rect 65890 383832 65946 383888
rect 65890 373940 65892 373960
rect 65892 373940 65944 373960
rect 65944 373940 65946 373960
rect 65890 373904 65946 373940
rect 67638 575728 67694 575784
rect 67730 575048 67786 575104
rect 67638 574368 67694 574424
rect 67638 573416 67694 573472
rect 68650 580624 68706 580680
rect 68650 576408 68706 576464
rect 68282 571648 68338 571704
rect 68466 571648 68522 571704
rect 67638 570016 67694 570072
rect 67638 568656 67694 568712
rect 67730 567568 67786 567624
rect 67638 567160 67694 567216
rect 67638 566208 67694 566264
rect 67638 564848 67694 564904
rect 67730 563488 67786 563544
rect 67638 563116 67640 563136
rect 67640 563116 67692 563136
rect 67692 563116 67694 563136
rect 67638 563080 67694 563116
rect 67638 562300 67640 562320
rect 67640 562300 67692 562320
rect 67692 562300 67694 562320
rect 67638 562264 67694 562300
rect 67638 562128 67694 562184
rect 67730 560768 67786 560824
rect 67638 560360 67694 560416
rect 67638 559408 67694 559464
rect 67638 557540 67640 557560
rect 67640 557540 67692 557560
rect 67692 557540 67694 557560
rect 67638 557504 67694 557540
rect 68282 557368 68338 557424
rect 67730 556688 67786 556744
rect 67638 556144 67694 556200
rect 67730 555328 67786 555384
rect 67638 554820 67640 554840
rect 67640 554820 67692 554840
rect 67692 554820 67694 554840
rect 67638 554784 67694 554820
rect 67638 553444 67694 553480
rect 67638 553424 67640 553444
rect 67640 553424 67692 553444
rect 67692 553424 67694 553444
rect 67638 552084 67694 552120
rect 67638 552064 67640 552084
rect 67640 552064 67692 552084
rect 67692 552064 67694 552084
rect 67638 551248 67694 551304
rect 67638 549888 67694 549944
rect 67730 548528 67786 548584
rect 67638 548004 67694 548040
rect 67638 547984 67640 548004
rect 67640 547984 67692 548004
rect 67692 547984 67694 548004
rect 67730 547168 67786 547224
rect 67638 546508 67694 546544
rect 67638 546488 67640 546508
rect 67640 546488 67692 546508
rect 67692 546488 67694 546508
rect 68098 545264 68154 545320
rect 68006 543904 68062 543960
rect 68006 543224 68062 543280
rect 67638 542544 67694 542600
rect 67638 541184 67694 541240
rect 67638 540096 67694 540152
rect 68926 572464 68982 572520
rect 68926 571784 68982 571840
rect 68834 558864 68890 558920
rect 68834 550704 68890 550760
rect 68742 544448 68798 544504
rect 67638 489812 67640 489832
rect 67640 489812 67692 489832
rect 67692 489812 67694 489832
rect 67638 489776 67694 489812
rect 67638 487212 67694 487248
rect 67638 487192 67640 487212
rect 67640 487192 67692 487212
rect 67692 487192 67694 487212
rect 67638 486512 67694 486568
rect 67638 485852 67694 485888
rect 67638 485832 67640 485852
rect 67640 485832 67692 485852
rect 67692 485832 67694 485852
rect 67638 485152 67694 485208
rect 67638 483928 67694 483984
rect 67638 482568 67694 482624
rect 67638 481208 67694 481264
rect 68006 481072 68062 481128
rect 67638 480156 67640 480176
rect 67640 480156 67692 480176
rect 67692 480156 67694 480176
rect 67638 480120 67694 480156
rect 67546 478488 67602 478544
rect 67546 477672 67602 477728
rect 67638 476312 67694 476368
rect 68650 484628 68706 484664
rect 68650 484608 68652 484628
rect 68652 484608 68704 484628
rect 68704 484608 68706 484628
rect 68374 476992 68430 477048
rect 68558 476992 68614 477048
rect 67730 476176 67786 476232
rect 67638 475632 67694 475688
rect 67638 474952 67694 475008
rect 67454 474272 67510 474328
rect 67454 473320 67510 473376
rect 67638 472640 67694 472696
rect 67638 471588 67640 471608
rect 67640 471588 67692 471608
rect 67692 471588 67694 471608
rect 67638 471552 67694 471588
rect 67638 471008 67694 471064
rect 67638 469648 67694 469704
rect 67730 469532 67786 469568
rect 67730 469512 67732 469532
rect 67732 469512 67784 469532
rect 67784 469512 67786 469532
rect 67730 468288 67786 468344
rect 67638 468188 67640 468208
rect 67640 468188 67692 468208
rect 67692 468188 67694 468208
rect 67638 468152 67694 468188
rect 67638 466812 67694 466848
rect 67638 466792 67640 466812
rect 67640 466792 67692 466812
rect 67692 466792 67694 466812
rect 67730 466112 67786 466168
rect 67638 465568 67694 465624
rect 67822 464072 67878 464128
rect 67638 463664 67694 463720
rect 67638 463392 67694 463448
rect 67730 462848 67786 462904
rect 67638 461352 67694 461408
rect 67638 460672 67694 460728
rect 67730 460164 67732 460184
rect 67732 460164 67784 460184
rect 67784 460164 67786 460184
rect 67730 460128 67786 460164
rect 67638 458804 67640 458824
rect 67640 458804 67692 458824
rect 67692 458804 67694 458824
rect 67362 369688 67418 369744
rect 67638 458768 67694 458804
rect 67638 458632 67694 458688
rect 67638 457952 67694 458008
rect 67730 457408 67786 457464
rect 67638 455912 67694 455968
rect 67638 455232 67694 455288
rect 67638 453872 67694 453928
rect 67638 453192 67694 453248
rect 67638 449948 67694 449984
rect 67638 449928 67640 449948
rect 67640 449928 67692 449948
rect 67692 449928 67694 449948
rect 67730 449248 67786 449304
rect 67638 449148 67640 449168
rect 67640 449148 67692 449168
rect 67692 449148 67694 449168
rect 67638 449112 67694 449148
rect 67730 448568 67786 448624
rect 67730 447752 67786 447808
rect 67638 447228 67694 447264
rect 67638 447208 67640 447228
rect 67640 447208 67692 447228
rect 67692 447208 67694 447228
rect 67730 446528 67786 446584
rect 67638 446412 67694 446448
rect 67638 446392 67640 446412
rect 67640 446392 67692 446412
rect 67692 446392 67694 446412
rect 68190 445440 68246 445496
rect 67638 443692 67694 443728
rect 67638 443672 67640 443692
rect 67640 443672 67692 443692
rect 67692 443672 67694 443692
rect 67638 442448 67694 442504
rect 67638 442312 67694 442368
rect 67638 441088 67694 441144
rect 67638 440988 67640 441008
rect 67640 440988 67692 441008
rect 67692 440988 67694 441008
rect 67638 440952 67694 440988
rect 67454 362344 67510 362400
rect 66074 331744 66130 331800
rect 67638 382472 67694 382528
rect 67638 380704 67694 380760
rect 67638 379752 67694 379808
rect 67638 377304 67694 377360
rect 67638 374448 67694 374504
rect 67730 371900 67732 371920
rect 67732 371900 67784 371920
rect 67784 371900 67786 371920
rect 67730 371864 67786 371900
rect 67638 371728 67694 371784
rect 67638 369008 67694 369064
rect 67638 366424 67694 366480
rect 68006 366016 68062 366072
rect 67638 364404 67694 364440
rect 67638 364384 67640 364404
rect 67640 364384 67692 364404
rect 67692 364384 67694 364404
rect 67730 364284 67732 364304
rect 67732 364284 67784 364304
rect 67784 364284 67786 364304
rect 67730 364248 67786 364284
rect 67638 363604 67640 363624
rect 67640 363604 67692 363624
rect 67692 363604 67694 363624
rect 67638 363568 67694 363604
rect 67638 360848 67694 360904
rect 67638 359216 67694 359272
rect 67730 358128 67786 358184
rect 67638 358028 67640 358048
rect 67640 358028 67692 358048
rect 67692 358028 67694 358048
rect 67638 357992 67694 358028
rect 67638 355816 67694 355872
rect 67730 355408 67786 355464
rect 67638 353776 67694 353832
rect 67638 352588 67640 352608
rect 67640 352588 67692 352608
rect 67692 352588 67694 352608
rect 67638 352552 67694 352588
rect 67914 351212 67970 351248
rect 67914 351192 67916 351212
rect 67916 351192 67968 351212
rect 67968 351192 67970 351212
rect 67638 350376 67694 350432
rect 67638 349052 67640 349072
rect 67640 349052 67692 349072
rect 67692 349052 67694 349072
rect 67638 349016 67694 349052
rect 67638 347112 67694 347168
rect 67730 346976 67786 347032
rect 68282 444216 68338 444272
rect 68926 543904 68982 543960
rect 68742 451288 68798 451344
rect 68558 445440 68614 445496
rect 69202 582392 69258 582448
rect 69018 543224 69074 543280
rect 69202 545264 69258 545320
rect 69202 541728 69258 541784
rect 69202 525716 69204 525736
rect 69204 525716 69256 525736
rect 69256 525716 69258 525736
rect 69202 525680 69258 525716
rect 69110 482840 69166 482896
rect 68926 444216 68982 444272
rect 68742 383424 68798 383480
rect 68374 370132 68376 370152
rect 68376 370132 68428 370152
rect 68428 370132 68430 370152
rect 68374 370096 68430 370132
rect 75090 583888 75146 583944
rect 82542 583888 82598 583944
rect 81438 583752 81494 583808
rect 82082 583752 82138 583808
rect 91650 586336 91706 586392
rect 94134 586336 94190 586392
rect 101402 584296 101458 584352
rect 103886 583752 103942 583808
rect 102598 581712 102654 581768
rect 106186 577768 106242 577824
rect 105726 548392 105782 548448
rect 74538 529080 74594 529136
rect 71778 491816 71834 491872
rect 80334 537512 80390 537568
rect 80610 499568 80666 499624
rect 81622 537376 81678 537432
rect 82266 491544 82322 491600
rect 87142 536016 87198 536072
rect 84198 494672 84254 494728
rect 88062 538056 88118 538112
rect 87418 500112 87474 500168
rect 92570 534656 92626 534712
rect 97722 500248 97778 500304
rect 96434 491444 96436 491464
rect 96436 491444 96488 491464
rect 96488 491444 96490 491464
rect 96434 491408 96490 491444
rect 96434 491272 96490 491328
rect 100942 537376 100998 537432
rect 99746 535336 99802 535392
rect 99286 491816 99342 491872
rect 99286 489368 99342 489424
rect 69202 451832 69258 451888
rect 69110 437552 69166 437608
rect 69018 434716 69074 434752
rect 69018 434696 69020 434716
rect 69020 434696 69072 434716
rect 69072 434696 69074 434716
rect 69018 433744 69074 433800
rect 99286 443672 99342 443728
rect 71042 438912 71098 438968
rect 69110 375944 69166 376000
rect 69110 374584 69166 374640
rect 68374 349732 68376 349752
rect 68376 349732 68428 349752
rect 68428 349732 68430 349752
rect 68374 349696 68430 349732
rect 68190 346332 68192 346352
rect 68192 346332 68244 346352
rect 68244 346332 68246 346352
rect 68190 346296 68246 346332
rect 68926 353096 68982 353152
rect 68742 351192 68798 351248
rect 68650 344936 68706 344992
rect 67638 343712 67694 343768
rect 67638 342896 67694 342952
rect 68650 341672 68706 341728
rect 67546 341536 67602 341592
rect 67914 340196 67970 340232
rect 67914 340176 67916 340196
rect 67916 340176 67968 340196
rect 67968 340176 67970 340196
rect 68834 349696 68890 349752
rect 68742 329024 68798 329080
rect 68834 322088 68890 322144
rect 65614 302096 65670 302152
rect 69202 370096 69258 370152
rect 73802 437552 73858 437608
rect 74538 433200 74594 433256
rect 73526 387776 73582 387832
rect 73802 387776 73858 387832
rect 75458 438132 75460 438152
rect 75460 438132 75512 438152
rect 75512 438132 75514 438152
rect 75458 438096 75514 438132
rect 78586 434716 78642 434752
rect 78586 434696 78588 434716
rect 78588 434696 78640 434716
rect 78640 434696 78642 434716
rect 76654 386416 76710 386472
rect 80978 437416 81034 437472
rect 80058 436464 80114 436520
rect 80978 436464 81034 436520
rect 80150 386960 80206 387016
rect 84198 438912 84254 438968
rect 88982 439456 89038 439512
rect 90086 397976 90142 398032
rect 93674 437416 93730 437472
rect 96618 438912 96674 438968
rect 97722 439728 97778 439784
rect 97722 438912 97778 438968
rect 96434 389816 96490 389872
rect 95882 389136 95938 389192
rect 96434 389136 96490 389192
rect 98366 437824 98422 437880
rect 99286 437824 99342 437880
rect 98642 397976 98698 398032
rect 99654 484608 99710 484664
rect 99470 443128 99526 443184
rect 99562 442448 99618 442504
rect 100758 440272 100814 440328
rect 101494 451152 101550 451208
rect 103518 537920 103574 537976
rect 102046 491408 102102 491464
rect 101954 447072 102010 447128
rect 102138 485152 102194 485208
rect 102322 484336 102378 484392
rect 102138 483792 102194 483848
rect 102138 482568 102194 482624
rect 102138 481752 102194 481808
rect 102138 481208 102194 481264
rect 102322 481072 102378 481128
rect 103426 489232 103482 489288
rect 103426 488452 103428 488472
rect 103428 488452 103480 488472
rect 103480 488452 103482 488472
rect 103426 488416 103482 488452
rect 103426 487872 103482 487928
rect 103426 486648 103482 486704
rect 103426 486512 103482 486568
rect 102138 479848 102194 479904
rect 102138 479732 102194 479768
rect 102138 479712 102140 479732
rect 102140 479712 102192 479732
rect 102192 479712 102194 479732
rect 102138 477808 102194 477864
rect 102138 476992 102194 477048
rect 102138 475632 102194 475688
rect 102138 474272 102194 474328
rect 102138 472912 102194 472968
rect 102138 471552 102194 471608
rect 102138 470192 102194 470248
rect 102138 466792 102194 466848
rect 102138 466112 102194 466168
rect 102138 465568 102194 465624
rect 102414 477128 102470 477184
rect 102322 476448 102378 476504
rect 102322 475088 102378 475144
rect 102322 472368 102378 472424
rect 102322 470872 102378 470928
rect 102874 469648 102930 469704
rect 103150 466928 103206 466984
rect 102138 464752 102194 464808
rect 102138 464108 102140 464128
rect 102140 464108 102192 464128
rect 102192 464108 102194 464128
rect 102138 464072 102194 464108
rect 102138 463392 102194 463448
rect 102138 462032 102194 462088
rect 102230 461488 102286 461544
rect 102230 460672 102286 460728
rect 102138 460128 102194 460184
rect 102138 459312 102194 459368
rect 103242 458632 103298 458688
rect 102138 457952 102194 458008
rect 102138 456592 102194 456648
rect 102230 456048 102286 456104
rect 102138 455232 102194 455288
rect 102138 454552 102194 454608
rect 102874 453348 102930 453384
rect 102874 453328 102876 453348
rect 102876 453328 102928 453348
rect 102928 453328 102930 453348
rect 102138 453228 102140 453248
rect 102140 453228 102192 453248
rect 102192 453228 102194 453248
rect 102138 453192 102194 453228
rect 102138 452548 102140 452568
rect 102140 452548 102192 452568
rect 102192 452548 102194 452568
rect 102138 452512 102194 452548
rect 102138 449248 102194 449304
rect 102138 448452 102194 448488
rect 102138 448432 102140 448452
rect 102140 448432 102192 448452
rect 102192 448432 102194 448452
rect 102230 447888 102286 447944
rect 103150 445068 103152 445088
rect 103152 445068 103204 445088
rect 103204 445068 103206 445088
rect 103150 445032 103206 445068
rect 102598 443128 102654 443184
rect 102690 442448 102746 442504
rect 103150 441768 103206 441824
rect 103150 440816 103206 440872
rect 102138 440292 102194 440328
rect 102138 440272 102140 440292
rect 102140 440272 102192 440292
rect 102192 440272 102194 440292
rect 103610 468968 103666 469024
rect 103610 450608 103666 450664
rect 103702 449792 103758 449848
rect 104806 538056 104862 538112
rect 104254 449792 104310 449848
rect 104162 444352 104218 444408
rect 103426 391176 103482 391232
rect 104990 479732 105046 479768
rect 104990 479712 104992 479732
rect 104992 479712 105044 479732
rect 105044 479712 105046 479732
rect 106370 564440 106426 564496
rect 106278 560360 106334 560416
rect 106922 583888 106978 583944
rect 108210 580080 108266 580136
rect 108854 579400 108910 579456
rect 108946 578720 109002 578776
rect 108762 577360 108818 577416
rect 108946 576000 109002 576056
rect 108946 574640 109002 574696
rect 108946 573960 109002 574016
rect 107658 573280 107714 573336
rect 108670 573280 108726 573336
rect 108946 572756 109002 572792
rect 108946 572736 108948 572756
rect 108948 572736 109000 572756
rect 109000 572736 109002 572756
rect 108946 571920 109002 571976
rect 108946 570016 109002 570072
rect 107658 569200 107714 569256
rect 108946 567840 109002 567896
rect 108946 567196 108948 567216
rect 108948 567196 109000 567216
rect 109000 567196 109002 567216
rect 108946 567160 109002 567196
rect 108854 566480 108910 566536
rect 108946 565836 108948 565856
rect 108948 565836 109000 565856
rect 109000 565836 109002 565856
rect 108946 565800 109002 565836
rect 108854 565120 108910 565176
rect 108946 563896 109002 563952
rect 108946 562400 109002 562456
rect 108946 561040 109002 561096
rect 107658 560380 107714 560416
rect 107658 560360 107660 560380
rect 107660 560360 107712 560380
rect 107712 560360 107714 560380
rect 108854 559680 108910 559736
rect 108946 559020 109002 559056
rect 108946 559000 108948 559020
rect 108948 559000 109000 559020
rect 109000 559000 109002 559020
rect 108946 558320 109002 558376
rect 107750 557640 107806 557696
rect 107014 552200 107070 552256
rect 106922 542000 106978 542056
rect 106462 540640 106518 540696
rect 106830 540640 106886 540696
rect 107658 551520 107714 551576
rect 107658 546760 107714 546816
rect 107566 470620 107622 470656
rect 107566 470600 107568 470620
rect 107568 470600 107620 470620
rect 107620 470600 107622 470620
rect 108946 556960 109002 557016
rect 107934 556280 107990 556336
rect 107842 543360 107898 543416
rect 107842 542272 107898 542328
rect 108854 555736 108910 555792
rect 108946 554240 109002 554296
rect 108946 552880 109002 552936
rect 108946 550840 109002 550896
rect 108854 550160 108910 550216
rect 108946 549480 109002 549536
rect 108946 547440 109002 547496
rect 108946 546080 109002 546136
rect 108946 545400 109002 545456
rect 108946 544720 109002 544776
rect 108946 544040 109002 544096
rect 108302 539960 108358 540016
rect 109130 581712 109186 581768
rect 109682 537784 109738 537840
rect 109314 491544 109370 491600
rect 109038 489368 109094 489424
rect 107474 449384 107530 449440
rect 107474 448568 107530 448624
rect 111890 584296 111946 584352
rect 112074 584296 112130 584352
rect 112350 545708 112352 545728
rect 112352 545708 112404 545728
rect 112404 545708 112406 545728
rect 112350 545672 112406 545708
rect 113086 545672 113142 545728
rect 111798 485696 111854 485752
rect 112442 488008 112498 488064
rect 114834 500384 114890 500440
rect 111798 386960 111854 387016
rect 115110 491136 115166 491192
rect 115846 477400 115902 477456
rect 115110 400152 115166 400208
rect 114190 390632 114246 390688
rect 114190 387912 114246 387968
rect 114926 389136 114982 389192
rect 112810 385328 112866 385384
rect 115846 388320 115902 388376
rect 115938 383968 115994 384024
rect 115294 359488 115350 359544
rect 115294 349152 115350 349208
rect 70306 345888 70362 345944
rect 70398 341672 70454 341728
rect 70490 340176 70546 340232
rect 66166 302096 66222 302152
rect 68926 299512 68982 299568
rect 67730 291080 67786 291136
rect 67638 290808 67694 290864
rect 67638 289176 67694 289232
rect 67822 288088 67878 288144
rect 67822 287428 67878 287464
rect 67822 287408 67824 287428
rect 67824 287408 67876 287428
rect 67876 287408 67878 287428
rect 67546 287000 67602 287056
rect 68926 286048 68982 286104
rect 68282 284416 68338 284472
rect 67638 283328 67694 283384
rect 67730 280472 67786 280528
rect 67638 280336 67694 280392
rect 68006 279656 68062 279712
rect 67638 279248 67694 279304
rect 67730 277752 67786 277808
rect 67638 277616 67694 277672
rect 67730 276392 67786 276448
rect 67638 276256 67694 276312
rect 67730 275168 67786 275224
rect 67638 274896 67694 274952
rect 68006 274216 68062 274272
rect 67638 273536 67694 273592
rect 67638 272312 67694 272368
rect 68190 272176 68246 272232
rect 67638 270952 67694 271008
rect 66902 270816 66958 270872
rect 68926 283736 68982 283792
rect 67730 269592 67786 269648
rect 67638 269456 67694 269512
rect 67730 268232 67786 268288
rect 67638 268096 67694 268152
rect 67638 267028 67694 267064
rect 67638 267008 67640 267028
rect 67640 267008 67692 267028
rect 67692 267008 67694 267028
rect 67638 266364 67640 266384
rect 67640 266364 67692 266384
rect 67692 266364 67694 266384
rect 67638 266328 67694 266364
rect 67730 265512 67786 265568
rect 67822 265376 67878 265432
rect 67638 264868 67640 264888
rect 67640 264868 67692 264888
rect 67692 264868 67694 264888
rect 67638 264832 67694 264868
rect 67638 263628 67694 263664
rect 67638 263608 67640 263628
rect 67640 263608 67692 263628
rect 67692 263608 67694 263628
rect 67730 262792 67786 262848
rect 67638 262268 67694 262304
rect 67638 262248 67640 262268
rect 67640 262248 67692 262268
rect 67692 262248 67694 262268
rect 67730 261432 67786 261488
rect 67638 260924 67640 260944
rect 67640 260924 67692 260944
rect 67692 260924 67694 260944
rect 67638 260888 67694 260924
rect 67638 260788 67640 260808
rect 67640 260788 67692 260808
rect 67692 260788 67694 260808
rect 67638 260752 67694 260788
rect 67638 259528 67694 259584
rect 67730 258712 67786 258768
rect 67638 258168 67694 258224
rect 67914 257216 67970 257272
rect 67638 256808 67694 256864
rect 67638 255856 67694 255912
rect 67730 255332 67786 255368
rect 67730 255312 67732 255332
rect 67732 255312 67784 255332
rect 67784 255312 67786 255332
rect 67638 255212 67640 255232
rect 67640 255212 67692 255232
rect 67692 255212 67694 255232
rect 67638 255176 67694 255212
rect 67638 253972 67694 254008
rect 67638 253952 67640 253972
rect 67640 253952 67692 253972
rect 67692 253952 67694 253972
rect 67638 253136 67694 253192
rect 67730 251776 67786 251832
rect 67638 251368 67694 251424
rect 68650 250416 68706 250472
rect 67638 249872 67694 249928
rect 67730 249056 67786 249112
rect 67638 248512 67694 248568
rect 67730 247696 67786 247752
rect 67638 247172 67694 247208
rect 67638 247152 67640 247172
rect 67640 247152 67692 247172
rect 67692 247152 67694 247172
rect 67730 246336 67786 246392
rect 67638 245792 67694 245848
rect 67454 244296 67510 244352
rect 67546 243616 67602 243672
rect 67638 243072 67694 243128
rect 67638 241848 67694 241904
rect 68650 239400 68706 239456
rect 70398 302232 70454 302288
rect 73894 338000 73950 338056
rect 74446 338000 74502 338056
rect 71042 301416 71098 301472
rect 71134 292304 71190 292360
rect 75918 339632 75974 339688
rect 75274 318008 75330 318064
rect 74446 315288 74502 315344
rect 77114 339632 77170 339688
rect 73250 300872 73306 300928
rect 75826 294072 75882 294128
rect 79414 316648 79470 316704
rect 91006 333240 91062 333296
rect 91282 294480 91338 294536
rect 102138 338136 102194 338192
rect 101586 297336 101642 297392
rect 96710 295976 96766 296032
rect 95790 294208 95846 294264
rect 97078 292576 97134 292632
rect 100942 295432 100998 295488
rect 109958 339360 110014 339416
rect 108026 293936 108082 293992
rect 111246 295296 111302 295352
rect 113178 296792 113234 296848
rect 111890 292712 111946 292768
rect 117410 489132 117412 489152
rect 117412 489132 117464 489152
rect 117464 489132 117466 489152
rect 117410 489096 117466 489132
rect 117042 481480 117098 481536
rect 116030 370368 116086 370424
rect 116214 391176 116270 391232
rect 117686 477400 117742 477456
rect 117318 379480 117374 379536
rect 116214 371320 116270 371376
rect 116214 370640 116270 370696
rect 117318 368600 117374 368656
rect 117318 367920 117374 367976
rect 117410 367240 117466 367296
rect 117318 365880 117374 365936
rect 117318 365200 117374 365256
rect 117318 362480 117374 362536
rect 117318 361800 117374 361856
rect 117318 361120 117374 361176
rect 116122 357040 116178 357096
rect 118790 488552 118846 488608
rect 121550 583752 121606 583808
rect 117686 386280 117742 386336
rect 118514 384920 118570 384976
rect 118606 383596 118608 383616
rect 118608 383596 118660 383616
rect 118660 383596 118662 383616
rect 118606 383560 118662 383596
rect 118606 381540 118662 381576
rect 118606 381520 118608 381540
rect 118608 381520 118660 381540
rect 118660 381520 118662 381540
rect 118606 380860 118662 380896
rect 118606 380840 118608 380860
rect 118608 380840 118660 380860
rect 118660 380840 118662 380860
rect 118330 379480 118386 379536
rect 118606 378836 118608 378856
rect 118608 378836 118660 378856
rect 118660 378836 118662 378856
rect 118606 378800 118662 378836
rect 118606 378156 118608 378176
rect 118608 378156 118660 378176
rect 118660 378156 118662 378176
rect 118606 378120 118662 378156
rect 118422 376780 118478 376816
rect 118422 376760 118424 376780
rect 118424 376760 118476 376780
rect 118476 376760 118478 376780
rect 117778 376080 117834 376136
rect 118606 375400 118662 375456
rect 118606 374040 118662 374096
rect 118606 373360 118662 373416
rect 117870 370640 117926 370696
rect 118054 369960 118110 370016
rect 117686 363160 117742 363216
rect 117870 359080 117926 359136
rect 118606 358400 118662 358456
rect 118146 357040 118202 357096
rect 118606 356360 118662 356416
rect 117594 355680 117650 355736
rect 118606 355680 118662 355736
rect 118606 354320 118662 354376
rect 118514 353640 118570 353696
rect 118606 352960 118662 353016
rect 117502 351600 117558 351656
rect 118606 351600 118662 351656
rect 118054 350920 118110 350976
rect 118606 350240 118662 350296
rect 117870 348880 117926 348936
rect 118606 348200 118662 348256
rect 117410 347520 117466 347576
rect 118514 346160 118570 346216
rect 118606 345480 118662 345536
rect 118606 344800 118662 344856
rect 118606 343440 118662 343496
rect 117778 342760 117834 342816
rect 118606 342080 118662 342136
rect 117502 340720 117558 340776
rect 117318 340040 117374 340096
rect 118422 340040 118478 340096
rect 114558 291896 114614 291952
rect 119066 364792 119122 364848
rect 118882 359760 118938 359816
rect 119342 338000 119398 338056
rect 117318 327664 117374 327720
rect 118882 307672 118938 307728
rect 119894 295568 119950 295624
rect 118330 292848 118386 292904
rect 69846 288768 69902 288824
rect 69110 286728 69166 286784
rect 69018 282104 69074 282160
rect 69018 274216 69074 274272
rect 68926 232600 68982 232656
rect 69110 252592 69166 252648
rect 122102 572736 122158 572792
rect 120262 386960 120318 387016
rect 120170 338000 120226 338056
rect 122746 485696 122802 485752
rect 120170 256400 120226 256456
rect 120170 250960 120226 251016
rect 120078 247560 120134 247616
rect 69202 244976 69258 245032
rect 72606 238584 72662 238640
rect 80150 229744 80206 229800
rect 84290 220088 84346 220144
rect 90362 237904 90418 237960
rect 97078 177656 97134 177712
rect 106922 197920 106978 197976
rect 102046 177656 102102 177712
rect 106186 177656 106242 177712
rect 108118 176976 108174 177032
rect 110694 177656 110750 177712
rect 100666 176704 100722 176760
rect 103334 176704 103390 176760
rect 107014 176704 107070 176760
rect 109958 176704 110014 176760
rect 113822 238584 113878 238640
rect 114650 226208 114706 226264
rect 117042 238448 117098 238504
rect 119342 235864 119398 235920
rect 122930 483248 122986 483304
rect 122102 387640 122158 387696
rect 122838 387640 122894 387696
rect 122102 386572 122158 386608
rect 122102 386552 122104 386572
rect 122104 386552 122156 386572
rect 122156 386552 122158 386572
rect 122194 380160 122250 380216
rect 121550 291780 121606 291816
rect 121550 291760 121552 291780
rect 121552 291760 121604 291780
rect 121604 291760 121606 291780
rect 121550 291080 121606 291136
rect 121550 287680 121606 287736
rect 121550 287020 121606 287056
rect 121734 289040 121790 289096
rect 121826 288360 121882 288416
rect 121550 287000 121552 287020
rect 121552 287000 121604 287020
rect 121604 287000 121606 287020
rect 121550 286340 121606 286376
rect 121550 286320 121552 286340
rect 121552 286320 121604 286340
rect 121604 286320 121606 286340
rect 121550 284960 121606 285016
rect 121642 284316 121644 284336
rect 121644 284316 121696 284336
rect 121696 284316 121698 284336
rect 121642 284280 121698 284316
rect 121550 283620 121606 283656
rect 121550 283600 121552 283620
rect 121552 283600 121604 283620
rect 121604 283600 121606 283620
rect 121550 282940 121606 282976
rect 121550 282920 121552 282940
rect 121552 282920 121604 282940
rect 121604 282920 121606 282940
rect 121642 282240 121698 282296
rect 121550 281580 121606 281616
rect 121550 281560 121552 281580
rect 121552 281560 121604 281580
rect 121604 281560 121606 281580
rect 121642 280880 121698 280936
rect 121550 280236 121552 280256
rect 121552 280236 121604 280256
rect 121604 280236 121606 280256
rect 121550 280200 121606 280236
rect 121642 279520 121698 279576
rect 121550 278860 121606 278896
rect 121550 278840 121552 278860
rect 121552 278840 121604 278860
rect 121604 278840 121606 278860
rect 121550 277480 121606 277536
rect 121734 276800 121790 276856
rect 121550 276120 121606 276176
rect 121642 275440 121698 275496
rect 121550 274760 121606 274816
rect 121550 274080 121606 274136
rect 121550 273400 121606 273456
rect 121550 272720 121606 272776
rect 121550 272040 121606 272096
rect 121550 271360 121606 271416
rect 121642 270000 121698 270056
rect 121550 269320 121606 269376
rect 121642 268640 121698 268696
rect 121550 267960 121606 268016
rect 121642 267280 121698 267336
rect 121550 266600 121606 266656
rect 121642 265920 121698 265976
rect 121550 265240 121606 265296
rect 121734 264560 121790 264616
rect 121550 263880 121606 263936
rect 121550 263200 121606 263256
rect 121550 262520 121606 262576
rect 121734 261840 121790 261896
rect 121642 261160 121698 261216
rect 121550 260480 121606 260536
rect 121550 259800 121606 259856
rect 121550 259120 121606 259176
rect 121642 258440 121698 258496
rect 121642 257760 121698 257816
rect 121550 257080 121606 257136
rect 121642 256400 121698 256456
rect 121550 254360 121606 254416
rect 121550 253680 121606 253736
rect 121642 253000 121698 253056
rect 121550 252320 121606 252376
rect 121550 251640 121606 251696
rect 122562 314200 122618 314256
rect 124402 553968 124458 554024
rect 123758 438948 123760 438968
rect 123760 438948 123812 438968
rect 123812 438948 123814 438968
rect 123758 438912 123814 438948
rect 123022 378936 123078 378992
rect 124954 541592 125010 541648
rect 122378 289448 122434 289504
rect 122746 285640 122802 285696
rect 122286 255040 122342 255096
rect 122102 250960 122158 251016
rect 121550 250280 121606 250336
rect 121550 248920 121606 248976
rect 121458 248240 121514 248296
rect 121642 247560 121698 247616
rect 121550 246880 121606 246936
rect 121458 246200 121514 246256
rect 121642 245520 121698 245576
rect 121550 244840 121606 244896
rect 121458 244160 121514 244216
rect 121458 242836 121460 242856
rect 121460 242836 121512 242856
rect 121512 242836 121514 242856
rect 121458 242800 121514 242836
rect 121366 241440 121422 241496
rect 121458 240760 121514 240816
rect 121734 243516 121736 243536
rect 121736 243516 121788 243536
rect 121788 243516 121790 243536
rect 121734 243480 121790 243516
rect 121458 240080 121514 240136
rect 124034 248240 124090 248296
rect 125598 453348 125654 453384
rect 125598 453328 125600 453348
rect 125600 453328 125652 453348
rect 125652 453328 125654 453348
rect 124954 444896 125010 444952
rect 124402 315988 124458 316024
rect 124402 315968 124404 315988
rect 124404 315968 124456 315988
rect 124456 315968 124458 315988
rect 126150 342372 126206 342408
rect 126150 342352 126152 342372
rect 126152 342352 126204 342372
rect 126204 342352 126206 342372
rect 128450 498788 128452 498808
rect 128452 498788 128504 498808
rect 128504 498788 128506 498808
rect 128450 498752 128506 498788
rect 127254 312432 127310 312488
rect 127622 238448 127678 238504
rect 129830 388320 129886 388376
rect 130382 388320 130438 388376
rect 128450 238584 128506 238640
rect 131670 319368 131726 319424
rect 131118 297336 131174 297392
rect 134522 385600 134578 385656
rect 133878 296928 133934 296984
rect 114374 177656 114430 177712
rect 118514 177656 118570 177712
rect 114006 176976 114062 177032
rect 115846 176976 115902 177032
rect 121458 179424 121514 179480
rect 121366 177656 121422 177712
rect 126886 177656 126942 177712
rect 124126 177112 124182 177168
rect 136914 390496 136970 390552
rect 137098 326440 137154 326496
rect 136638 226208 136694 226264
rect 136638 225664 136694 225720
rect 299478 541592 299534 541648
rect 143538 385600 143594 385656
rect 144918 448568 144974 448624
rect 146206 374584 146262 374640
rect 144182 283464 144238 283520
rect 150530 368328 150586 368384
rect 151818 373224 151874 373280
rect 150990 368328 151046 368384
rect 150990 367648 151046 367704
rect 147034 193840 147090 193896
rect 152462 291896 152518 291952
rect 130750 177656 130806 177712
rect 132406 177656 132462 177712
rect 162122 177248 162178 177304
rect 119526 176704 119582 176760
rect 122102 176704 122158 176760
rect 124494 176704 124550 176760
rect 127898 176704 127954 176760
rect 133142 176724 133198 176760
rect 133142 176704 133144 176724
rect 133144 176704 133196 176724
rect 133196 176704 133198 176724
rect 134430 176704 134486 176760
rect 136086 176740 136088 176760
rect 136088 176740 136140 176760
rect 136140 176740 136142 176760
rect 136086 176704 136142 176740
rect 104622 175480 104678 175536
rect 116950 175480 117006 175536
rect 128174 175480 128230 175536
rect 129462 175480 129518 175536
rect 148230 175480 148286 175536
rect 158902 175480 158958 175536
rect 164882 173984 164938 174040
rect 165618 173984 165674 174040
rect 66074 129240 66130 129296
rect 65522 128016 65578 128072
rect 65982 102312 66038 102368
rect 67362 126248 67418 126304
rect 66166 125160 66222 125216
rect 66074 94696 66130 94752
rect 67546 123528 67602 123584
rect 67454 122576 67510 122632
rect 67362 94832 67418 94888
rect 67454 91024 67510 91080
rect 67638 120808 67694 120864
rect 67546 89664 67602 89720
rect 67730 100680 67786 100736
rect 167642 171536 167698 171592
rect 126518 94152 126574 94208
rect 152094 94172 152150 94208
rect 152094 94152 152096 94172
rect 152096 94152 152148 94172
rect 152148 94152 152150 94172
rect 112350 94016 112406 94072
rect 126702 94036 126758 94072
rect 126702 94016 126704 94036
rect 126704 94016 126756 94036
rect 126756 94016 126758 94036
rect 96158 93900 96214 93936
rect 96158 93880 96160 93900
rect 96160 93880 96212 93900
rect 96212 93880 96214 93900
rect 100942 93472 100998 93528
rect 109222 93472 109278 93528
rect 116766 93472 116822 93528
rect 121734 93472 121790 93528
rect 133142 93492 133198 93528
rect 133142 93472 133144 93492
rect 133144 93472 133196 93492
rect 133196 93472 133198 93492
rect 103334 93200 103390 93256
rect 151726 93472 151782 93528
rect 74814 92384 74870 92440
rect 85854 92384 85910 92440
rect 88062 92384 88118 92440
rect 88982 92420 88984 92440
rect 88984 92420 89036 92440
rect 89036 92420 89038 92440
rect 88982 92384 89038 92420
rect 97538 92384 97594 92440
rect 98826 92384 98882 92440
rect 85486 91160 85542 91216
rect 66166 84088 66222 84144
rect 86774 91160 86830 91216
rect 90730 91704 90786 91760
rect 95054 91296 95110 91352
rect 92386 91160 92442 91216
rect 93766 91160 93822 91216
rect 95146 91160 95202 91216
rect 97814 91160 97870 91216
rect 103242 92248 103298 92304
rect 99194 91296 99250 91352
rect 100574 91296 100630 91352
rect 101862 91296 101918 91352
rect 99286 91160 99342 91216
rect 99194 82728 99250 82784
rect 100666 91160 100722 91216
rect 102046 91160 102102 91216
rect 99286 80008 99342 80064
rect 110142 93200 110198 93256
rect 106094 91296 106150 91352
rect 107566 91296 107622 91352
rect 104254 91160 104310 91216
rect 104806 91160 104862 91216
rect 106186 91160 106242 91216
rect 107474 91160 107530 91216
rect 107934 91160 107990 91216
rect 108946 91160 109002 91216
rect 106186 81368 106242 81424
rect 114466 92384 114522 92440
rect 114926 92384 114982 92440
rect 115478 92384 115534 92440
rect 118054 92404 118110 92440
rect 118054 92384 118056 92404
rect 118056 92384 118108 92404
rect 118108 92384 118110 92404
rect 110326 91160 110382 91216
rect 110694 91160 110750 91216
rect 111706 91160 111762 91216
rect 113086 91160 113142 91216
rect 113362 91160 113418 91216
rect 114374 91160 114430 91216
rect 108946 79872 109002 79928
rect 110694 88168 110750 88224
rect 132406 92384 132462 92440
rect 151542 92384 151598 92440
rect 122838 92112 122894 92168
rect 119802 91568 119858 91624
rect 115754 91160 115810 91216
rect 117134 91160 117190 91216
rect 118606 91160 118662 91216
rect 120722 91296 120778 91352
rect 119986 91160 120042 91216
rect 121366 91160 121422 91216
rect 136454 91568 136510 91624
rect 124034 91296 124090 91352
rect 125414 91296 125470 91352
rect 124126 91160 124182 91216
rect 125506 91160 125562 91216
rect 126518 91160 126574 91216
rect 129462 91160 129518 91216
rect 130750 91160 130806 91216
rect 135166 91160 135222 91216
rect 130750 85448 130806 85504
rect 151634 92112 151690 92168
rect 67638 64096 67694 64152
rect 167642 108704 167698 108760
rect 168010 111732 168012 111752
rect 168012 111732 168064 111752
rect 168064 111732 168066 111752
rect 168010 111696 168066 111732
rect 168102 110064 168158 110120
rect 170494 90888 170550 90944
rect 170402 84768 170458 84824
rect 173438 94696 173494 94752
rect 178774 294208 178830 294264
rect 184294 177248 184350 177304
rect 188434 294072 188490 294128
rect 188434 93472 188490 93528
rect 198094 86128 198150 86184
rect 202234 292712 202290 292768
rect 202234 90344 202290 90400
rect 203614 93608 203670 93664
rect 206558 94832 206614 94888
rect 209226 89664 209282 89720
rect 213918 176160 213974 176216
rect 213274 175344 213330 175400
rect 213918 175072 213974 175128
rect 214010 174664 214066 174720
rect 213918 173712 213974 173768
rect 214010 173304 214066 173360
rect 214102 172352 214158 172408
rect 213918 171944 213974 172000
rect 213918 171028 213920 171048
rect 213920 171028 213972 171048
rect 213972 171028 213974 171048
rect 213918 170992 213974 171028
rect 213918 169652 213974 169688
rect 213918 169632 213920 169652
rect 213920 169632 213972 169652
rect 213972 169632 213974 169652
rect 214010 169360 214066 169416
rect 213918 168000 213974 168056
rect 214010 167864 214066 167920
rect 213918 166640 213974 166696
rect 213366 166096 213422 166152
rect 213918 165280 213974 165336
rect 214010 164736 214066 164792
rect 213918 163920 213974 163976
rect 213918 162560 213974 162616
rect 213918 161372 213920 161392
rect 213920 161372 213972 161392
rect 213972 161372 213974 161392
rect 213918 161336 213974 161372
rect 214746 170720 214802 170776
rect 214654 166912 214710 166968
rect 214562 160792 214618 160848
rect 214102 160656 214158 160712
rect 213918 159840 213974 159896
rect 214010 159432 214066 159488
rect 213918 158652 213920 158672
rect 213920 158652 213972 158672
rect 213972 158652 213974 158672
rect 213918 158616 213974 158652
rect 214102 158072 214158 158128
rect 213918 157276 213974 157312
rect 213918 157256 213920 157276
rect 213920 157256 213972 157276
rect 213972 157256 213974 157276
rect 214010 156848 214066 156904
rect 213274 155896 213330 155952
rect 213918 155488 213974 155544
rect 214010 153856 214066 153912
rect 213918 153332 213974 153368
rect 213918 153312 213920 153332
rect 213920 153312 213972 153332
rect 213972 153312 213974 153332
rect 214010 152632 214066 152688
rect 213918 151952 213974 152008
rect 213458 151816 213514 151872
rect 213274 142296 213330 142352
rect 215022 150728 215078 150784
rect 213918 150592 213974 150648
rect 213918 150048 213974 150104
rect 214010 149504 214066 149560
rect 213918 148824 213974 148880
rect 213918 148008 213974 148064
rect 214010 146648 214066 146704
rect 213918 146376 213974 146432
rect 214654 145288 214710 145344
rect 214010 143928 214066 143984
rect 213918 143520 213974 143576
rect 213918 142704 213974 142760
rect 214010 141344 214066 141400
rect 213918 140820 213974 140856
rect 213918 140800 213920 140820
rect 213920 140800 213972 140820
rect 213972 140800 213974 140820
rect 214562 139984 214618 140040
rect 213918 139460 213974 139496
rect 213918 139440 213920 139460
rect 213920 139440 213972 139460
rect 213972 139440 213974 139460
rect 214010 138760 214066 138816
rect 213918 138100 213974 138136
rect 213918 138080 213920 138100
rect 213920 138080 213972 138100
rect 213972 138080 213974 138100
rect 213918 137400 213974 137456
rect 214010 136740 214066 136776
rect 214010 136720 214012 136740
rect 214012 136720 214064 136740
rect 214064 136720 214066 136740
rect 214010 136040 214066 136096
rect 213918 135380 213974 135416
rect 213918 135360 213920 135380
rect 213920 135360 213972 135380
rect 213972 135360 213974 135380
rect 213918 134000 213974 134056
rect 213918 132524 213974 132560
rect 213918 132504 213920 132524
rect 213920 132504 213972 132524
rect 213972 132504 213974 132524
rect 213918 131164 213974 131200
rect 213918 131144 213920 131164
rect 213920 131144 213972 131164
rect 213972 131144 213974 131164
rect 213918 129804 213974 129840
rect 213918 129784 213920 129804
rect 213920 129784 213972 129804
rect 213972 129784 213974 129804
rect 213918 128832 213974 128888
rect 213918 127064 213974 127120
rect 214010 126112 214066 126168
rect 213918 125724 213974 125760
rect 213918 125704 213920 125724
rect 213920 125704 213972 125724
rect 213972 125704 213974 125724
rect 214010 124752 214066 124808
rect 213918 124344 213974 124400
rect 214010 123528 214066 123584
rect 213918 123120 213974 123176
rect 214010 122168 214066 122224
rect 213918 121508 213974 121544
rect 213918 121488 213920 121508
rect 213920 121488 213972 121508
rect 213972 121488 213974 121508
rect 213918 120808 213974 120864
rect 214010 120264 214066 120320
rect 214010 119584 214066 119640
rect 213918 118904 213974 118960
rect 214102 119040 214158 119096
rect 214010 117544 214066 117600
rect 213918 117308 213920 117328
rect 213920 117308 213972 117328
rect 213972 117308 213974 117328
rect 213918 117272 213974 117308
rect 214010 116184 214066 116240
rect 213918 115948 213920 115968
rect 213920 115948 213972 115968
rect 213972 115948 213974 115968
rect 213918 115912 213974 115948
rect 214010 114960 214066 115016
rect 213918 114572 213974 114608
rect 213918 114552 213920 114572
rect 213920 114552 213972 114572
rect 213972 114552 213974 114572
rect 214010 113600 214066 113656
rect 213918 113212 213974 113248
rect 213918 113192 213920 113212
rect 213920 113192 213972 113212
rect 213972 113192 213974 113212
rect 213458 112240 213514 112296
rect 213918 111852 213974 111888
rect 213918 111832 213920 111852
rect 213920 111832 213972 111852
rect 213972 111832 213974 111852
rect 214010 110880 214066 110936
rect 213918 110508 213920 110528
rect 213920 110508 213972 110528
rect 213972 110508 213974 110528
rect 213918 110472 213974 110508
rect 213918 109248 213974 109304
rect 214010 108296 214066 108352
rect 213918 107888 213974 107944
rect 214010 106936 214066 106992
rect 213918 106412 213974 106448
rect 213918 106392 213920 106412
rect 213920 106392 213972 106412
rect 213972 106392 213974 106412
rect 214010 105712 214066 105768
rect 213918 105052 213974 105088
rect 213918 105032 213920 105052
rect 213920 105032 213972 105052
rect 213972 105032 213974 105052
rect 214102 105168 214158 105224
rect 213918 103808 213974 103864
rect 213918 102584 213974 102640
rect 214746 135496 214802 135552
rect 214654 130056 214710 130112
rect 214746 109656 214802 109712
rect 214562 101360 214618 101416
rect 213918 100816 213974 100872
rect 214102 99728 214158 99784
rect 214010 98368 214066 98424
rect 213918 97960 213974 98016
rect 214286 99456 214342 99512
rect 214654 96600 214710 96656
rect 214562 95784 214618 95840
rect 214838 101088 214894 101144
rect 216678 97008 216734 97064
rect 220082 180104 220138 180160
rect 224222 179968 224278 180024
rect 272522 369008 272578 369064
rect 228362 177384 228418 177440
rect 222842 177248 222898 177304
rect 238022 177520 238078 177576
rect 242162 181328 242218 181384
rect 247682 178608 247738 178664
rect 246486 176568 246542 176624
rect 228454 175888 228510 175944
rect 249154 175208 249210 175264
rect 249154 174648 249210 174704
rect 249338 175616 249394 175672
rect 249246 173304 249302 173360
rect 249430 172760 249486 172816
rect 249798 168136 249854 168192
rect 250074 171400 250130 171456
rect 249982 160520 250038 160576
rect 249890 154400 249946 154456
rect 250442 144608 250498 144664
rect 246486 94424 246542 94480
rect 246394 77832 246450 77888
rect 250810 153720 250866 153776
rect 250626 144064 250682 144120
rect 250534 136584 250590 136640
rect 249798 97008 249854 97064
rect 251270 157800 251326 157856
rect 252466 172352 252522 172408
rect 252374 171808 252430 171864
rect 252466 170856 252522 170912
rect 252374 170448 252430 170504
rect 252466 170076 252468 170096
rect 252468 170076 252520 170096
rect 252520 170076 252522 170096
rect 252466 170040 252522 170076
rect 252466 169088 252522 169144
rect 252374 168544 252430 168600
rect 252374 167592 252430 167648
rect 252466 167184 252522 167240
rect 252466 166640 252522 166696
rect 252466 165688 252522 165744
rect 252282 164736 252338 164792
rect 252466 165280 252522 165336
rect 252374 164328 252430 164384
rect 252466 163920 252522 163976
rect 252374 163376 252430 163432
rect 252282 162968 252338 163024
rect 252558 162424 252614 162480
rect 252466 162016 252522 162072
rect 252374 161472 252430 161528
rect 252466 160248 252522 160304
rect 251730 159568 251786 159624
rect 252466 158752 252522 158808
rect 252466 158208 252522 158264
rect 251362 156304 251418 156360
rect 251178 147872 251234 147928
rect 251454 146920 251510 146976
rect 251178 145016 251234 145072
rect 250810 141752 250866 141808
rect 251178 140800 251234 140856
rect 252466 156848 252522 156904
rect 252650 155896 252706 155952
rect 252466 155352 252522 155408
rect 252374 154944 252430 155000
rect 252466 153992 252522 154048
rect 252098 153448 252154 153504
rect 252282 153040 252338 153096
rect 252466 152632 252522 152688
rect 252374 152088 252430 152144
rect 252466 151716 252468 151736
rect 252468 151716 252520 151736
rect 252520 151716 252522 151736
rect 252466 151680 252522 151716
rect 252466 151136 252522 151192
rect 252282 150728 252338 150784
rect 252282 149776 252338 149832
rect 252466 150184 252522 150240
rect 252374 149232 252430 149288
rect 252466 148824 252522 148880
rect 252374 148280 252430 148336
rect 252466 147500 252468 147520
rect 252468 147500 252520 147520
rect 252520 147500 252522 147520
rect 252466 147464 252522 147500
rect 252374 146512 252430 146568
rect 252466 145968 252522 146024
rect 252374 145560 252430 145616
rect 251822 138488 251878 138544
rect 251178 111152 251234 111208
rect 251730 109248 251786 109304
rect 250718 105984 250774 106040
rect 252466 143656 252522 143712
rect 252466 143112 252522 143168
rect 252374 142704 252430 142760
rect 252834 169496 252890 169552
rect 252466 141344 252522 141400
rect 252466 140392 252522 140448
rect 252374 139848 252430 139904
rect 252558 139440 252614 139496
rect 252466 138896 252522 138952
rect 252466 137964 252522 138000
rect 252466 137944 252468 137964
rect 252468 137944 252520 137964
rect 252520 137944 252522 137964
rect 252098 131416 252154 131472
rect 252006 124752 252062 124808
rect 252466 136176 252522 136232
rect 252374 135632 252430 135688
rect 252282 135224 252338 135280
rect 252466 134680 252522 134736
rect 252374 134272 252430 134328
rect 252466 133748 252522 133784
rect 252466 133728 252468 133748
rect 252468 133728 252520 133748
rect 252520 133728 252522 133748
rect 252374 133320 252430 133376
rect 252282 132776 252338 132832
rect 252466 132388 252522 132424
rect 252466 132368 252468 132388
rect 252468 132368 252520 132388
rect 252520 132368 252522 132388
rect 252374 131824 252430 131880
rect 252374 130872 252430 130928
rect 252466 130464 252522 130520
rect 252282 130056 252338 130112
rect 252466 129512 252522 129568
rect 252374 129104 252430 129160
rect 252282 128560 252338 128616
rect 252466 128152 252522 128208
rect 252282 127608 252338 127664
rect 252374 127200 252430 127256
rect 252466 126656 252522 126712
rect 252374 126248 252430 126304
rect 252282 125704 252338 125760
rect 252466 125296 252522 125352
rect 252190 124344 252246 124400
rect 252466 123936 252522 123992
rect 252374 123392 252430 123448
rect 252282 122984 252338 123040
rect 252466 122440 252522 122496
rect 252374 122032 252430 122088
rect 252282 121488 252338 121544
rect 252098 121080 252154 121136
rect 252466 120536 252522 120592
rect 251914 120128 251970 120184
rect 251914 107888 251970 107944
rect 252282 119176 252338 119232
rect 252466 119584 252522 119640
rect 252374 118768 252430 118824
rect 252466 118224 252522 118280
rect 252374 117816 252430 117872
rect 252282 117272 252338 117328
rect 252466 116320 252522 116376
rect 252374 115912 252430 115968
rect 252466 115368 252522 115424
rect 252374 114960 252430 115016
rect 252466 114452 252468 114472
rect 252468 114452 252520 114472
rect 252520 114452 252522 114472
rect 252466 114416 252522 114452
rect 253202 114008 253258 114064
rect 252282 113464 252338 113520
rect 252282 113076 252338 113112
rect 252282 113056 252284 113076
rect 252284 113056 252336 113076
rect 252336 113056 252338 113076
rect 252374 112648 252430 112704
rect 252466 112104 252522 112160
rect 252374 111716 252430 111752
rect 252374 111696 252376 111716
rect 252376 111696 252428 111716
rect 252428 111696 252430 111716
rect 252466 110744 252522 110800
rect 252466 110200 252522 110256
rect 252466 108876 252468 108896
rect 252468 108876 252520 108896
rect 252520 108876 252522 108896
rect 252466 108840 252522 108876
rect 252374 108296 252430 108352
rect 252466 107480 252522 107536
rect 252374 106936 252430 106992
rect 252466 106528 252522 106584
rect 252282 105576 252338 105632
rect 252006 105032 252062 105088
rect 252282 104624 252338 104680
rect 252374 104080 252430 104136
rect 252466 103672 252522 103728
rect 251822 102720 251878 102776
rect 252466 103128 252522 103184
rect 252374 102176 252430 102232
rect 251730 101360 251786 101416
rect 251362 97960 251418 98016
rect 252466 101768 252522 101824
rect 252374 100816 252430 100872
rect 252282 99864 252338 99920
rect 252466 100408 252522 100464
rect 252374 99456 252430 99512
rect 252466 98912 252522 98968
rect 252374 98504 252430 98560
rect 252190 97552 252246 97608
rect 252466 97280 252522 97336
rect 252466 96600 252522 96656
rect 251178 96192 251234 96248
rect 251178 86128 251234 86184
rect 242898 10920 242954 10976
rect 243542 10920 243598 10976
rect 258906 139984 258962 140040
rect 259550 65612 259606 65648
rect 259550 65592 259552 65612
rect 259552 65592 259604 65612
rect 259604 65592 259606 65612
rect 258446 10940 258502 10976
rect 258446 10920 258448 10940
rect 258448 10920 258500 10940
rect 258500 10920 258502 10940
rect 263506 81504 263562 81560
rect 260746 11736 260802 11792
rect 258262 3440 258318 3496
rect 259366 3440 259422 3496
rect 259458 3304 259514 3360
rect 260746 3304 260802 3360
rect 263598 56480 263654 56536
rect 263690 24148 263692 24168
rect 263692 24148 263744 24168
rect 263744 24148 263746 24168
rect 263690 24112 263746 24148
rect 264610 11736 264666 11792
rect 262954 3440 263010 3496
rect 263506 3440 263562 3496
rect 267646 81368 267702 81424
rect 267738 57976 267794 58032
rect 269118 47524 269174 47560
rect 269118 47504 269120 47524
rect 269120 47504 269172 47524
rect 269172 47504 269174 47524
rect 268382 12280 268438 12336
rect 266542 3440 266598 3496
rect 267646 3440 267702 3496
rect 270590 26968 270646 27024
rect 270314 11736 270370 11792
rect 273258 41248 273314 41304
rect 271786 12688 271842 12744
rect 271234 3440 271290 3496
rect 271786 3440 271842 3496
rect 274178 71032 274234 71088
rect 274178 41248 274234 41304
rect 283562 367648 283618 367704
rect 276754 149640 276810 149696
rect 278318 137264 278374 137320
rect 280894 330384 280950 330440
rect 284390 49020 284446 49056
rect 284390 49000 284392 49020
rect 284392 49000 284444 49020
rect 284444 49000 284446 49020
rect 286322 67496 286378 67552
rect 286966 67496 287022 67552
rect 285586 11736 285642 11792
rect 284298 3440 284354 3496
rect 285586 3440 285642 3496
rect 293222 335960 293278 336016
rect 289174 177384 289230 177440
rect 293406 111016 293462 111072
rect 301502 370504 301558 370560
rect 298190 43288 298246 43344
rect 299662 39364 299718 39400
rect 299662 39344 299664 39364
rect 299664 39344 299716 39364
rect 299716 39344 299718 39364
rect 299386 11736 299442 11792
rect 304262 184184 304318 184240
rect 304354 175752 304410 175808
rect 300766 11736 300822 11792
rect 300122 9560 300178 9616
rect 300674 9560 300730 9616
rect 299662 3576 299718 3632
rect 298466 3440 298522 3496
rect 299386 3440 299442 3496
rect 300766 3576 300822 3632
rect 302238 40724 302294 40760
rect 302238 40704 302240 40724
rect 302240 40704 302292 40724
rect 302292 40704 302294 40724
rect 303526 11736 303582 11792
rect 305734 173984 305790 174040
rect 306562 172216 306618 172272
rect 307390 175208 307446 175264
rect 307482 174800 307538 174856
rect 307390 173984 307446 174040
rect 307666 174392 307722 174448
rect 307574 174020 307576 174040
rect 307576 174020 307628 174040
rect 307628 174020 307630 174040
rect 307574 173984 307630 174020
rect 307574 173576 307630 173632
rect 307482 173168 307538 173224
rect 307666 172624 307722 172680
rect 307666 171808 307722 171864
rect 307298 171400 307354 171456
rect 307298 170992 307354 171048
rect 307114 170176 307170 170232
rect 307574 170584 307630 170640
rect 307666 169788 307722 169824
rect 307666 169768 307668 169788
rect 307668 169768 307720 169788
rect 307720 169768 307722 169788
rect 307482 169224 307538 169280
rect 307666 168816 307722 168872
rect 307574 168408 307630 168464
rect 307482 168000 307538 168056
rect 307666 167592 307722 167648
rect 307574 167184 307630 167240
rect 306746 166776 306802 166832
rect 307482 166368 307538 166424
rect 307390 165416 307446 165472
rect 307206 165008 307262 165064
rect 307114 162968 307170 163024
rect 307114 159568 307170 159624
rect 306746 159024 306802 159080
rect 306562 158208 306618 158264
rect 306562 155624 306618 155680
rect 306930 154400 306986 154456
rect 306746 153992 306802 154048
rect 306654 151816 306710 151872
rect 307114 152632 307170 152688
rect 306838 152224 306894 152280
rect 306562 145832 306618 145888
rect 307114 148416 307170 148472
rect 307022 148008 307078 148064
rect 306562 144608 306618 144664
rect 306562 142976 306618 143032
rect 306930 142024 306986 142080
rect 307022 141616 307078 141672
rect 306562 140392 306618 140448
rect 306562 139032 306618 139088
rect 306930 138624 306986 138680
rect 306562 136176 306618 136232
rect 307114 137400 307170 137456
rect 307114 135224 307170 135280
rect 307022 134000 307078 134056
rect 306930 133592 306986 133648
rect 306562 133184 306618 133240
rect 306930 128832 306986 128888
rect 306746 122032 306802 122088
rect 306562 119992 306618 120048
rect 305734 118904 305790 118960
rect 305826 117544 305882 117600
rect 306562 114416 306618 114472
rect 306746 111016 306802 111072
rect 306930 109792 306986 109848
rect 305918 107888 305974 107944
rect 306746 106800 306802 106856
rect 306746 105440 306802 105496
rect 306930 104216 306986 104272
rect 306746 103808 306802 103864
rect 306562 102448 306618 102504
rect 306562 102040 306618 102096
rect 307298 161608 307354 161664
rect 307298 160792 307354 160848
rect 307666 165824 307722 165880
rect 307574 164600 307630 164656
rect 307666 164228 307668 164248
rect 307668 164228 307720 164248
rect 307720 164228 307722 164248
rect 307666 164192 307722 164228
rect 307574 163784 307630 163840
rect 307666 163376 307722 163432
rect 307574 162424 307630 162480
rect 307666 162016 307722 162072
rect 307574 161200 307630 161256
rect 307666 160384 307722 160440
rect 307666 159976 307722 160032
rect 307574 158616 307630 158672
rect 307390 157800 307446 157856
rect 307666 157428 307668 157448
rect 307668 157428 307720 157448
rect 307720 157428 307722 157448
rect 307666 157392 307722 157428
rect 307482 156984 307538 157040
rect 307574 156576 307630 156632
rect 307666 156168 307722 156224
rect 307666 155216 307722 155272
rect 307482 154808 307538 154864
rect 307666 153584 307722 153640
rect 307666 153176 307722 153232
rect 307482 151408 307538 151464
rect 307666 151000 307722 151056
rect 307574 150592 307630 150648
rect 307574 150184 307630 150240
rect 307666 149232 307722 149288
rect 307390 148824 307446 148880
rect 307298 145424 307354 145480
rect 307482 147600 307538 147656
rect 307574 147192 307630 147248
rect 307666 146784 307722 146840
rect 307666 146396 307722 146432
rect 307666 146376 307668 146396
rect 307668 146376 307720 146396
rect 307720 146376 307722 146396
rect 307482 144200 307538 144256
rect 307666 143792 307722 143848
rect 307574 143384 307630 143440
rect 307666 142432 307722 142488
rect 307574 141208 307630 141264
rect 307666 140820 307722 140856
rect 307666 140800 307668 140820
rect 307668 140800 307720 140820
rect 307720 140800 307722 140820
rect 307666 139576 307722 139632
rect 307666 138216 307722 138272
rect 307666 137808 307722 137864
rect 307482 136584 307538 136640
rect 307666 135632 307722 135688
rect 307574 134816 307630 134872
rect 307666 134408 307722 134464
rect 307482 132232 307538 132288
rect 307574 131824 307630 131880
rect 307666 131416 307722 131472
rect 307482 131008 307538 131064
rect 307574 129920 307630 129976
rect 307666 129784 307722 129840
rect 307666 129240 307722 129296
rect 307482 128016 307538 128072
rect 307574 127608 307630 127664
rect 307666 127200 307722 127256
rect 307574 126792 307630 126848
rect 307666 125704 307722 125760
rect 307482 125432 307538 125488
rect 307574 125024 307630 125080
rect 307666 124616 307722 124672
rect 307666 124228 307722 124264
rect 307666 124208 307668 124228
rect 307668 124208 307720 124228
rect 307720 124208 307722 124228
rect 307574 123392 307630 123448
rect 307666 122984 307722 123040
rect 307574 122440 307630 122496
rect 307666 121624 307722 121680
rect 307298 121216 307354 121272
rect 307574 120808 307630 120864
rect 307666 120400 307722 120456
rect 307666 119584 307722 119640
rect 307574 118632 307630 118688
rect 307298 118224 307354 118280
rect 307666 117408 307722 117464
rect 307482 117000 307538 117056
rect 307574 116592 307630 116648
rect 307666 116184 307722 116240
rect 307298 115640 307354 115696
rect 307574 115232 307630 115288
rect 307666 114824 307722 114880
rect 307666 113212 307722 113248
rect 307666 113192 307668 113212
rect 307668 113192 307720 113212
rect 307720 113192 307722 113212
rect 307482 112648 307538 112704
rect 307574 112240 307630 112296
rect 307666 111832 307722 111888
rect 307298 111424 307354 111480
rect 307666 110608 307722 110664
rect 307574 110200 307630 110256
rect 307666 109248 307722 109304
rect 307482 108840 307538 108896
rect 307574 107752 307630 107808
rect 307666 107616 307722 107672
rect 307666 107208 307722 107264
rect 307482 106412 307538 106448
rect 307482 106392 307484 106412
rect 307484 106392 307536 106412
rect 307536 106392 307538 106412
rect 307574 105848 307630 105904
rect 307666 105032 307722 105088
rect 307482 104624 307538 104680
rect 307574 103400 307630 103456
rect 307666 102992 307722 103048
rect 307482 101632 307538 101688
rect 307574 101224 307630 101280
rect 307666 100816 307722 100872
rect 307482 100408 307538 100464
rect 307574 100000 307630 100056
rect 307666 99592 307722 99648
rect 307574 99048 307630 99104
rect 307298 98232 307354 98288
rect 307666 98640 307722 98696
rect 307206 97824 307262 97880
rect 307574 97416 307630 97472
rect 307390 97008 307446 97064
rect 307666 96600 307722 96656
rect 307666 96192 307722 96248
rect 337382 349696 337438 349752
rect 309322 114008 309378 114064
rect 309322 113056 309378 113112
rect 309138 101768 309194 101824
rect 313922 293936 313978 293992
rect 312634 177384 312690 177440
rect 318062 178608 318118 178664
rect 316038 176704 316094 176760
rect 318246 175888 318302 175944
rect 321466 175208 321522 175264
rect 321282 172624 321338 172680
rect 321558 141888 321614 141944
rect 321650 119856 321706 119912
rect 321834 170584 321890 170640
rect 322938 160112 322994 160168
rect 323030 137808 323086 137864
rect 324318 173984 324374 174040
rect 324318 173168 324374 173224
rect 324318 170856 324374 170912
rect 324502 168544 324558 168600
rect 324410 167728 324466 167784
rect 324318 167048 324374 167104
rect 324318 166232 324374 166288
rect 324318 165452 324320 165472
rect 324320 165452 324372 165472
rect 324372 165452 324374 165472
rect 324318 165416 324374 165452
rect 324410 164736 324466 164792
rect 324318 163920 324374 163976
rect 324410 163104 324466 163160
rect 324318 162424 324374 162480
rect 324410 161608 324466 161664
rect 324318 160792 324374 160848
rect 324318 159296 324374 159352
rect 324318 158480 324374 158536
rect 324410 157800 324466 157856
rect 324318 156984 324374 157040
rect 324318 156304 324374 156360
rect 324318 155488 324374 155544
rect 324410 154672 324466 154728
rect 324318 153992 324374 154048
rect 324410 153176 324466 153232
rect 324318 152360 324374 152416
rect 324318 151716 324320 151736
rect 324320 151716 324372 151736
rect 324372 151716 324374 151736
rect 324318 151680 324374 151716
rect 324410 150864 324466 150920
rect 324318 150048 324374 150104
rect 324318 149368 324374 149424
rect 324318 148552 324374 148608
rect 323214 147736 323270 147792
rect 324318 147056 324374 147112
rect 324318 146260 324374 146296
rect 324318 146240 324320 146260
rect 324320 146240 324372 146260
rect 324372 146240 324374 146260
rect 324410 145424 324466 145480
rect 324318 143928 324374 143984
rect 324318 143112 324374 143168
rect 325606 142432 325662 142488
rect 324318 140800 324374 140856
rect 324318 140120 324374 140176
rect 324318 139324 324374 139360
rect 324318 139304 324320 139324
rect 324320 139304 324372 139324
rect 324372 139304 324374 139324
rect 324410 138488 324466 138544
rect 324318 136992 324374 137048
rect 324318 136312 324374 136368
rect 325606 136040 325662 136096
rect 324318 133184 324374 133240
rect 324318 132388 324374 132424
rect 324318 132368 324320 132388
rect 324320 132368 324372 132388
rect 324372 132368 324374 132388
rect 324410 131688 324466 131744
rect 324318 130872 324374 130928
rect 324410 130056 324466 130112
rect 324318 129376 324374 129432
rect 324410 128560 324466 128616
rect 324318 127744 324374 127800
rect 324410 127064 324466 127120
rect 324318 125432 324374 125488
rect 324410 124752 324466 124808
rect 324318 123936 324374 123992
rect 324962 123120 325018 123176
rect 324318 122440 324374 122496
rect 323122 121624 323178 121680
rect 324318 120808 324374 120864
rect 324410 120128 324466 120184
rect 324318 118496 324374 118552
rect 324410 117816 324466 117872
rect 324318 116320 324374 116376
rect 324318 115504 324374 115560
rect 324410 114688 324466 114744
rect 321834 113600 321890 113656
rect 321742 104488 321798 104544
rect 321742 102176 321798 102232
rect 321650 101088 321706 101144
rect 321374 99592 321430 99648
rect 321466 97280 321522 97336
rect 321558 96600 321614 96656
rect 311898 90380 311900 90400
rect 311900 90380 311952 90400
rect 311952 90380 311954 90400
rect 311898 90344 311954 90380
rect 310518 77988 310574 78024
rect 310518 77968 310520 77988
rect 310520 77968 310572 77988
rect 310572 77968 310574 77988
rect 312634 11736 312690 11792
rect 311438 11600 311494 11656
rect 318890 43424 318946 43480
rect 320086 43460 320088 43480
rect 320088 43460 320140 43480
rect 320140 43460 320142 43480
rect 320086 43424 320142 43460
rect 324318 113192 324374 113248
rect 326066 178608 326122 178664
rect 326066 171264 326122 171320
rect 324318 112376 324374 112432
rect 322938 111696 322994 111752
rect 321926 102720 321982 102776
rect 324318 109384 324374 109440
rect 324318 108568 324374 108624
rect 325606 107752 325662 107808
rect 324318 105440 324374 105496
rect 323030 104760 323086 104816
rect 324410 100816 324466 100872
rect 332598 66816 332654 66872
rect 335542 175888 335598 175944
rect 334070 46180 334072 46200
rect 334072 46180 334124 46200
rect 334124 46180 334126 46200
rect 334070 46144 334126 46180
rect 342258 296792 342314 296848
rect 340878 295296 340934 295352
rect 335082 11736 335138 11792
rect 342350 87644 342406 87680
rect 342350 87624 342352 87644
rect 342352 87624 342404 87644
rect 342404 87624 342406 87644
rect 343362 11736 343418 11792
rect 340970 3440 341026 3496
rect 342074 3460 342130 3496
rect 342074 3440 342076 3460
rect 342076 3440 342128 3460
rect 342128 3440 342130 3460
rect 348422 174528 348478 174584
rect 416778 178608 416834 178664
rect 416778 176976 416834 177032
rect 416778 175208 416834 175264
rect 416778 171808 416834 171864
rect 416778 170176 416834 170232
rect 416778 165008 416834 165064
rect 416778 161744 416834 161800
rect 416778 159976 416834 160032
rect 416778 158344 416834 158400
rect 416778 156576 416834 156632
rect 416778 154944 416834 155000
rect 416778 153212 416780 153232
rect 416780 153212 416832 153232
rect 416832 153212 416834 153232
rect 416778 153176 416834 153212
rect 416778 151544 416834 151600
rect 416778 149776 416834 149832
rect 416778 148144 416834 148200
rect 416778 146512 416834 146568
rect 416778 144744 416834 144800
rect 416778 143112 416834 143168
rect 416778 141344 416834 141400
rect 416778 139712 416834 139768
rect 416778 137944 416834 138000
rect 416778 136312 416834 136368
rect 417330 134544 417386 134600
rect 416778 129512 416834 129568
rect 416778 119312 416834 119368
rect 416962 117680 417018 117736
rect 416778 114280 416834 114336
rect 416778 112648 416834 112704
rect 416778 110880 416834 110936
rect 417514 177248 417570 177304
rect 419170 134544 419226 134600
rect 417606 131280 417662 131336
rect 418526 126112 418582 126168
rect 418526 124480 418582 124536
rect 417514 121080 417570 121136
rect 417422 109248 417478 109304
rect 416778 107480 416834 107536
rect 416778 105848 416834 105904
rect 416778 104080 416834 104136
rect 416778 102448 416834 102504
rect 416778 100816 416834 100872
rect 419354 132912 419410 132968
rect 436098 292576 436154 292632
rect 455418 232464 455474 232520
rect 462318 225528 462374 225584
rect 491298 179288 491354 179344
rect 494150 170992 494206 171048
rect 419722 131280 419778 131336
rect 419538 122748 419540 122768
rect 419540 122748 419592 122768
rect 419592 122748 419594 122768
rect 419538 122712 419594 122748
rect 419814 127880 419870 127936
rect 373998 8880 374054 8936
rect 477498 67496 477554 67552
rect 494058 100000 494114 100056
rect 494242 132096 494298 132152
rect 494426 171672 494482 171728
rect 494334 131008 494390 131064
rect 495530 168816 495586 168872
rect 495438 132912 495494 132968
rect 495438 104896 495494 104952
rect 495438 102720 495494 102776
rect 495714 147600 495770 147656
rect 495622 121760 495678 121816
rect 496818 140800 496874 140856
rect 496818 139712 496874 139768
rect 496818 138624 496874 138680
rect 496818 137400 496874 137456
rect 496818 136312 496874 136368
rect 496818 134136 496874 134192
rect 497002 177792 497058 177848
rect 497002 176724 497058 176760
rect 497002 176704 497004 176724
rect 497004 176704 497056 176724
rect 497056 176704 497058 176724
rect 498106 175616 498162 175672
rect 497002 174392 497058 174448
rect 497002 169904 497058 169960
rect 497002 167728 497058 167784
rect 497002 166640 497058 166696
rect 497002 165416 497058 165472
rect 497094 164328 497150 164384
rect 497002 163240 497058 163296
rect 497002 162152 497058 162208
rect 497002 160928 497058 160984
rect 497002 159840 497058 159896
rect 497094 158752 497150 158808
rect 497002 157664 497058 157720
rect 497002 156440 497058 156496
rect 497002 155352 497058 155408
rect 497002 154264 497058 154320
rect 497094 153176 497150 153232
rect 497002 152088 497058 152144
rect 497002 150864 497058 150920
rect 497002 149776 497058 149832
rect 497002 148688 497058 148744
rect 497002 146376 497058 146432
rect 497002 145288 497058 145344
rect 497094 144200 497150 144256
rect 497002 143112 497058 143168
rect 497002 141888 497058 141944
rect 497002 135224 497058 135280
rect 496818 129684 496820 129704
rect 496820 129684 496872 129704
rect 496872 129684 496874 129704
rect 496818 129648 496874 129684
rect 496910 128424 496966 128480
rect 496818 126248 496874 126304
rect 496818 125160 496874 125216
rect 496818 124108 496820 124128
rect 496820 124108 496872 124128
rect 496872 124108 496874 124128
rect 496818 124072 496874 124108
rect 496910 122848 496966 122904
rect 496818 120672 496874 120728
rect 496818 119584 496874 119640
rect 496818 118360 496874 118416
rect 496910 117272 496966 117328
rect 497002 116184 497058 116240
rect 496818 115096 496874 115152
rect 496818 113872 496874 113928
rect 496818 112784 496874 112840
rect 496818 111716 496874 111752
rect 496818 111696 496820 111716
rect 496820 111696 496872 111716
rect 496872 111696 496874 111716
rect 496910 110608 496966 110664
rect 496818 109384 496874 109440
rect 497002 108296 497058 108352
rect 496818 106120 496874 106176
rect 496910 103808 496966 103864
rect 497094 107208 497150 107264
rect 495714 93744 495770 93800
rect 498382 101632 498438 101688
rect 503810 188264 503866 188320
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580906 670692 580908 670712
rect 580908 670692 580960 670712
rect 580960 670692 580962 670712
rect 580906 670656 580962 670692
rect 582378 670656 582434 670712
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 582392 580226 582448
rect 580170 577632 580226 577688
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 579802 524456 579858 524512
rect 580170 511264 580226 511320
rect 580354 490456 580410 490512
rect 580354 484608 580410 484664
rect 579894 471416 579950 471472
rect 579618 458088 579674 458144
rect 579802 431568 579858 431624
rect 579986 418240 580042 418296
rect 579618 404912 579674 404968
rect 580354 378392 580410 378448
rect 580262 365064 580318 365120
rect 579618 351872 579674 351928
rect 580262 325216 580318 325272
rect 580170 312024 580226 312080
rect 580906 298696 580962 298752
rect 579802 272176 579858 272232
rect 580170 258848 580226 258904
rect 579986 245520 580042 245576
rect 580262 232328 580318 232384
rect 580170 219000 580226 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 580262 179152 580318 179208
rect 580170 165824 580226 165880
rect 579802 152632 579858 152688
rect 580170 139304 580226 139360
rect 580170 125976 580226 126032
rect 580262 112784 580318 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580262 33088 580318 33144
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580901 670714 580967 670717
rect 582373 670714 582439 670717
rect 583520 670714 584960 670804
rect 580901 670712 584960 670714
rect 580901 670656 580906 670712
rect 580962 670656 582378 670712
rect 582434 670656 584960 670712
rect 580901 670654 584960 670656
rect 580901 670651 580967 670654
rect 582373 670651 582439 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 644058 584960 644148
rect 583342 643998 584960 644058
rect 583342 643922 583402 643998
rect 583520 643922 584960 643998
rect 583342 643908 584960 643922
rect 583342 643862 583586 643908
rect 111558 643180 111564 643244
rect 111628 643242 111634 643244
rect 583526 643242 583586 643862
rect 111628 643182 583586 643242
rect 111628 643180 111634 643182
rect -960 632090 480 632180
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 114502 586468 114508 586532
rect 114572 586468 114578 586532
rect 53598 586332 53604 586396
rect 53668 586394 53674 586396
rect 91645 586394 91711 586397
rect 53668 586392 91711 586394
rect 53668 586336 91650 586392
rect 91706 586336 91711 586392
rect 53668 586334 91711 586336
rect 53668 586332 53674 586334
rect 91645 586331 91711 586334
rect 94129 586394 94195 586397
rect 114510 586394 114570 586468
rect 94129 586392 114570 586394
rect 94129 586336 94134 586392
rect 94190 586336 114570 586392
rect 94129 586334 114570 586336
rect 94129 586331 94195 586334
rect 101397 584354 101463 584357
rect 111885 584354 111951 584357
rect 112069 584354 112135 584357
rect 101397 584352 112135 584354
rect 101397 584296 101402 584352
rect 101458 584296 111890 584352
rect 111946 584296 112074 584352
rect 112130 584296 112135 584352
rect 101397 584294 112135 584296
rect 101397 584291 101463 584294
rect 111885 584291 111951 584294
rect 112069 584291 112135 584294
rect 57646 583884 57652 583948
rect 57716 583946 57722 583948
rect 75085 583946 75151 583949
rect 57716 583944 75151 583946
rect 57716 583888 75090 583944
rect 75146 583888 75151 583944
rect 57716 583886 75151 583888
rect 57716 583884 57722 583886
rect 75085 583883 75151 583886
rect 82537 583946 82603 583949
rect 106917 583946 106983 583949
rect 82537 583944 106983 583946
rect 82537 583888 82542 583944
rect 82598 583888 106922 583944
rect 106978 583888 106983 583944
rect 82537 583886 106983 583888
rect 82537 583883 82603 583886
rect 106917 583883 106983 583886
rect 54937 583810 55003 583813
rect 81433 583810 81499 583813
rect 82077 583810 82143 583813
rect 54937 583808 82143 583810
rect 54937 583752 54942 583808
rect 54998 583752 81438 583808
rect 81494 583752 82082 583808
rect 82138 583752 82143 583808
rect 54937 583750 82143 583752
rect 54937 583747 55003 583750
rect 81433 583747 81499 583750
rect 82077 583747 82143 583750
rect 103881 583810 103947 583813
rect 121545 583810 121611 583813
rect 103881 583808 121611 583810
rect 103881 583752 103886 583808
rect 103942 583752 121550 583808
rect 121606 583752 121611 583808
rect 103881 583750 121611 583752
rect 103881 583747 103947 583750
rect 121545 583747 121611 583750
rect 69197 582450 69263 582453
rect 580165 582450 580231 582453
rect 69197 582448 580231 582450
rect 69197 582392 69202 582448
rect 69258 582392 580170 582448
rect 580226 582392 580231 582448
rect 69197 582390 580231 582392
rect 69197 582387 69263 582390
rect 580165 582387 580231 582390
rect 102593 581770 102659 581773
rect 109125 581770 109191 581773
rect 102593 581768 109191 581770
rect 102593 581712 102598 581768
rect 102654 581712 109130 581768
rect 109186 581712 109191 581768
rect 102593 581710 109191 581712
rect 102593 581707 102659 581710
rect 109125 581707 109191 581710
rect 67633 581362 67699 581365
rect 70166 581362 70226 581468
rect 67633 581360 70226 581362
rect 67633 581304 67638 581360
rect 67694 581304 70226 581360
rect 67633 581302 70226 581304
rect 67633 581299 67699 581302
rect 68645 580682 68711 580685
rect 70166 580682 70226 580788
rect 68645 580680 70226 580682
rect 68645 580624 68650 580680
rect 68706 580624 70226 580680
rect 68645 580622 70226 580624
rect 68645 580619 68711 580622
rect 105862 580546 105922 580788
rect 105862 580486 113190 580546
rect 108205 580138 108271 580141
rect 105892 580136 108271 580138
rect -960 580002 480 580092
rect 105892 580080 108210 580136
rect 108266 580080 108271 580136
rect 105892 580078 108271 580080
rect 108205 580075 108271 580078
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect 113130 580002 113190 580486
rect 117998 580002 118004 580004
rect 113130 579942 118004 580002
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 117998 579940 118004 579942
rect 118068 579940 118074 580004
rect 108849 579458 108915 579461
rect 105892 579456 108915 579458
rect 67725 579186 67791 579189
rect 70166 579186 70226 579428
rect 105892 579400 108854 579456
rect 108910 579400 108915 579456
rect 105892 579398 108915 579400
rect 108849 579395 108915 579398
rect 67725 579184 70226 579186
rect 67725 579128 67730 579184
rect 67786 579128 70226 579184
rect 67725 579126 70226 579128
rect 67725 579123 67791 579126
rect 108941 578778 109007 578781
rect 105892 578776 109007 578778
rect 67633 578506 67699 578509
rect 70166 578506 70226 578748
rect 105892 578720 108946 578776
rect 109002 578720 109007 578776
rect 105892 578718 109007 578720
rect 108941 578715 109007 578718
rect 67633 578504 70226 578506
rect 67633 578448 67638 578504
rect 67694 578448 70226 578504
rect 67633 578446 70226 578448
rect 67633 578443 67699 578446
rect 67633 577826 67699 577829
rect 70166 577826 70226 578068
rect 67633 577824 70226 577826
rect 67633 577768 67638 577824
rect 67694 577768 70226 577824
rect 67633 577766 70226 577768
rect 105862 577826 105922 578068
rect 106181 577826 106247 577829
rect 105862 577824 106247 577826
rect 105862 577768 106186 577824
rect 106242 577768 106247 577824
rect 105862 577766 106247 577768
rect 67633 577763 67699 577766
rect 106181 577763 106247 577766
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 108757 577418 108823 577421
rect 111742 577418 111748 577420
rect 105892 577416 111748 577418
rect 67541 577146 67607 577149
rect 70166 577146 70226 577388
rect 105892 577360 108762 577416
rect 108818 577360 111748 577416
rect 105892 577358 111748 577360
rect 108757 577355 108823 577358
rect 111742 577356 111748 577358
rect 111812 577356 111818 577420
rect 67541 577144 70226 577146
rect 67541 577088 67546 577144
rect 67602 577088 70226 577144
rect 67541 577086 70226 577088
rect 67541 577083 67607 577086
rect 107878 576738 107884 576740
rect 68645 576466 68711 576469
rect 70166 576466 70226 576708
rect 105892 576678 107884 576738
rect 107878 576676 107884 576678
rect 107948 576676 107954 576740
rect 68645 576464 70226 576466
rect 68645 576408 68650 576464
rect 68706 576408 70226 576464
rect 68645 576406 70226 576408
rect 68645 576403 68711 576406
rect 108941 576058 109007 576061
rect 105892 576056 109007 576058
rect 67633 575786 67699 575789
rect 70166 575786 70226 576028
rect 105892 576000 108946 576056
rect 109002 576000 109007 576056
rect 105892 575998 109007 576000
rect 108941 575995 109007 575998
rect 67633 575784 70226 575786
rect 67633 575728 67638 575784
rect 67694 575728 70226 575784
rect 67633 575726 70226 575728
rect 67633 575723 67699 575726
rect 67725 575106 67791 575109
rect 70166 575106 70226 575348
rect 67725 575104 70226 575106
rect 67725 575048 67730 575104
rect 67786 575048 70226 575104
rect 67725 575046 70226 575048
rect 67725 575043 67791 575046
rect 108941 574698 109007 574701
rect 105892 574696 109007 574698
rect 67633 574426 67699 574429
rect 70166 574426 70226 574668
rect 105892 574640 108946 574696
rect 109002 574640 109007 574696
rect 105892 574638 109007 574640
rect 108941 574635 109007 574638
rect 67633 574424 70226 574426
rect 67633 574368 67638 574424
rect 67694 574368 70226 574424
rect 67633 574366 70226 574368
rect 67633 574363 67699 574366
rect 108941 574018 109007 574021
rect 105892 574016 109007 574018
rect 67633 573474 67699 573477
rect 70166 573474 70226 573988
rect 105892 573960 108946 574016
rect 109002 573960 109007 574016
rect 105892 573958 109007 573960
rect 108941 573955 109007 573958
rect 67633 573472 70226 573474
rect 67633 573416 67638 573472
rect 67694 573416 70226 573472
rect 67633 573414 70226 573416
rect 67633 573411 67699 573414
rect 107653 573338 107719 573341
rect 108665 573338 108731 573341
rect 105892 573336 108731 573338
rect 105892 573280 107658 573336
rect 107714 573280 108670 573336
rect 108726 573280 108731 573336
rect 105892 573278 108731 573280
rect 107653 573275 107719 573278
rect 108665 573275 108731 573278
rect 67449 572794 67515 572797
rect 108941 572794 109007 572797
rect 67449 572792 70042 572794
rect 67449 572736 67454 572792
rect 67510 572736 70042 572792
rect 105892 572792 109007 572794
rect 67449 572734 70042 572736
rect 67449 572731 67515 572734
rect 69982 572730 70042 572734
rect 70166 572730 70226 572764
rect 105892 572736 108946 572792
rect 109002 572736 109007 572792
rect 105892 572734 109007 572736
rect 108941 572731 109007 572734
rect 121678 572732 121684 572796
rect 121748 572794 121754 572796
rect 122097 572794 122163 572797
rect 121748 572792 122163 572794
rect 121748 572736 122102 572792
rect 122158 572736 122163 572792
rect 121748 572734 122163 572736
rect 121748 572732 121754 572734
rect 122097 572731 122163 572734
rect 69982 572670 70226 572730
rect 68921 572522 68987 572525
rect 68921 572520 70226 572522
rect 68921 572464 68926 572520
rect 68982 572464 70226 572520
rect 68921 572462 70226 572464
rect 68921 572459 68987 572462
rect 70166 572084 70226 572462
rect 108941 571978 109007 571981
rect 105892 571976 109007 571978
rect 105892 571920 108946 571976
rect 109002 571920 109007 571976
rect 105892 571918 109007 571920
rect 108941 571915 109007 571918
rect 66478 571780 66484 571844
rect 66548 571842 66554 571844
rect 68921 571842 68987 571845
rect 66548 571840 68987 571842
rect 66548 571784 68926 571840
rect 68982 571784 68987 571840
rect 66548 571782 68987 571784
rect 66548 571780 66554 571782
rect 68921 571779 68987 571782
rect 68277 571706 68343 571709
rect 68461 571706 68527 571709
rect 68277 571704 70410 571706
rect 68277 571648 68282 571704
rect 68338 571648 68466 571704
rect 68522 571648 70410 571704
rect 68277 571646 70410 571648
rect 68277 571643 68343 571646
rect 68461 571643 68527 571646
rect 70350 571404 70410 571646
rect 105494 571164 105554 571268
rect 105486 571100 105492 571164
rect 105556 571100 105562 571164
rect 65926 570284 65932 570348
rect 65996 570346 66002 570348
rect 70166 570346 70226 570588
rect 65996 570286 70226 570346
rect 105862 570346 105922 570588
rect 129774 570346 129780 570348
rect 105862 570286 129780 570346
rect 65996 570284 66002 570286
rect 129774 570284 129780 570286
rect 129844 570284 129850 570348
rect 67633 570074 67699 570077
rect 108941 570074 109007 570077
rect 67633 570072 70042 570074
rect 67633 570016 67638 570072
rect 67694 570016 70042 570072
rect 67633 570014 70042 570016
rect 105892 570072 109007 570074
rect 105892 570016 108946 570072
rect 109002 570016 109007 570072
rect 105892 570014 109007 570016
rect 67633 570011 67699 570014
rect 69982 569802 70042 570014
rect 108941 570011 109007 570014
rect 70166 569802 70226 569908
rect 69982 569742 70226 569802
rect 107653 569258 107719 569261
rect 105892 569256 107719 569258
rect 66110 568924 66116 568988
rect 66180 568986 66186 568988
rect 70166 568986 70226 569228
rect 105892 569200 107658 569256
rect 107714 569200 107719 569256
rect 105892 569198 107719 569200
rect 107653 569195 107719 569198
rect 66180 568926 70226 568986
rect 66180 568924 66186 568926
rect 67633 568714 67699 568717
rect 67633 568712 70042 568714
rect 67633 568656 67638 568712
rect 67694 568656 70042 568712
rect 67633 568654 70042 568656
rect 67633 568651 67699 568654
rect 69982 568442 70042 568654
rect 70166 568442 70226 568548
rect 69982 568382 70226 568442
rect 108941 567898 109007 567901
rect 105892 567896 109007 567898
rect 67725 567626 67791 567629
rect 70166 567626 70226 567868
rect 105892 567840 108946 567896
rect 109002 567840 109007 567896
rect 105892 567838 109007 567840
rect 108941 567835 109007 567838
rect 67725 567624 70226 567626
rect 67725 567568 67730 567624
rect 67786 567568 70226 567624
rect 67725 567566 70226 567568
rect 67725 567563 67791 567566
rect 67633 567218 67699 567221
rect 108941 567218 109007 567221
rect 67633 567216 70042 567218
rect 67633 567160 67638 567216
rect 67694 567210 70042 567216
rect 105892 567216 109007 567218
rect 67694 567160 70226 567210
rect 67633 567158 70226 567160
rect 105892 567160 108946 567216
rect 109002 567160 109007 567216
rect 105892 567158 109007 567160
rect 67633 567155 67699 567158
rect 69982 567150 70226 567158
rect 108941 567155 109007 567158
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 108849 566538 108915 566541
rect 105892 566536 108915 566538
rect 105892 566480 108854 566536
rect 108910 566480 108915 566536
rect 105892 566478 108915 566480
rect 108849 566475 108915 566478
rect 67633 566266 67699 566269
rect 67633 566264 70410 566266
rect 67633 566208 67638 566264
rect 67694 566208 70410 566264
rect 67633 566206 70410 566208
rect 67633 566203 67699 566206
rect 70350 565964 70410 566206
rect 108941 565858 109007 565861
rect 105892 565856 109007 565858
rect 105892 565800 108946 565856
rect 109002 565800 109007 565856
rect 105892 565798 109007 565800
rect 108941 565795 109007 565798
rect 108849 565178 108915 565181
rect 105892 565176 108915 565178
rect 67633 564906 67699 564909
rect 70166 564906 70226 565148
rect 105892 565120 108854 565176
rect 108910 565120 108915 565176
rect 105892 565118 108915 565120
rect 108849 565115 108915 565118
rect 67633 564904 70226 564906
rect 67633 564848 67638 564904
rect 67694 564848 70226 564904
rect 67633 564846 70226 564848
rect 67633 564843 67699 564846
rect 67357 564498 67423 564501
rect 106365 564498 106431 564501
rect 67357 564496 70042 564498
rect 67357 564440 67362 564496
rect 67418 564440 70042 564496
rect 105892 564496 106431 564498
rect 67357 564438 70042 564440
rect 67357 564435 67423 564438
rect 69982 564362 70042 564438
rect 70166 564362 70226 564468
rect 105892 564440 106370 564496
rect 106426 564440 106431 564496
rect 105892 564438 106431 564440
rect 106365 564435 106431 564438
rect 69982 564302 70226 564362
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 108941 563954 109007 563957
rect 105892 563952 109007 563954
rect 105892 563896 108946 563952
rect 109002 563896 109007 563952
rect 105892 563894 109007 563896
rect 108941 563891 109007 563894
rect 67725 563546 67791 563549
rect 70166 563546 70226 563788
rect 67725 563544 70226 563546
rect 67725 563488 67730 563544
rect 67786 563488 70226 563544
rect 67725 563486 70226 563488
rect 67725 563483 67791 563486
rect 67633 563138 67699 563141
rect 107694 563138 107700 563140
rect 67633 563136 70042 563138
rect 67633 563080 67638 563136
rect 67694 563080 70042 563136
rect 67633 563078 70042 563080
rect 67633 563075 67699 563078
rect 69982 563002 70042 563078
rect 70166 563002 70226 563108
rect 105892 563078 107700 563138
rect 107694 563076 107700 563078
rect 107764 563076 107770 563140
rect 69982 562942 70226 563002
rect 108941 562458 109007 562461
rect 105892 562456 109007 562458
rect 67633 562322 67699 562325
rect 70166 562322 70226 562428
rect 105892 562400 108946 562456
rect 109002 562400 109007 562456
rect 105892 562398 109007 562400
rect 108941 562395 109007 562398
rect 67633 562320 70226 562322
rect 67633 562264 67638 562320
rect 67694 562264 70226 562320
rect 67633 562262 70226 562264
rect 67633 562259 67699 562262
rect 67633 562186 67699 562189
rect 67633 562184 70410 562186
rect 67633 562128 67638 562184
rect 67694 562128 70410 562184
rect 67633 562126 70410 562128
rect 67633 562123 67699 562126
rect 70350 561884 70410 562126
rect 108941 561098 109007 561101
rect 105892 561096 109007 561098
rect 67725 560826 67791 560829
rect 70166 560826 70226 561068
rect 105892 561040 108946 561096
rect 109002 561040 109007 561096
rect 105892 561038 109007 561040
rect 108941 561035 109007 561038
rect 67725 560824 70226 560826
rect 67725 560768 67730 560824
rect 67786 560768 70226 560824
rect 67725 560766 70226 560768
rect 67725 560763 67791 560766
rect 67633 560418 67699 560421
rect 106273 560418 106339 560421
rect 107653 560418 107719 560421
rect 67633 560416 70042 560418
rect 67633 560360 67638 560416
rect 67694 560360 70042 560416
rect 105892 560416 107719 560418
rect 67633 560358 70042 560360
rect 67633 560355 67699 560358
rect 69982 560282 70042 560358
rect 70166 560282 70226 560388
rect 105892 560360 106278 560416
rect 106334 560360 107658 560416
rect 107714 560360 107719 560416
rect 105892 560358 107719 560360
rect 106273 560355 106339 560358
rect 107653 560355 107719 560358
rect 69982 560222 70226 560282
rect 108849 559738 108915 559741
rect 105892 559736 108915 559738
rect 105892 559680 108854 559736
rect 108910 559680 108915 559736
rect 105892 559678 108915 559680
rect 108849 559675 108915 559678
rect 67633 559466 67699 559469
rect 67633 559464 70410 559466
rect 67633 559408 67638 559464
rect 67694 559408 70410 559464
rect 67633 559406 70410 559408
rect 67633 559403 67699 559406
rect 70350 559164 70410 559406
rect 108941 559058 109007 559061
rect 105892 559056 109007 559058
rect 105892 559000 108946 559056
rect 109002 559000 109007 559056
rect 105892 558998 109007 559000
rect 108941 558995 109007 558998
rect 68829 558922 68895 558925
rect 68829 558920 70226 558922
rect 68829 558864 68834 558920
rect 68890 558864 70226 558920
rect 68829 558862 70226 558864
rect 68829 558859 68895 558862
rect 70166 558484 70226 558862
rect 108941 558378 109007 558381
rect 105892 558376 109007 558378
rect 105892 558320 108946 558376
rect 109002 558320 109007 558376
rect 105892 558318 109007 558320
rect 108941 558315 109007 558318
rect 107745 557698 107811 557701
rect 105892 557696 107811 557698
rect 67633 557562 67699 557565
rect 70166 557562 70226 557668
rect 105892 557640 107750 557696
rect 107806 557640 107811 557696
rect 105892 557638 107811 557640
rect 107745 557635 107811 557638
rect 67633 557560 70226 557562
rect 67633 557504 67638 557560
rect 67694 557504 70226 557560
rect 67633 557502 70226 557504
rect 67633 557499 67699 557502
rect 68277 557426 68343 557429
rect 69974 557426 69980 557428
rect 68277 557424 69980 557426
rect 68277 557368 68282 557424
rect 68338 557368 69980 557424
rect 68277 557366 69980 557368
rect 68277 557363 68343 557366
rect 69974 557364 69980 557366
rect 70044 557364 70050 557428
rect 108941 557018 109007 557021
rect 105892 557016 109007 557018
rect 67725 556746 67791 556749
rect 70166 556746 70226 556988
rect 105892 556960 108946 557016
rect 109002 556960 109007 557016
rect 105892 556958 109007 556960
rect 108941 556955 109007 556958
rect 67725 556744 70226 556746
rect 67725 556688 67730 556744
rect 67786 556688 70226 556744
rect 67725 556686 70226 556688
rect 67725 556683 67791 556686
rect 107929 556338 107995 556341
rect 105892 556336 107995 556338
rect 67633 556202 67699 556205
rect 70166 556202 70226 556308
rect 105892 556280 107934 556336
rect 107990 556280 107995 556336
rect 105892 556278 107995 556280
rect 107929 556275 107995 556278
rect 67633 556200 70226 556202
rect 67633 556144 67638 556200
rect 67694 556144 70226 556200
rect 67633 556142 70226 556144
rect 67633 556139 67699 556142
rect 108849 555794 108915 555797
rect 105892 555792 108915 555794
rect 105892 555736 108854 555792
rect 108910 555736 108915 555792
rect 105892 555734 108915 555736
rect 108849 555731 108915 555734
rect 67725 555386 67791 555389
rect 70166 555386 70226 555628
rect 67725 555384 70226 555386
rect 67725 555328 67730 555384
rect 67786 555328 70226 555384
rect 67725 555326 70226 555328
rect 67725 555323 67791 555326
rect 67633 554842 67699 554845
rect 70166 554842 70226 554948
rect 67633 554840 70226 554842
rect 67633 554784 67638 554840
rect 67694 554784 70226 554840
rect 67633 554782 70226 554784
rect 67633 554779 67699 554782
rect 108941 554298 109007 554301
rect 105892 554296 109007 554298
rect -960 553890 480 553980
rect 68870 553964 68876 554028
rect 68940 554026 68946 554028
rect 70166 554026 70226 554268
rect 105892 554240 108946 554296
rect 109002 554240 109007 554296
rect 105892 554238 109007 554240
rect 108941 554235 109007 554238
rect 111558 554026 111564 554028
rect 68940 553966 70226 554026
rect 105862 553966 111564 554026
rect 68940 553964 68946 553966
rect 3509 553890 3575 553893
rect -960 553888 3575 553890
rect -960 553832 3514 553888
rect 3570 553832 3575 553888
rect -960 553830 3575 553832
rect -960 553740 480 553830
rect 3509 553827 3575 553830
rect 105862 553724 105922 553966
rect 111558 553964 111564 553966
rect 111628 554026 111634 554028
rect 124397 554026 124463 554029
rect 111628 554024 124463 554026
rect 111628 553968 124402 554024
rect 124458 553968 124463 554024
rect 111628 553966 124463 553968
rect 111628 553964 111634 553966
rect 124397 553963 124463 553966
rect 67633 553482 67699 553485
rect 70166 553482 70226 553588
rect 67633 553480 70226 553482
rect 67633 553424 67638 553480
rect 67694 553424 70226 553480
rect 67633 553422 70226 553424
rect 67633 553419 67699 553422
rect 108941 552938 109007 552941
rect 105892 552936 109007 552938
rect 105892 552880 108946 552936
rect 109002 552880 109007 552936
rect 105892 552878 109007 552880
rect 108941 552875 109007 552878
rect 107009 552258 107075 552261
rect 105892 552256 107075 552258
rect 67633 552122 67699 552125
rect 70166 552122 70226 552228
rect 105892 552200 107014 552256
rect 107070 552200 107075 552256
rect 105892 552198 107075 552200
rect 107009 552195 107075 552198
rect 67633 552120 70226 552122
rect 67633 552064 67638 552120
rect 67694 552064 70226 552120
rect 67633 552062 70226 552064
rect 67633 552059 67699 552062
rect 107653 551578 107719 551581
rect 105892 551576 107719 551578
rect 67633 551306 67699 551309
rect 70166 551306 70226 551548
rect 105892 551520 107658 551576
rect 107714 551520 107719 551576
rect 105892 551518 107719 551520
rect 107653 551515 107719 551518
rect 67633 551304 70226 551306
rect 67633 551248 67638 551304
rect 67694 551248 70226 551304
rect 67633 551246 70226 551248
rect 67633 551243 67699 551246
rect 583520 551020 584960 551260
rect 108941 550898 109007 550901
rect 105892 550896 109007 550898
rect 68829 550762 68895 550765
rect 70166 550762 70226 550868
rect 105892 550840 108946 550896
rect 109002 550840 109007 550896
rect 105892 550838 109007 550840
rect 108941 550835 109007 550838
rect 68829 550760 70226 550762
rect 68829 550704 68834 550760
rect 68890 550704 70226 550760
rect 68829 550702 70226 550704
rect 68829 550699 68895 550702
rect 108849 550218 108915 550221
rect 105892 550216 108915 550218
rect 67633 549946 67699 549949
rect 70166 549946 70226 550188
rect 105892 550160 108854 550216
rect 108910 550160 108915 550216
rect 105892 550158 108915 550160
rect 108849 550155 108915 550158
rect 67633 549944 70226 549946
rect 67633 549888 67638 549944
rect 67694 549888 70226 549944
rect 67633 549886 70226 549888
rect 67633 549883 67699 549886
rect 61878 549476 61884 549540
rect 61948 549538 61954 549540
rect 108941 549538 109007 549541
rect 61948 549478 64890 549538
rect 105892 549536 109007 549538
rect 61948 549476 61954 549478
rect 64830 549402 64890 549478
rect 70166 549402 70226 549508
rect 105892 549480 108946 549536
rect 109002 549480 109007 549536
rect 105892 549478 109007 549480
rect 108941 549475 109007 549478
rect 64830 549342 70226 549402
rect 67725 548586 67791 548589
rect 70166 548586 70226 548828
rect 67725 548584 70226 548586
rect 67725 548528 67730 548584
rect 67786 548528 70226 548584
rect 67725 548526 70226 548528
rect 67725 548523 67791 548526
rect 105678 548453 105738 548828
rect 105678 548448 105787 548453
rect 105678 548392 105726 548448
rect 105782 548392 105787 548448
rect 105678 548390 105787 548392
rect 105721 548387 105787 548390
rect 67633 548042 67699 548045
rect 70166 548042 70226 548148
rect 67633 548040 70226 548042
rect 67633 547984 67638 548040
rect 67694 547984 70226 548040
rect 67633 547982 70226 547984
rect 67633 547979 67699 547982
rect 108941 547498 109007 547501
rect 105892 547496 109007 547498
rect 67725 547226 67791 547229
rect 70166 547226 70226 547468
rect 105892 547440 108946 547496
rect 109002 547440 109007 547496
rect 105892 547438 109007 547440
rect 108941 547435 109007 547438
rect 67725 547224 70226 547226
rect 67725 547168 67730 547224
rect 67786 547168 70226 547224
rect 67725 547166 70226 547168
rect 67725 547163 67791 547166
rect 107653 546818 107719 546821
rect 105892 546816 107719 546818
rect 67633 546546 67699 546549
rect 70166 546546 70226 546788
rect 105892 546760 107658 546816
rect 107714 546760 107719 546816
rect 105892 546758 107719 546760
rect 107653 546755 107719 546758
rect 67633 546544 70226 546546
rect 67633 546488 67638 546544
rect 67694 546488 70226 546544
rect 67633 546486 70226 546488
rect 67633 546483 67699 546486
rect 108941 546138 109007 546141
rect 105892 546136 109007 546138
rect 105892 546080 108946 546136
rect 109002 546080 109007 546136
rect 105892 546078 109007 546080
rect 108941 546075 109007 546078
rect 112345 545730 112411 545733
rect 113081 545730 113147 545733
rect 125726 545730 125732 545732
rect 112345 545728 125732 545730
rect 112345 545672 112350 545728
rect 112406 545672 113086 545728
rect 113142 545672 125732 545728
rect 112345 545670 125732 545672
rect 112345 545667 112411 545670
rect 113081 545667 113147 545670
rect 125726 545668 125732 545670
rect 125796 545668 125802 545732
rect 108941 545458 109007 545461
rect 105892 545456 109007 545458
rect 68093 545322 68159 545325
rect 69197 545322 69263 545325
rect 70166 545322 70226 545428
rect 105892 545400 108946 545456
rect 109002 545400 109007 545456
rect 105892 545398 109007 545400
rect 108941 545395 109007 545398
rect 68093 545320 70226 545322
rect 68093 545264 68098 545320
rect 68154 545264 69202 545320
rect 69258 545264 70226 545320
rect 68093 545262 70226 545264
rect 68093 545259 68159 545262
rect 69197 545259 69263 545262
rect 108941 544778 109007 544781
rect 105892 544776 109007 544778
rect 68737 544506 68803 544509
rect 70166 544506 70226 544748
rect 105892 544720 108946 544776
rect 109002 544720 109007 544776
rect 105892 544718 109007 544720
rect 108941 544715 109007 544718
rect 68737 544504 70226 544506
rect 68737 544448 68742 544504
rect 68798 544448 70226 544504
rect 68737 544446 70226 544448
rect 68737 544443 68803 544446
rect 108941 544098 109007 544101
rect 105892 544096 109007 544098
rect 68001 543962 68067 543965
rect 68921 543962 68987 543965
rect 70166 543962 70226 544068
rect 105892 544040 108946 544096
rect 109002 544040 109007 544096
rect 105892 544038 109007 544040
rect 108941 544035 109007 544038
rect 68001 543960 70226 543962
rect 68001 543904 68006 543960
rect 68062 543904 68926 543960
rect 68982 543904 70226 543960
rect 68001 543902 70226 543904
rect 68001 543899 68067 543902
rect 68921 543899 68987 543902
rect 107837 543418 107903 543421
rect 105892 543416 107903 543418
rect 68001 543282 68067 543285
rect 69013 543282 69079 543285
rect 70166 543282 70226 543388
rect 105892 543360 107842 543416
rect 107898 543360 107903 543416
rect 105892 543358 107903 543360
rect 107837 543355 107903 543358
rect 68001 543280 70226 543282
rect 68001 543224 68006 543280
rect 68062 543224 69018 543280
rect 69074 543224 70226 543280
rect 68001 543222 70226 543224
rect 68001 543219 68067 543222
rect 69013 543219 69079 543222
rect 67633 542602 67699 542605
rect 70166 542602 70226 542708
rect 67633 542600 70226 542602
rect 67633 542544 67638 542600
rect 67694 542544 70226 542600
rect 67633 542542 70226 542544
rect 67633 542539 67699 542542
rect 105862 542466 105922 542708
rect 105862 542406 107762 542466
rect 107702 542330 107762 542406
rect 107837 542330 107903 542333
rect 107702 542328 107903 542330
rect 107702 542272 107842 542328
rect 107898 542272 107903 542328
rect 107702 542270 107903 542272
rect 107837 542267 107903 542270
rect 106917 542058 106983 542061
rect 105892 542056 106983 542058
rect 69197 541786 69263 541789
rect 70166 541786 70226 542028
rect 105892 542000 106922 542056
rect 106978 542000 106983 542056
rect 105892 541998 106983 542000
rect 106917 541995 106983 541998
rect 69197 541784 70226 541786
rect 69197 541728 69202 541784
rect 69258 541728 70226 541784
rect 69197 541726 70226 541728
rect 69197 541723 69263 541726
rect 124949 541650 125015 541653
rect 299473 541650 299539 541653
rect 122790 541648 299539 541650
rect 122790 541592 124954 541648
rect 125010 541592 299478 541648
rect 299534 541592 299539 541648
rect 122790 541590 299539 541592
rect 67633 541242 67699 541245
rect 70166 541242 70226 541348
rect 67633 541240 70226 541242
rect 67633 541184 67638 541240
rect 67694 541184 70226 541240
rect 67633 541182 70226 541184
rect 67633 541179 67699 541182
rect 109534 541044 109540 541108
rect 109604 541106 109610 541108
rect 122790 541106 122850 541590
rect 124949 541587 125015 541590
rect 299473 541587 299539 541590
rect 109604 541046 122850 541106
rect 109604 541044 109610 541046
rect -960 540684 480 540924
rect 106457 540698 106523 540701
rect 106825 540698 106891 540701
rect 105892 540696 106891 540698
rect 67633 540154 67699 540157
rect 70166 540154 70226 540668
rect 105892 540640 106462 540696
rect 106518 540640 106830 540696
rect 106886 540640 106891 540696
rect 105892 540638 106891 540640
rect 106457 540635 106523 540638
rect 106825 540635 106891 540638
rect 67633 540152 70226 540154
rect 67633 540096 67638 540152
rect 67694 540096 70226 540152
rect 67633 540094 70226 540096
rect 67633 540091 67699 540094
rect 107510 540018 107516 540020
rect 105892 539958 107516 540018
rect 107510 539956 107516 539958
rect 107580 540018 107586 540020
rect 108297 540018 108363 540021
rect 107580 540016 108363 540018
rect 107580 539960 108302 540016
rect 108358 539960 108363 540016
rect 107580 539958 108363 539960
rect 107580 539956 107586 539958
rect 108297 539955 108363 539958
rect 88057 538114 88123 538117
rect 88057 538112 99390 538114
rect 88057 538056 88062 538112
rect 88118 538056 99390 538112
rect 88057 538054 99390 538056
rect 88057 538051 88123 538054
rect 99330 537842 99390 538054
rect 103646 538052 103652 538116
rect 103716 538114 103722 538116
rect 104801 538114 104867 538117
rect 103716 538112 104867 538114
rect 103716 538056 104806 538112
rect 104862 538056 104867 538112
rect 103716 538054 104867 538056
rect 103716 538052 103722 538054
rect 104801 538051 104867 538054
rect 103513 537978 103579 537981
rect 109534 537978 109540 537980
rect 103513 537976 109540 537978
rect 103513 537920 103518 537976
rect 103574 537920 109540 537976
rect 103513 537918 109540 537920
rect 103513 537915 103579 537918
rect 109534 537916 109540 537918
rect 109604 537916 109610 537980
rect 109677 537842 109743 537845
rect 99330 537840 109743 537842
rect 99330 537784 109682 537840
rect 109738 537784 109743 537840
rect 99330 537782 109743 537784
rect 109677 537779 109743 537782
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 59118 537508 59124 537572
rect 59188 537570 59194 537572
rect 80329 537570 80395 537573
rect 59188 537568 80395 537570
rect 59188 537512 80334 537568
rect 80390 537512 80395 537568
rect 59188 537510 80395 537512
rect 59188 537508 59194 537510
rect 80329 537507 80395 537510
rect 57830 537372 57836 537436
rect 57900 537434 57906 537436
rect 81617 537434 81683 537437
rect 57900 537432 81683 537434
rect 57900 537376 81622 537432
rect 81678 537376 81683 537432
rect 57900 537374 81683 537376
rect 57900 537372 57906 537374
rect 81617 537371 81683 537374
rect 100937 537434 101003 537437
rect 101254 537434 101260 537436
rect 100937 537432 101260 537434
rect 100937 537376 100942 537432
rect 100998 537376 101260 537432
rect 100937 537374 101260 537376
rect 100937 537371 101003 537374
rect 101254 537372 101260 537374
rect 101324 537372 101330 537436
rect 53598 536012 53604 536076
rect 53668 536074 53674 536076
rect 87137 536074 87203 536077
rect 53668 536072 87203 536074
rect 53668 536016 87142 536072
rect 87198 536016 87203 536072
rect 53668 536014 87203 536016
rect 53668 536012 53674 536014
rect 87137 536011 87203 536014
rect 99741 535394 99807 535397
rect 107878 535394 107884 535396
rect 99741 535392 107884 535394
rect 99741 535336 99746 535392
rect 99802 535336 107884 535392
rect 99741 535334 107884 535336
rect 99741 535331 99807 535334
rect 107878 535332 107884 535334
rect 107948 535332 107954 535396
rect 92565 534714 92631 534717
rect 108798 534714 108804 534716
rect 92565 534712 108804 534714
rect 92565 534656 92570 534712
rect 92626 534656 108804 534712
rect 92565 534654 108804 534656
rect 92565 534651 92631 534654
rect 108798 534652 108804 534654
rect 108868 534652 108874 534716
rect 44030 529076 44036 529140
rect 44100 529138 44106 529140
rect 74533 529138 74599 529141
rect 44100 529136 74599 529138
rect 44100 529080 74538 529136
rect 74594 529080 74599 529136
rect 44100 529078 74599 529080
rect 44100 529076 44106 529078
rect 74533 529075 74599 529078
rect -960 527914 480 528004
rect 3141 527914 3207 527917
rect -960 527912 3207 527914
rect -960 527856 3146 527912
rect 3202 527856 3207 527912
rect -960 527854 3207 527856
rect -960 527764 480 527854
rect 3141 527851 3207 527854
rect 38561 525874 38627 525877
rect 38561 525872 64890 525874
rect 38561 525816 38566 525872
rect 38622 525816 64890 525872
rect 38561 525814 64890 525816
rect 38561 525811 38627 525814
rect 64830 525738 64890 525814
rect 69197 525738 69263 525741
rect 64830 525736 69263 525738
rect 64830 525680 69202 525736
rect 69258 525680 69263 525736
rect 64830 525678 69263 525680
rect 69197 525675 69263 525678
rect 579797 524514 579863 524517
rect 583520 524514 584960 524604
rect 579797 524512 584960 524514
rect 579797 524456 579802 524512
rect 579858 524456 584960 524512
rect 579797 524454 584960 524456
rect 579797 524451 579863 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3417 501802 3483 501805
rect -960 501800 3483 501802
rect -960 501744 3422 501800
rect 3478 501744 3483 501800
rect -960 501742 3483 501744
rect -960 501652 480 501742
rect 3417 501739 3483 501742
rect 114502 500380 114508 500444
rect 114572 500442 114578 500444
rect 114829 500442 114895 500445
rect 114572 500440 114895 500442
rect 114572 500384 114834 500440
rect 114890 500384 114895 500440
rect 114572 500382 114895 500384
rect 114572 500380 114578 500382
rect 114829 500379 114895 500382
rect 97717 500306 97783 500309
rect 114502 500306 114508 500308
rect 97717 500304 114508 500306
rect 97717 500248 97722 500304
rect 97778 500248 114508 500304
rect 97717 500246 114508 500248
rect 97717 500243 97783 500246
rect 114502 500244 114508 500246
rect 114572 500244 114578 500308
rect 87413 500170 87479 500173
rect 111926 500170 111932 500172
rect 87413 500168 111932 500170
rect 87413 500112 87418 500168
rect 87474 500112 111932 500168
rect 87413 500110 111932 500112
rect 87413 500107 87479 500110
rect 111926 500108 111932 500110
rect 111996 500108 112002 500172
rect 80605 499626 80671 499629
rect 110638 499626 110644 499628
rect 80605 499624 110644 499626
rect 80605 499568 80610 499624
rect 80666 499568 110644 499624
rect 80605 499566 110644 499568
rect 80605 499563 80671 499566
rect 110638 499564 110644 499566
rect 110708 499564 110714 499628
rect 128445 498810 128511 498813
rect 136582 498810 136588 498812
rect 128445 498808 136588 498810
rect 128445 498752 128450 498808
rect 128506 498752 136588 498808
rect 128445 498750 136588 498752
rect 128445 498747 128511 498750
rect 136582 498748 136588 498750
rect 136652 498748 136658 498812
rect 583520 497844 584960 498084
rect 60590 494668 60596 494732
rect 60660 494730 60666 494732
rect 84193 494730 84259 494733
rect 60660 494728 84259 494730
rect 60660 494672 84198 494728
rect 84254 494672 84259 494728
rect 60660 494670 84259 494672
rect 60660 494668 60666 494670
rect 84193 494667 84259 494670
rect 52310 493308 52316 493372
rect 52380 493370 52386 493372
rect 54109 493370 54175 493373
rect 52380 493368 54175 493370
rect 52380 493312 54114 493368
rect 54170 493312 54175 493368
rect 52380 493310 54175 493312
rect 52380 493308 52386 493310
rect 54109 493307 54175 493310
rect 50286 492628 50292 492692
rect 50356 492690 50362 492692
rect 50705 492690 50771 492693
rect 50356 492688 50771 492690
rect 50356 492632 50710 492688
rect 50766 492632 50771 492688
rect 50356 492630 50771 492632
rect 50356 492628 50362 492630
rect 50705 492627 50771 492630
rect 48078 491812 48084 491876
rect 48148 491874 48154 491876
rect 71773 491874 71839 491877
rect 48148 491872 71839 491874
rect 48148 491816 71778 491872
rect 71834 491816 71839 491872
rect 48148 491814 71839 491816
rect 48148 491812 48154 491814
rect 71773 491811 71839 491814
rect 99281 491874 99347 491877
rect 111006 491874 111012 491876
rect 99281 491872 111012 491874
rect 99281 491816 99286 491872
rect 99342 491816 111012 491872
rect 99281 491814 111012 491816
rect 99281 491811 99347 491814
rect 111006 491812 111012 491814
rect 111076 491812 111082 491876
rect 82261 491602 82327 491605
rect 109309 491602 109375 491605
rect 82261 491600 109375 491602
rect 82261 491544 82266 491600
rect 82322 491544 109314 491600
rect 109370 491544 109375 491600
rect 82261 491542 109375 491544
rect 82261 491539 82327 491542
rect 109309 491539 109375 491542
rect 96429 491466 96495 491469
rect 102041 491466 102107 491469
rect 96429 491464 102107 491466
rect 96429 491408 96434 491464
rect 96490 491408 102046 491464
rect 102102 491408 102107 491464
rect 96429 491406 102107 491408
rect 96429 491403 96495 491406
rect 102041 491403 102107 491406
rect 96429 491330 96495 491333
rect 99230 491330 99236 491332
rect 96429 491328 99236 491330
rect 96429 491272 96434 491328
rect 96490 491272 99236 491328
rect 96429 491270 99236 491272
rect 96429 491267 96495 491270
rect 99230 491268 99236 491270
rect 99300 491268 99306 491332
rect 115105 491196 115171 491197
rect 115054 491194 115060 491196
rect 115014 491134 115060 491194
rect 115124 491192 115171 491196
rect 115166 491136 115171 491192
rect 115054 491132 115060 491134
rect 115124 491132 115171 491136
rect 115105 491131 115171 491132
rect 65977 490514 66043 490517
rect 580349 490514 580415 490517
rect 65977 490512 580415 490514
rect 65977 490456 65982 490512
rect 66038 490456 580354 490512
rect 580410 490456 580415 490512
rect 65977 490454 580415 490456
rect 65977 490451 66043 490454
rect 580349 490451 580415 490454
rect 69982 489910 70226 489970
rect 67633 489834 67699 489837
rect 69982 489834 70042 489910
rect 67633 489832 70042 489834
rect 67633 489776 67638 489832
rect 67694 489776 70042 489832
rect 70166 489804 70226 489910
rect 67633 489774 70042 489776
rect 67633 489771 67699 489774
rect 99281 489426 99347 489429
rect 109033 489426 109099 489429
rect 99281 489424 109099 489426
rect 99281 489368 99286 489424
rect 99342 489368 109038 489424
rect 109094 489368 109099 489424
rect 99281 489366 109099 489368
rect 99281 489363 99347 489366
rect 109033 489363 109099 489366
rect 103421 489290 103487 489293
rect 99790 489288 103487 489290
rect 99790 489232 103426 489288
rect 103482 489232 103487 489288
rect 99790 489230 103487 489232
rect 99790 489124 99850 489230
rect 103421 489227 103487 489230
rect 117405 489154 117471 489157
rect 117998 489154 118004 489156
rect 117405 489152 118004 489154
rect 117405 489096 117410 489152
rect 117466 489096 118004 489152
rect 117405 489094 118004 489096
rect 117405 489091 117471 489094
rect 117998 489092 118004 489094
rect 118068 489092 118074 489156
rect -960 488596 480 488836
rect 118785 488612 118851 488613
rect 118734 488610 118740 488612
rect 118694 488550 118740 488610
rect 118804 488608 118851 488612
rect 118846 488552 118851 488608
rect 118734 488548 118740 488550
rect 118804 488548 118851 488552
rect 118785 488547 118851 488548
rect 103421 488474 103487 488477
rect 99974 488472 103487 488474
rect 99974 488440 103426 488472
rect 99790 488416 103426 488440
rect 103482 488416 103487 488472
rect 99790 488414 103487 488416
rect 99790 488380 100034 488414
rect 103421 488411 103487 488414
rect 99790 488308 99850 488380
rect 70166 487930 70226 488308
rect 99414 488004 99420 488068
rect 99484 488066 99490 488068
rect 112437 488066 112503 488069
rect 99484 488064 112503 488066
rect 99484 488008 112442 488064
rect 112498 488008 112503 488064
rect 99484 488006 112503 488008
rect 99484 488004 99490 488006
rect 112437 488003 112503 488006
rect 103421 487930 103487 487933
rect 64830 487870 70226 487930
rect 99790 487928 103487 487930
rect 99790 487872 103426 487928
rect 103482 487872 103487 487928
rect 99790 487870 103487 487872
rect 53598 487324 53604 487388
rect 53668 487386 53674 487388
rect 57646 487386 57652 487388
rect 53668 487326 57652 487386
rect 53668 487324 53674 487326
rect 57646 487324 57652 487326
rect 57716 487386 57722 487388
rect 64830 487386 64890 487870
rect 99790 487764 99850 487870
rect 103421 487867 103487 487870
rect 57716 487326 64890 487386
rect 57716 487324 57722 487326
rect 67633 487250 67699 487253
rect 70166 487250 70226 487628
rect 67633 487248 70226 487250
rect 67633 487192 67638 487248
rect 67694 487192 70226 487248
rect 67633 487190 70226 487192
rect 67633 487187 67699 487190
rect 67633 486570 67699 486573
rect 70166 486570 70226 486948
rect 99606 486706 99666 486948
rect 103421 486706 103487 486709
rect 99606 486704 103487 486706
rect 99606 486648 103426 486704
rect 103482 486648 103487 486704
rect 99606 486646 103487 486648
rect 103421 486643 103487 486646
rect 103421 486570 103487 486573
rect 67633 486568 70226 486570
rect 67633 486512 67638 486568
rect 67694 486512 70226 486568
rect 67633 486510 70226 486512
rect 99790 486568 103487 486570
rect 99790 486512 103426 486568
rect 103482 486512 103487 486568
rect 99790 486510 103487 486512
rect 67633 486507 67699 486510
rect 99790 486404 99850 486510
rect 103421 486507 103487 486510
rect 67633 485890 67699 485893
rect 70166 485890 70226 486268
rect 67633 485888 70226 485890
rect 67633 485832 67638 485888
rect 67694 485832 70226 485888
rect 67633 485830 70226 485832
rect 67633 485827 67699 485830
rect 111793 485756 111859 485757
rect 111742 485754 111748 485756
rect 111702 485694 111748 485754
rect 111812 485752 111859 485756
rect 111854 485696 111859 485752
rect 111742 485692 111748 485694
rect 111812 485692 111859 485696
rect 111793 485691 111859 485692
rect 122741 485754 122807 485757
rect 123334 485754 123340 485756
rect 122741 485752 123340 485754
rect 122741 485696 122746 485752
rect 122802 485696 123340 485752
rect 122741 485694 123340 485696
rect 122741 485691 122807 485694
rect 123334 485692 123340 485694
rect 123404 485692 123410 485756
rect 67633 485210 67699 485213
rect 70166 485210 70226 485588
rect 67633 485208 70226 485210
rect 67633 485152 67638 485208
rect 67694 485152 70226 485208
rect 67633 485150 70226 485152
rect 99790 485210 99850 485588
rect 102133 485210 102199 485213
rect 99790 485208 102199 485210
rect 99790 485152 102138 485208
rect 102194 485152 102199 485208
rect 99790 485150 102199 485152
rect 67633 485147 67699 485150
rect 102133 485147 102199 485150
rect 68645 484666 68711 484669
rect 70166 484666 70226 484908
rect 99606 484669 99666 484908
rect 70342 484666 70348 484668
rect 68645 484664 70348 484666
rect 68645 484608 68650 484664
rect 68706 484608 70348 484664
rect 68645 484606 70348 484608
rect 68645 484603 68711 484606
rect 70342 484604 70348 484606
rect 70412 484604 70418 484668
rect 99606 484664 99715 484669
rect 99606 484608 99654 484664
rect 99710 484608 99715 484664
rect 99606 484606 99715 484608
rect 99649 484603 99715 484606
rect 580349 484666 580415 484669
rect 583520 484666 584960 484756
rect 580349 484664 584960 484666
rect 580349 484608 580354 484664
rect 580410 484608 584960 484664
rect 580349 484606 584960 484608
rect 580349 484603 580415 484606
rect 583520 484516 584960 484606
rect 99966 484332 99972 484396
rect 100036 484394 100042 484396
rect 102317 484394 102383 484397
rect 100036 484392 102383 484394
rect 100036 484336 102322 484392
rect 102378 484336 102383 484392
rect 100036 484334 102383 484336
rect 100036 484332 100042 484334
rect 102317 484331 102383 484334
rect 67633 483986 67699 483989
rect 70166 483986 70226 484228
rect 67633 483984 70226 483986
rect 67633 483928 67638 483984
rect 67694 483928 70226 483984
rect 67633 483926 70226 483928
rect 67633 483923 67699 483926
rect 102133 483850 102199 483853
rect 99790 483848 102199 483850
rect 99790 483792 102138 483848
rect 102194 483792 102199 483848
rect 99790 483790 102199 483792
rect 99790 483684 99850 483790
rect 102133 483787 102199 483790
rect 122925 483306 122991 483309
rect 123334 483306 123340 483308
rect 122925 483304 123340 483306
rect 122925 483248 122930 483304
rect 122986 483248 123340 483304
rect 122925 483246 123340 483248
rect 122925 483243 122991 483246
rect 123334 483244 123340 483246
rect 123404 483244 123410 483308
rect 69982 483110 70226 483170
rect 69105 482898 69171 482901
rect 69982 482898 70042 483110
rect 70166 483004 70226 483110
rect 69105 482896 70042 482898
rect 69105 482840 69110 482896
rect 69166 482840 70042 482896
rect 69105 482838 70042 482840
rect 69105 482835 69171 482838
rect 67633 482626 67699 482629
rect 99606 482626 99666 482868
rect 102133 482626 102199 482629
rect 67633 482624 70226 482626
rect 67633 482568 67638 482624
rect 67694 482568 70226 482624
rect 67633 482566 70226 482568
rect 99606 482624 102199 482626
rect 99606 482568 102138 482624
rect 102194 482568 102199 482624
rect 99606 482566 102199 482568
rect 67633 482563 67699 482566
rect 70166 482324 70226 482566
rect 102133 482563 102199 482566
rect 99790 481810 99850 482188
rect 102133 481810 102199 481813
rect 99790 481808 102199 481810
rect 99790 481752 102138 481808
rect 102194 481752 102199 481808
rect 99790 481750 102199 481752
rect 102133 481747 102199 481750
rect 58065 481538 58131 481541
rect 59169 481538 59235 481541
rect 117037 481540 117103 481541
rect 117037 481538 117084 481540
rect 58065 481536 59235 481538
rect 58065 481480 58070 481536
rect 58126 481480 59174 481536
rect 59230 481480 59235 481536
rect 116956 481536 117084 481538
rect 117148 481538 117154 481540
rect 121678 481538 121684 481540
rect 58065 481478 59235 481480
rect 58065 481475 58131 481478
rect 59169 481475 59235 481478
rect 67633 481266 67699 481269
rect 70350 481266 70410 481508
rect 67633 481264 70410 481266
rect 67633 481208 67638 481264
rect 67694 481208 70410 481264
rect 67633 481206 70410 481208
rect 99790 481266 99850 481508
rect 116956 481480 117042 481536
rect 116956 481478 117084 481480
rect 117037 481476 117084 481478
rect 117148 481478 121684 481538
rect 117148 481476 117154 481478
rect 121678 481476 121684 481478
rect 121748 481476 121754 481540
rect 117037 481475 117103 481476
rect 102133 481266 102199 481269
rect 99790 481264 102199 481266
rect 99790 481208 102138 481264
rect 102194 481208 102199 481264
rect 99790 481206 102199 481208
rect 67633 481203 67699 481206
rect 102133 481203 102199 481206
rect 68001 481130 68067 481133
rect 69054 481130 69060 481132
rect 68001 481128 69060 481130
rect 68001 481072 68006 481128
rect 68062 481072 69060 481128
rect 68001 481070 69060 481072
rect 68001 481067 68067 481070
rect 69054 481068 69060 481070
rect 69124 481130 69130 481132
rect 102317 481130 102383 481133
rect 69124 481070 70226 481130
rect 69124 481068 69130 481070
rect 70166 480964 70226 481070
rect 99790 481128 102383 481130
rect 99790 481072 102322 481128
rect 102378 481072 102383 481128
rect 99790 481070 102383 481072
rect 99790 480964 99850 481070
rect 102317 481067 102383 481070
rect 54937 480314 55003 480317
rect 59169 480314 59235 480317
rect 54937 480312 59235 480314
rect 54937 480256 54942 480312
rect 54998 480256 59174 480312
rect 59230 480256 59235 480312
rect 54937 480254 59235 480256
rect 54937 480251 55003 480254
rect 59169 480251 59235 480254
rect 69982 480210 70226 480270
rect 61694 480116 61700 480180
rect 61764 480178 61770 480180
rect 64505 480178 64571 480181
rect 67633 480178 67699 480181
rect 69982 480178 70042 480210
rect 61764 480176 64890 480178
rect 61764 480120 64510 480176
rect 64566 480120 64890 480176
rect 61764 480118 64890 480120
rect 61764 480116 61770 480118
rect 64505 480115 64571 480118
rect 64830 479906 64890 480118
rect 67633 480176 70042 480178
rect 67633 480120 67638 480176
rect 67694 480120 70042 480176
rect 70166 480148 70226 480210
rect 67633 480118 70042 480120
rect 67633 480115 67699 480118
rect 99606 479906 99666 480148
rect 102133 479906 102199 479909
rect 64830 479846 70226 479906
rect 99606 479904 102199 479906
rect 99606 479848 102138 479904
rect 102194 479848 102199 479904
rect 99606 479846 102199 479848
rect 70166 479604 70226 479846
rect 102133 479843 102199 479846
rect 102133 479770 102199 479773
rect 104985 479772 105051 479773
rect 104934 479770 104940 479772
rect 99790 479768 102199 479770
rect 99790 479712 102138 479768
rect 102194 479712 102199 479768
rect 99790 479710 102199 479712
rect 104894 479710 104940 479770
rect 105004 479768 105051 479772
rect 105046 479712 105051 479768
rect 99790 479604 99850 479710
rect 102133 479707 102199 479710
rect 104934 479708 104940 479710
rect 105004 479708 105051 479712
rect 104985 479707 105051 479708
rect 67541 478546 67607 478549
rect 70350 478546 70410 478788
rect 67541 478544 70410 478546
rect 67541 478488 67546 478544
rect 67602 478488 70410 478544
rect 67541 478486 70410 478488
rect 67541 478483 67607 478486
rect 99790 477866 99850 478108
rect 102133 477866 102199 477869
rect 99790 477864 102199 477866
rect 99790 477808 102138 477864
rect 102194 477808 102199 477864
rect 99790 477806 102199 477808
rect 102133 477803 102199 477806
rect 65742 477668 65748 477732
rect 65812 477730 65818 477732
rect 67541 477730 67607 477733
rect 65812 477728 67607 477730
rect 65812 477672 67546 477728
rect 67602 477672 67607 477728
rect 65812 477670 67607 477672
rect 65812 477668 65818 477670
rect 67541 477667 67607 477670
rect 64965 477594 65031 477597
rect 65926 477594 65932 477596
rect 64965 477592 65932 477594
rect 64965 477536 64970 477592
rect 65026 477536 65932 477592
rect 64965 477534 65932 477536
rect 64965 477531 65031 477534
rect 65926 477532 65932 477534
rect 65996 477532 66002 477596
rect 62982 477396 62988 477460
rect 63052 477458 63058 477460
rect 63217 477458 63283 477461
rect 63052 477456 63283 477458
rect 63052 477400 63222 477456
rect 63278 477400 63283 477456
rect 115841 477458 115907 477461
rect 117681 477458 117747 477461
rect 129774 477458 129780 477460
rect 115841 477456 129780 477458
rect 63052 477398 63283 477400
rect 63052 477396 63058 477398
rect 63217 477395 63283 477398
rect 68369 477050 68435 477053
rect 68553 477050 68619 477053
rect 70166 477050 70226 477428
rect 99790 477186 99850 477428
rect 115841 477400 115846 477456
rect 115902 477400 117686 477456
rect 117742 477400 129780 477456
rect 115841 477398 129780 477400
rect 115841 477395 115907 477398
rect 117681 477395 117747 477398
rect 129774 477396 129780 477398
rect 129844 477396 129850 477460
rect 102409 477186 102475 477189
rect 99790 477184 102475 477186
rect 99790 477128 102414 477184
rect 102470 477128 102475 477184
rect 99790 477126 102475 477128
rect 102409 477123 102475 477126
rect 102133 477050 102199 477053
rect 68369 477048 70226 477050
rect 68369 476992 68374 477048
rect 68430 476992 68558 477048
rect 68614 476992 70226 477048
rect 68369 476990 70226 476992
rect 99790 477048 102199 477050
rect 99790 476992 102138 477048
rect 102194 476992 102199 477048
rect 99790 476990 102199 476992
rect 68369 476987 68435 476990
rect 68553 476987 68619 476990
rect 99790 476884 99850 476990
rect 102133 476987 102199 476990
rect 67633 476370 67699 476373
rect 70534 476370 70594 476748
rect 102317 476506 102383 476509
rect 67633 476368 70594 476370
rect 67633 476312 67638 476368
rect 67694 476312 70594 476368
rect 67633 476310 70594 476312
rect 99790 476504 102383 476506
rect 99790 476448 102322 476504
rect 102378 476448 102383 476504
rect 99790 476446 102383 476448
rect 67633 476307 67699 476310
rect 67725 476234 67791 476237
rect 67725 476232 70042 476234
rect 67725 476176 67730 476232
rect 67786 476176 70042 476232
rect 99790 476204 99850 476446
rect 102317 476443 102383 476446
rect 67725 476174 70042 476176
rect 67725 476171 67791 476174
rect 69982 476130 70042 476174
rect 106774 476172 106780 476236
rect 106844 476234 106850 476236
rect 108982 476234 108988 476236
rect 106844 476174 108988 476234
rect 106844 476172 106850 476174
rect 108982 476172 108988 476174
rect 109052 476172 109058 476236
rect 69982 476070 70226 476130
rect 70166 476068 70226 476070
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 67633 475690 67699 475693
rect 102133 475690 102199 475693
rect 67633 475688 70226 475690
rect 67633 475632 67638 475688
rect 67694 475632 70226 475688
rect 67633 475630 70226 475632
rect 67633 475627 67699 475630
rect 70166 475524 70226 475630
rect 99790 475688 102199 475690
rect 99790 475632 102138 475688
rect 102194 475632 102199 475688
rect 99790 475630 102199 475632
rect 99790 475524 99850 475630
rect 102133 475627 102199 475630
rect 102317 475146 102383 475149
rect 99790 475144 102383 475146
rect 99790 475088 102322 475144
rect 102378 475088 102383 475144
rect 99790 475086 102383 475088
rect 67633 475010 67699 475013
rect 67633 475008 70226 475010
rect 67633 474952 67638 475008
rect 67694 474952 70226 475008
rect 67633 474950 70226 474952
rect 67633 474947 67699 474950
rect 70166 474844 70226 474950
rect 99790 474844 99850 475086
rect 102317 475083 102383 475086
rect 49601 474738 49667 474741
rect 55949 474738 56015 474741
rect 49601 474736 56015 474738
rect 49601 474680 49606 474736
rect 49662 474680 55954 474736
rect 56010 474680 56015 474736
rect 49601 474678 56015 474680
rect 49601 474675 49667 474678
rect 55949 474675 56015 474678
rect 67449 474330 67515 474333
rect 102133 474330 102199 474333
rect 67449 474328 70226 474330
rect 67449 474272 67454 474328
rect 67510 474272 70226 474328
rect 67449 474270 70226 474272
rect 67449 474267 67515 474270
rect 70166 474164 70226 474270
rect 99790 474328 102199 474330
rect 99790 474272 102138 474328
rect 102194 474272 102199 474328
rect 99790 474270 102199 474272
rect 99790 474164 99850 474270
rect 102133 474267 102199 474270
rect 55070 473996 55076 474060
rect 55140 474058 55146 474060
rect 66478 474058 66484 474060
rect 55140 473998 66484 474058
rect 55140 473996 55146 473998
rect 66478 473996 66484 473998
rect 66548 473996 66554 474060
rect 66478 473724 66484 473788
rect 66548 473786 66554 473788
rect 66548 473726 70226 473786
rect 66548 473724 66554 473726
rect 70166 473484 70226 473726
rect 66662 473316 66668 473380
rect 66732 473378 66738 473380
rect 67449 473378 67515 473381
rect 66732 473376 67515 473378
rect 66732 473320 67454 473376
rect 67510 473320 67515 473376
rect 66732 473318 67515 473320
rect 66732 473316 66738 473318
rect 67449 473315 67515 473318
rect 102133 472970 102199 472973
rect 99790 472968 102199 472970
rect 99790 472912 102138 472968
rect 102194 472912 102199 472968
rect 99790 472910 102199 472912
rect 99790 472804 99850 472910
rect 102133 472907 102199 472910
rect 67633 472698 67699 472701
rect 67633 472696 70226 472698
rect 67633 472640 67638 472696
rect 67694 472640 70226 472696
rect 67633 472638 70226 472640
rect 67633 472635 67699 472638
rect 70166 472124 70226 472638
rect 102317 472426 102383 472429
rect 99790 472424 102383 472426
rect 99790 472368 102322 472424
rect 102378 472368 102383 472424
rect 99790 472366 102383 472368
rect 99790 472124 99850 472366
rect 102317 472363 102383 472366
rect 67633 471610 67699 471613
rect 102133 471610 102199 471613
rect 67633 471608 70226 471610
rect 67633 471552 67638 471608
rect 67694 471552 70226 471608
rect 67633 471550 70226 471552
rect 67633 471547 67699 471550
rect 70166 471444 70226 471550
rect 99790 471608 102199 471610
rect 99790 471552 102138 471608
rect 102194 471552 102199 471608
rect 99790 471550 102199 471552
rect 99790 471444 99850 471550
rect 102133 471547 102199 471550
rect 579889 471474 579955 471477
rect 583520 471474 584960 471564
rect 579889 471472 584960 471474
rect 579889 471416 579894 471472
rect 579950 471416 584960 471472
rect 579889 471414 584960 471416
rect 579889 471411 579955 471414
rect 583520 471324 584960 471414
rect 67633 471066 67699 471069
rect 67633 471064 70226 471066
rect 67633 471008 67638 471064
rect 67694 471008 70226 471064
rect 67633 471006 70226 471008
rect 67633 471003 67699 471006
rect 70166 470764 70226 471006
rect 102317 470930 102383 470933
rect 99790 470928 102383 470930
rect 99790 470872 102322 470928
rect 102378 470872 102383 470928
rect 99790 470870 102383 470872
rect 99790 470764 99850 470870
rect 102317 470867 102383 470870
rect 107561 470658 107627 470661
rect 107694 470658 107700 470660
rect 107561 470656 107700 470658
rect 107561 470600 107566 470656
rect 107622 470600 107700 470656
rect 107561 470598 107700 470600
rect 107561 470595 107627 470598
rect 107694 470596 107700 470598
rect 107764 470596 107770 470660
rect 66069 470524 66135 470525
rect 66069 470520 66116 470524
rect 66180 470522 66186 470524
rect 66069 470464 66074 470520
rect 66069 470460 66116 470464
rect 66180 470462 66226 470522
rect 66180 470460 66186 470462
rect 66069 470459 66135 470460
rect 102133 470250 102199 470253
rect 99790 470248 102199 470250
rect 99790 470192 102138 470248
rect 102194 470192 102199 470248
rect 99790 470190 102199 470192
rect 99790 470084 99850 470190
rect 102133 470187 102199 470190
rect 67633 469706 67699 469709
rect 70350 469706 70410 469948
rect 102869 469706 102935 469709
rect 67633 469704 70410 469706
rect 67633 469648 67638 469704
rect 67694 469648 70410 469704
rect 67633 469646 70410 469648
rect 99790 469704 102935 469706
rect 99790 469648 102874 469704
rect 102930 469648 102935 469704
rect 99790 469646 102935 469648
rect 67633 469643 67699 469646
rect 67725 469570 67791 469573
rect 67725 469568 70226 469570
rect 67725 469512 67730 469568
rect 67786 469512 70226 469568
rect 67725 469510 70226 469512
rect 67725 469507 67791 469510
rect 70166 469404 70226 469510
rect 99790 469404 99850 469646
rect 102869 469643 102935 469646
rect 103605 469026 103671 469029
rect 99790 469024 103671 469026
rect 99790 468968 103610 469024
rect 103666 468968 103671 469024
rect 99790 468966 103671 468968
rect 99790 468724 99850 468966
rect 103605 468963 103671 468966
rect 67725 468346 67791 468349
rect 70166 468346 70226 468588
rect 67725 468344 70226 468346
rect 67725 468288 67730 468344
rect 67786 468288 70226 468344
rect 67725 468286 70226 468288
rect 67725 468283 67791 468286
rect 67633 468210 67699 468213
rect 67633 468208 70226 468210
rect 67633 468152 67638 468208
rect 67694 468152 70226 468208
rect 67633 468150 70226 468152
rect 67633 468147 67699 468150
rect 70166 468044 70226 468150
rect 99790 466986 99850 467228
rect 103145 466986 103211 466989
rect 99790 466984 103211 466986
rect 99790 466928 103150 466984
rect 103206 466928 103211 466984
rect 99790 466926 103211 466928
rect 103145 466923 103211 466926
rect 67633 466850 67699 466853
rect 102133 466850 102199 466853
rect 67633 466848 70226 466850
rect 67633 466792 67638 466848
rect 67694 466792 70226 466848
rect 67633 466790 70226 466792
rect 67633 466787 67699 466790
rect 70166 466684 70226 466790
rect 99790 466848 102199 466850
rect 99790 466792 102138 466848
rect 102194 466792 102199 466848
rect 99790 466790 102199 466792
rect 99790 466684 99850 466790
rect 102133 466787 102199 466790
rect 67725 466170 67791 466173
rect 102133 466170 102199 466173
rect 67725 466168 70226 466170
rect 67725 466112 67730 466168
rect 67786 466112 70226 466168
rect 67725 466110 70226 466112
rect 67725 466107 67791 466110
rect 70166 466004 70226 466110
rect 99790 466168 102199 466170
rect 99790 466112 102138 466168
rect 102194 466112 102199 466168
rect 99790 466110 102199 466112
rect 99790 466004 99850 466110
rect 102133 466107 102199 466110
rect 67633 465626 67699 465629
rect 102133 465626 102199 465629
rect 67633 465624 70410 465626
rect 67633 465568 67638 465624
rect 67694 465568 70410 465624
rect 67633 465566 70410 465568
rect 67633 465563 67699 465566
rect 70350 465324 70410 465566
rect 99790 465624 102199 465626
rect 99790 465568 102138 465624
rect 102194 465568 102199 465624
rect 99790 465566 102199 465568
rect 99790 465324 99850 465566
rect 102133 465563 102199 465566
rect 102133 464810 102199 464813
rect 99790 464808 102199 464810
rect 99790 464752 102138 464808
rect 102194 464752 102199 464808
rect 99790 464750 102199 464752
rect 99790 464644 99850 464750
rect 102133 464747 102199 464750
rect 67817 464130 67883 464133
rect 70166 464130 70226 464508
rect 102133 464130 102199 464133
rect 67817 464128 70226 464130
rect 67817 464072 67822 464128
rect 67878 464072 70226 464128
rect 67817 464070 70226 464072
rect 99790 464128 102199 464130
rect 99790 464072 102138 464128
rect 102194 464072 102199 464128
rect 99790 464070 102199 464072
rect 67817 464067 67883 464070
rect 99790 463964 99850 464070
rect 102133 464067 102199 464070
rect 67633 463722 67699 463725
rect 67633 463720 69858 463722
rect 67633 463664 67638 463720
rect 67694 463664 69858 463720
rect 67633 463662 69858 463664
rect 67633 463659 67699 463662
rect 69798 463586 69858 463662
rect 70350 463586 70410 463828
rect 69798 463526 70410 463586
rect 67633 463450 67699 463453
rect 102133 463450 102199 463453
rect 67633 463448 70226 463450
rect 67633 463392 67638 463448
rect 67694 463392 70226 463448
rect 67633 463390 70226 463392
rect 67633 463387 67699 463390
rect 70166 463284 70226 463390
rect 99790 463448 102199 463450
rect 99790 463392 102138 463448
rect 102194 463392 102199 463448
rect 99790 463390 102199 463392
rect 99790 463284 99850 463390
rect 102133 463387 102199 463390
rect 67725 462906 67791 462909
rect 67725 462904 70410 462906
rect 67725 462848 67730 462904
rect 67786 462848 70410 462904
rect 67725 462846 70410 462848
rect 67725 462843 67791 462846
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect 70350 462604 70410 462846
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 102133 462090 102199 462093
rect 99790 462088 102199 462090
rect 99790 462032 102138 462088
rect 102194 462032 102199 462088
rect 99790 462030 102199 462032
rect 99790 461924 99850 462030
rect 102133 462027 102199 462030
rect 102225 461546 102291 461549
rect 99790 461544 102291 461546
rect 99790 461488 102230 461544
rect 102286 461488 102291 461544
rect 99790 461486 102291 461488
rect 67633 461410 67699 461413
rect 67633 461408 70226 461410
rect 67633 461352 67638 461408
rect 67694 461352 70226 461408
rect 67633 461350 70226 461352
rect 67633 461347 67699 461350
rect 70166 461244 70226 461350
rect 99790 461244 99850 461486
rect 102225 461483 102291 461486
rect 67633 460730 67699 460733
rect 102225 460730 102291 460733
rect 67633 460728 70226 460730
rect 67633 460672 67638 460728
rect 67694 460672 70226 460728
rect 67633 460670 70226 460672
rect 67633 460667 67699 460670
rect 70166 460564 70226 460670
rect 99790 460728 102291 460730
rect 99790 460672 102230 460728
rect 102286 460672 102291 460728
rect 99790 460670 102291 460672
rect 99790 460564 99850 460670
rect 102225 460667 102291 460670
rect 67725 460186 67791 460189
rect 102133 460186 102199 460189
rect 67725 460184 70226 460186
rect 67725 460128 67730 460184
rect 67786 460128 70226 460184
rect 67725 460126 70226 460128
rect 67725 460123 67791 460126
rect 70166 459884 70226 460126
rect 99606 460184 102199 460186
rect 99606 460128 102138 460184
rect 102194 460128 102199 460184
rect 99606 460126 102199 460128
rect 99606 459884 99666 460126
rect 102133 460123 102199 460126
rect 102133 459370 102199 459373
rect 99790 459368 102199 459370
rect 99790 459312 102138 459368
rect 102194 459312 102199 459368
rect 99790 459310 102199 459312
rect 99790 459204 99850 459310
rect 102133 459307 102199 459310
rect 67633 458826 67699 458829
rect 70350 458826 70410 459068
rect 67633 458824 70410 458826
rect 67633 458768 67638 458824
rect 67694 458768 70410 458824
rect 67633 458766 70410 458768
rect 67633 458763 67699 458766
rect 67633 458690 67699 458693
rect 103237 458690 103303 458693
rect 67633 458688 70226 458690
rect 67633 458632 67638 458688
rect 67694 458632 70226 458688
rect 67633 458630 70226 458632
rect 67633 458627 67699 458630
rect 70166 458524 70226 458630
rect 99790 458688 103303 458690
rect 99790 458632 103242 458688
rect 103298 458632 103303 458688
rect 99790 458630 103303 458632
rect 99790 458524 99850 458630
rect 103237 458627 103303 458630
rect 579613 458146 579679 458149
rect 583520 458146 584960 458236
rect 579613 458144 584960 458146
rect 579613 458088 579618 458144
rect 579674 458088 584960 458144
rect 579613 458086 584960 458088
rect 579613 458083 579679 458086
rect 67633 458010 67699 458013
rect 102133 458010 102199 458013
rect 67633 458008 70226 458010
rect 67633 457952 67638 458008
rect 67694 457952 70226 458008
rect 67633 457950 70226 457952
rect 67633 457947 67699 457950
rect 70166 457844 70226 457950
rect 99790 458008 102199 458010
rect 99790 457952 102138 458008
rect 102194 457952 102199 458008
rect 583520 457996 584960 458086
rect 99790 457950 102199 457952
rect 99790 457844 99850 457950
rect 102133 457947 102199 457950
rect 67725 457466 67791 457469
rect 67725 457464 70226 457466
rect 67725 457408 67730 457464
rect 67786 457408 70226 457464
rect 67725 457406 70226 457408
rect 67725 457403 67791 457406
rect 70166 457164 70226 457406
rect 102133 456650 102199 456653
rect 99790 456648 102199 456650
rect 99790 456592 102138 456648
rect 102194 456592 102199 456648
rect 99790 456590 102199 456592
rect 99790 456484 99850 456590
rect 102133 456587 102199 456590
rect 102225 456106 102291 456109
rect 99790 456104 102291 456106
rect 99790 456048 102230 456104
rect 102286 456048 102291 456104
rect 99790 456046 102291 456048
rect 67633 455970 67699 455973
rect 67633 455968 70226 455970
rect 67633 455912 67638 455968
rect 67694 455912 70226 455968
rect 67633 455910 70226 455912
rect 67633 455907 67699 455910
rect 70166 455804 70226 455910
rect 99790 455804 99850 456046
rect 102225 456043 102291 456046
rect 67633 455290 67699 455293
rect 102133 455290 102199 455293
rect 67633 455288 70226 455290
rect 67633 455232 67638 455288
rect 67694 455232 70226 455288
rect 67633 455230 70226 455232
rect 67633 455227 67699 455230
rect 70166 455124 70226 455230
rect 99790 455288 102199 455290
rect 99790 455232 102138 455288
rect 102194 455232 102199 455288
rect 99790 455230 102199 455232
rect 99790 455124 99850 455230
rect 102133 455227 102199 455230
rect 68134 454684 68140 454748
rect 68204 454746 68210 454748
rect 68870 454746 68876 454748
rect 68204 454686 68876 454746
rect 68204 454684 68210 454686
rect 68870 454684 68876 454686
rect 68940 454746 68946 454748
rect 68940 454686 70226 454746
rect 68940 454684 68946 454686
rect 70166 454444 70226 454686
rect 102133 454610 102199 454613
rect 99790 454608 102199 454610
rect 99790 454552 102138 454608
rect 102194 454552 102199 454608
rect 99790 454550 102199 454552
rect 99790 454444 99850 454550
rect 102133 454547 102199 454550
rect 67633 453930 67699 453933
rect 67633 453928 70226 453930
rect 67633 453872 67638 453928
rect 67694 453872 70226 453928
rect 67633 453870 70226 453872
rect 67633 453867 67699 453870
rect 70166 453764 70226 453870
rect 99790 453386 99850 453628
rect 102869 453386 102935 453389
rect 99790 453384 102935 453386
rect 99790 453328 102874 453384
rect 102930 453328 102935 453384
rect 99790 453326 102935 453328
rect 102869 453323 102935 453326
rect 125593 453386 125659 453389
rect 125726 453386 125732 453388
rect 125593 453384 125732 453386
rect 125593 453328 125598 453384
rect 125654 453328 125732 453384
rect 125593 453326 125732 453328
rect 125593 453323 125659 453326
rect 125726 453324 125732 453326
rect 125796 453324 125802 453388
rect 67633 453250 67699 453253
rect 102133 453250 102199 453253
rect 67633 453248 70226 453250
rect 67633 453192 67638 453248
rect 67694 453192 70226 453248
rect 67633 453190 70226 453192
rect 67633 453187 67699 453190
rect 70166 453084 70226 453190
rect 99790 453248 102199 453250
rect 99790 453192 102138 453248
rect 102194 453192 102199 453248
rect 99790 453190 102199 453192
rect 99790 453084 99850 453190
rect 102133 453187 102199 453190
rect 102133 452570 102199 452573
rect 99790 452568 102199 452570
rect 99790 452512 102138 452568
rect 102194 452512 102199 452568
rect 99790 452510 102199 452512
rect 99790 452404 99850 452510
rect 102133 452507 102199 452510
rect 69197 451890 69263 451893
rect 70166 451890 70226 452268
rect 69197 451888 70226 451890
rect 69197 451832 69202 451888
rect 69258 451832 70226 451888
rect 69197 451830 70226 451832
rect 69197 451827 69263 451830
rect 68737 451346 68803 451349
rect 70350 451346 70410 451588
rect 68737 451344 70410 451346
rect 68737 451288 68742 451344
rect 68798 451288 70410 451344
rect 68737 451286 70410 451288
rect 68737 451283 68803 451286
rect 101489 451210 101555 451213
rect 99790 451208 101555 451210
rect 99790 451152 101494 451208
rect 101550 451152 101555 451208
rect 99790 451150 101555 451152
rect 99790 451044 99850 451150
rect 101489 451147 101555 451150
rect 103605 450666 103671 450669
rect 99790 450664 103671 450666
rect 99790 450608 103610 450664
rect 103666 450608 103671 450664
rect 99790 450606 103671 450608
rect 99790 450364 99850 450606
rect 103605 450603 103671 450606
rect 67633 449986 67699 449989
rect 70166 449986 70226 450228
rect 67633 449984 70226 449986
rect 67633 449928 67638 449984
rect 67694 449928 70226 449984
rect 67633 449926 70226 449928
rect 67633 449923 67699 449926
rect 103697 449850 103763 449853
rect 104249 449850 104315 449853
rect 99790 449848 104315 449850
rect 99790 449792 103702 449848
rect 103758 449792 104254 449848
rect 104310 449792 104315 449848
rect 99790 449790 104315 449792
rect 99790 449684 99850 449790
rect 103697 449787 103763 449790
rect 104249 449787 104315 449790
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 67725 449306 67791 449309
rect 70166 449306 70226 449548
rect 107469 449444 107535 449445
rect 107469 449440 107516 449444
rect 107580 449442 107586 449444
rect 107469 449384 107474 449440
rect 107469 449380 107516 449384
rect 107580 449382 107626 449442
rect 107580 449380 107586 449382
rect 107469 449379 107535 449380
rect 102133 449306 102199 449309
rect 67725 449304 70226 449306
rect 67725 449248 67730 449304
rect 67786 449248 70226 449304
rect 67725 449246 70226 449248
rect 99790 449304 102199 449306
rect 99790 449248 102138 449304
rect 102194 449248 102199 449304
rect 99790 449246 102199 449248
rect 67725 449243 67791 449246
rect 67633 449170 67699 449173
rect 67633 449168 70226 449170
rect 67633 449112 67638 449168
rect 67694 449112 70226 449168
rect 67633 449110 70226 449112
rect 67633 449107 67699 449110
rect 70166 449004 70226 449110
rect 99790 449004 99850 449246
rect 102133 449243 102199 449246
rect 61878 448564 61884 448628
rect 61948 448626 61954 448628
rect 63309 448626 63375 448629
rect 67725 448626 67791 448629
rect 61948 448624 67791 448626
rect 61948 448568 63314 448624
rect 63370 448568 67730 448624
rect 67786 448568 67791 448624
rect 61948 448566 67791 448568
rect 61948 448564 61954 448566
rect 63309 448563 63375 448566
rect 67725 448563 67791 448566
rect 107469 448626 107535 448629
rect 144913 448626 144979 448629
rect 107469 448624 144979 448626
rect 107469 448568 107474 448624
rect 107530 448568 144918 448624
rect 144974 448568 144979 448624
rect 107469 448566 144979 448568
rect 107469 448563 107535 448566
rect 144913 448563 144979 448566
rect 102133 448490 102199 448493
rect 99790 448488 102199 448490
rect 99790 448432 102138 448488
rect 102194 448432 102199 448488
rect 99790 448430 102199 448432
rect 99790 448324 99850 448430
rect 102133 448427 102199 448430
rect 67725 447810 67791 447813
rect 70166 447810 70226 448188
rect 102225 447946 102291 447949
rect 67725 447808 70226 447810
rect 67725 447752 67730 447808
rect 67786 447752 70226 447808
rect 67725 447750 70226 447752
rect 99790 447944 102291 447946
rect 99790 447888 102230 447944
rect 102286 447888 102291 447944
rect 99790 447886 102291 447888
rect 67725 447747 67791 447750
rect 99790 447644 99850 447886
rect 102225 447883 102291 447886
rect 67633 447266 67699 447269
rect 70166 447266 70226 447508
rect 67633 447264 70226 447266
rect 67633 447208 67638 447264
rect 67694 447208 70226 447264
rect 67633 447206 70226 447208
rect 67633 447203 67699 447206
rect 101949 447130 102015 447133
rect 99790 447128 102015 447130
rect 99790 447072 101954 447128
rect 102010 447072 102015 447128
rect 99790 447070 102015 447072
rect 99790 446964 99850 447070
rect 101949 447067 102015 447070
rect 67725 446586 67791 446589
rect 70166 446586 70226 446828
rect 67725 446584 70226 446586
rect 67725 446528 67730 446584
rect 67786 446528 70226 446584
rect 67725 446526 70226 446528
rect 67725 446523 67791 446526
rect 67633 446450 67699 446453
rect 67633 446448 70226 446450
rect 67633 446392 67638 446448
rect 67694 446392 70226 446448
rect 67633 446390 70226 446392
rect 67633 446387 67699 446390
rect 70166 446284 70226 446390
rect 103830 445770 103836 445772
rect 99790 445710 103836 445770
rect 99790 445604 99850 445710
rect 103830 445708 103836 445710
rect 103900 445708 103906 445772
rect 68185 445498 68251 445501
rect 68553 445498 68619 445501
rect 68185 445496 70226 445498
rect 68185 445440 68190 445496
rect 68246 445440 68558 445496
rect 68614 445440 70226 445496
rect 68185 445438 70226 445440
rect 68185 445435 68251 445438
rect 68553 445435 68619 445438
rect 70166 444924 70226 445438
rect 103145 445090 103211 445093
rect 99790 445088 103211 445090
rect 99790 445032 103150 445088
rect 103206 445032 103211 445088
rect 99790 445030 103211 445032
rect 99790 444924 99850 445030
rect 103145 445027 103211 445030
rect 124949 444954 125015 444957
rect 128670 444954 128676 444956
rect 108990 444952 128676 444954
rect 108990 444896 124954 444952
rect 125010 444896 128676 444952
rect 108990 444894 128676 444896
rect 108990 444546 109050 444894
rect 124949 444891 125015 444894
rect 128670 444892 128676 444894
rect 128740 444892 128746 444956
rect 583520 444668 584960 444908
rect 103470 444486 109050 444546
rect 69982 444350 70226 444410
rect 68277 444274 68343 444277
rect 68921 444274 68987 444277
rect 69982 444274 70042 444350
rect 68277 444272 70042 444274
rect 68277 444216 68282 444272
rect 68338 444216 68926 444272
rect 68982 444216 70042 444272
rect 70166 444244 70226 444350
rect 99790 444390 100034 444410
rect 99790 444350 100218 444390
rect 99790 444244 99850 444350
rect 99974 444330 100218 444350
rect 100158 444274 100218 444330
rect 103470 444274 103530 444486
rect 103830 444348 103836 444412
rect 103900 444410 103906 444412
rect 104157 444410 104223 444413
rect 103900 444408 104223 444410
rect 103900 444352 104162 444408
rect 104218 444352 104223 444408
rect 103900 444350 104223 444352
rect 103900 444348 103906 444350
rect 104157 444347 104223 444350
rect 68277 444214 70042 444216
rect 100158 444214 103530 444274
rect 68277 444211 68343 444214
rect 68921 444211 68987 444214
rect 67633 443730 67699 443733
rect 99281 443730 99347 443733
rect 114502 443730 114508 443732
rect 67633 443728 70226 443730
rect 67633 443672 67638 443728
rect 67694 443672 70226 443728
rect 67633 443670 70226 443672
rect 67633 443667 67699 443670
rect 70166 443564 70226 443670
rect 99281 443728 114508 443730
rect 99281 443672 99286 443728
rect 99342 443672 114508 443728
rect 99281 443670 114508 443672
rect 99281 443667 99347 443670
rect 114502 443668 114508 443670
rect 114572 443668 114578 443732
rect 99465 443186 99531 443189
rect 99606 443186 99666 443428
rect 102593 443186 102659 443189
rect 99465 443184 102659 443186
rect 99465 443128 99470 443184
rect 99526 443128 102598 443184
rect 102654 443128 102659 443184
rect 99465 443126 102659 443128
rect 99465 443123 99531 443126
rect 102593 443123 102659 443126
rect 67633 442506 67699 442509
rect 70350 442506 70410 442748
rect 99606 442509 99666 442748
rect 99557 442506 99666 442509
rect 102685 442506 102751 442509
rect 67633 442504 70410 442506
rect 67633 442448 67638 442504
rect 67694 442448 70410 442504
rect 67633 442446 70410 442448
rect 99476 442504 102751 442506
rect 99476 442448 99562 442504
rect 99618 442448 102690 442504
rect 102746 442448 102751 442504
rect 99476 442446 102751 442448
rect 67633 442443 67699 442446
rect 99557 442443 99623 442446
rect 102685 442443 102751 442446
rect 67633 442370 67699 442373
rect 67633 442368 70226 442370
rect 67633 442312 67638 442368
rect 67694 442312 70226 442368
rect 67633 442310 70226 442312
rect 67633 442307 67699 442310
rect 70166 442204 70226 442310
rect 99414 442308 99420 442372
rect 99484 442370 99490 442372
rect 110638 442370 110644 442372
rect 99484 442310 110644 442370
rect 99484 442308 99490 442310
rect 110638 442308 110644 442310
rect 110708 442308 110714 442372
rect 99606 441826 99666 442068
rect 101254 441826 101260 441828
rect 99606 441766 101260 441826
rect 101254 441764 101260 441766
rect 101324 441826 101330 441828
rect 103145 441826 103211 441829
rect 101324 441824 103211 441826
rect 101324 441768 103150 441824
rect 103206 441768 103211 441824
rect 101324 441766 103211 441768
rect 101324 441764 101330 441766
rect 103145 441763 103211 441766
rect 67633 441146 67699 441149
rect 70350 441146 70410 441388
rect 67633 441144 70410 441146
rect 67633 441088 67638 441144
rect 67694 441088 70410 441144
rect 67633 441086 70410 441088
rect 67633 441083 67699 441086
rect 67633 441010 67699 441013
rect 67633 441008 70226 441010
rect 67633 440952 67638 441008
rect 67694 440952 70226 441008
rect 67633 440950 70226 440952
rect 67633 440947 67699 440950
rect 70166 440844 70226 440950
rect 99790 440874 99850 441388
rect 103145 440874 103211 440877
rect 99790 440872 103211 440874
rect 99790 440816 103150 440872
rect 103206 440816 103211 440872
rect 99790 440814 103211 440816
rect 103145 440811 103211 440814
rect 100753 440330 100819 440333
rect 102133 440330 102199 440333
rect 99790 440328 102199 440330
rect 99790 440272 100758 440328
rect 100814 440272 102138 440328
rect 102194 440272 102199 440328
rect 99790 440270 102199 440272
rect 99790 440164 99850 440270
rect 100753 440267 100819 440270
rect 102133 440267 102199 440270
rect 97717 439786 97783 439789
rect 99966 439786 99972 439788
rect 97717 439784 99972 439786
rect 97717 439728 97722 439784
rect 97778 439728 99972 439784
rect 97717 439726 99972 439728
rect 97717 439723 97783 439726
rect 99966 439724 99972 439726
rect 100036 439724 100042 439788
rect 60590 439452 60596 439516
rect 60660 439514 60666 439516
rect 70342 439514 70348 439516
rect 60660 439454 70348 439514
rect 60660 439452 60666 439454
rect 70342 439452 70348 439454
rect 70412 439514 70418 439516
rect 88977 439514 89043 439517
rect 111926 439514 111932 439516
rect 70412 439454 74550 439514
rect 70412 439452 70418 439454
rect 69054 438908 69060 438972
rect 69124 438970 69130 438972
rect 71037 438970 71103 438973
rect 69124 438968 71103 438970
rect 69124 438912 71042 438968
rect 71098 438912 71103 438968
rect 69124 438910 71103 438912
rect 74490 438970 74550 439454
rect 88977 439512 111932 439514
rect 88977 439456 88982 439512
rect 89038 439456 111932 439512
rect 88977 439454 111932 439456
rect 88977 439451 89043 439454
rect 111926 439452 111932 439454
rect 111996 439452 112002 439516
rect 84193 438970 84259 438973
rect 74490 438968 84259 438970
rect 74490 438912 84198 438968
rect 84254 438912 84259 438968
rect 74490 438910 84259 438912
rect 69124 438908 69130 438910
rect 71037 438907 71103 438910
rect 84193 438907 84259 438910
rect 96613 438970 96679 438973
rect 97717 438970 97783 438973
rect 96613 438968 97783 438970
rect 96613 438912 96618 438968
rect 96674 438912 97722 438968
rect 97778 438912 97783 438968
rect 96613 438910 97783 438912
rect 96613 438907 96679 438910
rect 97717 438907 97783 438910
rect 123753 438970 123819 438973
rect 124806 438970 124812 438972
rect 123753 438968 124812 438970
rect 123753 438912 123758 438968
rect 123814 438912 124812 438968
rect 123753 438910 124812 438912
rect 123753 438907 123819 438910
rect 124806 438908 124812 438910
rect 124876 438908 124882 438972
rect 57830 438092 57836 438156
rect 57900 438154 57906 438156
rect 75453 438154 75519 438157
rect 57900 438152 75519 438154
rect 57900 438096 75458 438152
rect 75514 438096 75519 438152
rect 57900 438094 75519 438096
rect 57900 438092 57906 438094
rect 75453 438091 75519 438094
rect 98361 437882 98427 437885
rect 99281 437882 99347 437885
rect 98361 437880 99347 437882
rect 98361 437824 98366 437880
rect 98422 437824 99286 437880
rect 99342 437824 99347 437880
rect 98361 437822 99347 437824
rect 98361 437819 98427 437822
rect 99281 437819 99347 437822
rect 69105 437610 69171 437613
rect 73797 437610 73863 437613
rect 69105 437608 73863 437610
rect 69105 437552 69110 437608
rect 69166 437552 73802 437608
rect 73858 437552 73863 437608
rect 69105 437550 73863 437552
rect 69105 437547 69171 437550
rect 73797 437547 73863 437550
rect 59118 437412 59124 437476
rect 59188 437474 59194 437476
rect 80973 437474 81039 437477
rect 59188 437472 81039 437474
rect 59188 437416 80978 437472
rect 81034 437416 81039 437472
rect 59188 437414 81039 437416
rect 59188 437412 59194 437414
rect 80973 437411 81039 437414
rect 93669 437474 93735 437477
rect 106774 437474 106780 437476
rect 93669 437472 106780 437474
rect 93669 437416 93674 437472
rect 93730 437416 106780 437472
rect 93669 437414 106780 437416
rect 93669 437411 93735 437414
rect 106774 437412 106780 437414
rect 106844 437412 106850 437476
rect -960 436508 480 436748
rect 80053 436522 80119 436525
rect 80973 436522 81039 436525
rect 80053 436520 81039 436522
rect 80053 436464 80058 436520
rect 80114 436464 80978 436520
rect 81034 436464 81039 436520
rect 80053 436462 81039 436464
rect 80053 436459 80119 436462
rect 80973 436459 81039 436462
rect 69013 434754 69079 434757
rect 78581 434754 78647 434757
rect 69013 434752 78647 434754
rect 69013 434696 69018 434752
rect 69074 434696 78586 434752
rect 78642 434696 78647 434752
rect 69013 434694 78647 434696
rect 69013 434691 69079 434694
rect 78581 434691 78647 434694
rect 69013 433804 69079 433805
rect 69013 433800 69060 433804
rect 69124 433802 69130 433804
rect 69013 433744 69018 433800
rect 69013 433740 69060 433744
rect 69124 433742 69170 433802
rect 69124 433740 69130 433742
rect 69013 433739 69079 433740
rect 42701 433258 42767 433261
rect 44030 433258 44036 433260
rect 42701 433256 44036 433258
rect 42701 433200 42706 433256
rect 42762 433200 44036 433256
rect 42701 433198 44036 433200
rect 42701 433195 42767 433198
rect 44030 433196 44036 433198
rect 44100 433258 44106 433260
rect 74533 433258 74599 433261
rect 44100 433256 74599 433258
rect 44100 433200 74538 433256
rect 74594 433200 74599 433256
rect 44100 433198 74599 433200
rect 44100 433196 44106 433198
rect 74533 433195 74599 433198
rect 579797 431626 579863 431629
rect 583520 431626 584960 431716
rect 579797 431624 584960 431626
rect 579797 431568 579802 431624
rect 579858 431568 584960 431624
rect 579797 431566 584960 431568
rect 579797 431563 579863 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 579981 418298 580047 418301
rect 583520 418298 584960 418388
rect 579981 418296 584960 418298
rect 579981 418240 579986 418296
rect 580042 418240 584960 418296
rect 579981 418238 584960 418240
rect 579981 418235 580047 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 579613 404970 579679 404973
rect 583520 404970 584960 405060
rect 579613 404968 584960 404970
rect 579613 404912 579618 404968
rect 579674 404912 584960 404968
rect 579613 404910 584960 404912
rect 579613 404907 579679 404910
rect 583520 404820 584960 404910
rect 115105 400212 115171 400213
rect 115054 400210 115060 400212
rect 115014 400150 115060 400210
rect 115124 400208 115171 400212
rect 115166 400152 115171 400208
rect 115054 400148 115060 400150
rect 115124 400148 115171 400152
rect 115105 400147 115171 400148
rect 48078 397972 48084 398036
rect 48148 398034 48154 398036
rect 90081 398034 90147 398037
rect 48148 398032 90147 398034
rect 48148 397976 90086 398032
rect 90142 397976 90147 398032
rect 48148 397974 90147 397976
rect 48148 397972 48154 397974
rect 90081 397971 90147 397974
rect 98637 398034 98703 398037
rect 99046 398034 99052 398036
rect 98637 398032 99052 398034
rect 98637 397976 98642 398032
rect 98698 397976 99052 398032
rect 98637 397974 99052 397976
rect 98637 397971 98703 397974
rect 99046 397972 99052 397974
rect 99116 397972 99122 398036
rect -960 397490 480 397580
rect 3141 397490 3207 397493
rect -960 397488 3207 397490
rect -960 397432 3146 397488
rect 3202 397432 3207 397488
rect -960 397430 3207 397432
rect -960 397340 480 397430
rect 3141 397427 3207 397430
rect 583520 391628 584960 391868
rect 103421 391234 103487 391237
rect 116209 391234 116275 391237
rect 103421 391232 116275 391234
rect 103421 391176 103426 391232
rect 103482 391176 116214 391232
rect 116270 391176 116275 391232
rect 103421 391174 116275 391176
rect 103421 391171 103487 391174
rect 116209 391171 116275 391174
rect 111006 390628 111012 390692
rect 111076 390690 111082 390692
rect 114185 390690 114251 390693
rect 111076 390688 114251 390690
rect 111076 390632 114190 390688
rect 114246 390632 114251 390688
rect 111076 390630 114251 390632
rect 111076 390628 111082 390630
rect 114185 390627 114251 390630
rect 53598 390492 53604 390556
rect 53668 390554 53674 390556
rect 57237 390554 57303 390557
rect 53668 390552 57303 390554
rect 53668 390496 57242 390552
rect 57298 390496 57303 390552
rect 53668 390494 57303 390496
rect 53668 390492 53674 390494
rect 57237 390491 57303 390494
rect 136582 390492 136588 390556
rect 136652 390554 136658 390556
rect 136909 390554 136975 390557
rect 136652 390552 136975 390554
rect 136652 390496 136914 390552
rect 136970 390496 136975 390552
rect 136652 390494 136975 390496
rect 136652 390492 136658 390494
rect 136909 390491 136975 390494
rect 96429 389874 96495 389877
rect 118734 389874 118740 389876
rect 96429 389872 118740 389874
rect 96429 389816 96434 389872
rect 96490 389816 118740 389872
rect 96429 389814 118740 389816
rect 96429 389811 96495 389814
rect 118734 389812 118740 389814
rect 118804 389812 118810 389876
rect 53598 389132 53604 389196
rect 53668 389194 53674 389196
rect 95877 389194 95943 389197
rect 96429 389194 96495 389197
rect 53668 389192 96495 389194
rect 53668 389136 95882 389192
rect 95938 389136 96434 389192
rect 96490 389136 96495 389192
rect 53668 389134 96495 389136
rect 53668 389132 53674 389134
rect 95877 389131 95943 389134
rect 96429 389131 96495 389134
rect 114921 389194 114987 389197
rect 268326 389194 268332 389196
rect 114921 389192 268332 389194
rect 114921 389136 114926 389192
rect 114982 389136 268332 389192
rect 114921 389134 268332 389136
rect 114921 389131 114987 389134
rect 268326 389132 268332 389134
rect 268396 389132 268402 389196
rect 58525 388380 58591 388381
rect 52310 388316 52316 388380
rect 52380 388378 52386 388380
rect 58525 388378 58572 388380
rect 52380 388376 58572 388378
rect 58636 388378 58642 388380
rect 115841 388378 115907 388381
rect 129825 388378 129891 388381
rect 130377 388378 130443 388381
rect 52380 388320 58530 388376
rect 52380 388318 58572 388320
rect 52380 388316 52386 388318
rect 58525 388316 58572 388318
rect 58636 388318 58718 388378
rect 115841 388376 130443 388378
rect 115841 388320 115846 388376
rect 115902 388320 129830 388376
rect 129886 388320 130382 388376
rect 130438 388320 130443 388376
rect 115841 388318 130443 388320
rect 58636 388316 58642 388318
rect 58525 388315 58591 388316
rect 115841 388315 115907 388318
rect 129825 388315 129891 388318
rect 130377 388315 130443 388318
rect 114185 387970 114251 387973
rect 119286 387970 119292 387972
rect 114185 387968 119292 387970
rect 114185 387912 114190 387968
rect 114246 387912 119292 387968
rect 114185 387910 119292 387912
rect 114185 387907 114251 387910
rect 119286 387908 119292 387910
rect 119356 387908 119362 387972
rect 73521 387834 73587 387837
rect 73797 387834 73863 387837
rect 119470 387834 119476 387836
rect 73521 387832 119476 387834
rect 73521 387776 73526 387832
rect 73582 387776 73802 387832
rect 73858 387776 119476 387832
rect 73521 387774 119476 387776
rect 73521 387771 73587 387774
rect 73797 387771 73863 387774
rect 119470 387772 119476 387774
rect 119540 387772 119546 387836
rect 50286 387636 50292 387700
rect 50356 387698 50362 387700
rect 50889 387698 50955 387701
rect 50356 387696 50955 387698
rect 50356 387640 50894 387696
rect 50950 387640 50955 387696
rect 50356 387638 50955 387640
rect 50356 387636 50362 387638
rect 50889 387635 50955 387638
rect 122097 387698 122163 387701
rect 122833 387698 122899 387701
rect 122097 387696 122899 387698
rect 122097 387640 122102 387696
rect 122158 387640 122838 387696
rect 122894 387640 122899 387696
rect 122097 387638 122899 387640
rect 122097 387635 122163 387638
rect 122833 387635 122899 387638
rect 54886 386956 54892 387020
rect 54956 387018 54962 387020
rect 80145 387018 80211 387021
rect 54956 387016 80211 387018
rect 54956 386960 80150 387016
rect 80206 386960 80211 387016
rect 54956 386958 80211 386960
rect 54956 386956 54962 386958
rect 80145 386955 80211 386958
rect 111793 387018 111859 387021
rect 120022 387018 120028 387020
rect 111793 387016 120028 387018
rect 111793 386960 111798 387016
rect 111854 386960 120028 387016
rect 111793 386958 120028 386960
rect 111793 386955 111859 386958
rect 120022 386956 120028 386958
rect 120092 386956 120098 387020
rect 120257 387018 120323 387021
rect 299606 387018 299612 387020
rect 120257 387016 299612 387018
rect 120257 386960 120262 387016
rect 120318 386960 299612 387016
rect 120257 386958 299612 386960
rect 120257 386955 120323 386958
rect 299606 386956 299612 386958
rect 299676 386956 299682 387020
rect 122097 386610 122163 386613
rect 122598 386610 122604 386612
rect 122097 386608 122604 386610
rect 122097 386552 122102 386608
rect 122158 386552 122604 386608
rect 122097 386550 122604 386552
rect 122097 386547 122163 386550
rect 122598 386548 122604 386550
rect 122668 386548 122674 386612
rect 76649 386474 76715 386477
rect 262990 386474 262996 386476
rect 76649 386472 262996 386474
rect 76649 386416 76654 386472
rect 76710 386416 262996 386472
rect 76649 386414 262996 386416
rect 76649 386411 76715 386414
rect 262990 386412 262996 386414
rect 263060 386412 263066 386476
rect 117681 386338 117747 386341
rect 117814 386338 117820 386340
rect 117681 386336 117820 386338
rect 117681 386280 117686 386336
rect 117742 386280 117820 386336
rect 117681 386278 117820 386280
rect 117681 386275 117747 386278
rect 117814 386276 117820 386278
rect 117884 386276 117890 386340
rect 134517 385658 134583 385661
rect 143533 385658 143599 385661
rect 122790 385656 143599 385658
rect 70166 385250 70226 385628
rect 122790 385600 134522 385656
rect 134578 385600 143538 385656
rect 143594 385600 143599 385656
rect 122790 385598 143599 385600
rect 112805 385386 112871 385389
rect 122790 385386 122850 385598
rect 134517 385595 134583 385598
rect 143533 385595 143599 385598
rect 112805 385384 122850 385386
rect 112805 385328 112810 385384
rect 112866 385328 122850 385384
rect 112805 385326 122850 385328
rect 112805 385323 112871 385326
rect 115790 385250 115796 385252
rect 64830 385190 74550 385250
rect 61694 385052 61700 385116
rect 61764 385114 61770 385116
rect 64830 385114 64890 385190
rect 61764 385054 64890 385114
rect 74490 385114 74550 385190
rect 103470 385190 115796 385250
rect 103470 385114 103530 385190
rect 115790 385188 115796 385190
rect 115860 385188 115866 385252
rect 74490 385054 103530 385114
rect 61764 385052 61770 385054
rect 117998 384978 118004 384980
rect 65926 384780 65932 384844
rect 65996 384842 66002 384844
rect 70166 384842 70226 384948
rect 115828 384918 118004 384978
rect 117998 384916 118004 384918
rect 118068 384978 118074 384980
rect 118509 384978 118575 384981
rect 118068 384976 118575 384978
rect 118068 384920 118514 384976
rect 118570 384920 118575 384976
rect 118068 384918 118575 384920
rect 118068 384916 118074 384918
rect 118509 384915 118575 384918
rect 65996 384782 70226 384842
rect 65996 384780 66002 384782
rect -960 384284 480 384524
rect 115790 384508 115796 384572
rect 115860 384570 115866 384572
rect 259494 384570 259500 384572
rect 115860 384510 259500 384570
rect 115860 384508 115866 384510
rect 259494 384508 259500 384510
rect 259564 384508 259570 384572
rect 115798 384026 115858 384268
rect 115933 384026 115999 384029
rect 115798 384024 115999 384026
rect 115798 383968 115938 384024
rect 115994 383968 115999 384024
rect 115798 383966 115999 383968
rect 115933 383963 115999 383966
rect 65885 383892 65951 383893
rect 65885 383890 65932 383892
rect 65840 383888 65932 383890
rect 65840 383832 65890 383888
rect 65840 383830 65932 383832
rect 65885 383828 65932 383830
rect 65996 383828 66002 383892
rect 65885 383827 65951 383828
rect 118601 383618 118667 383621
rect 115828 383616 118667 383618
rect 68737 383482 68803 383485
rect 70166 383482 70226 383588
rect 115828 383560 118606 383616
rect 118662 383560 118667 383616
rect 115828 383558 118667 383560
rect 118601 383555 118667 383558
rect 68737 383480 70226 383482
rect 68737 383424 68742 383480
rect 68798 383424 70226 383480
rect 68737 383422 70226 383424
rect 68737 383419 68803 383422
rect 67633 382530 67699 382533
rect 70166 382530 70226 382908
rect 67633 382528 70226 382530
rect 67633 382472 67638 382528
rect 67694 382472 70226 382528
rect 67633 382470 70226 382472
rect 67633 382467 67699 382470
rect 122046 382258 122052 382260
rect 70166 381578 70226 382228
rect 115828 382198 122052 382258
rect 122046 382196 122052 382198
rect 122116 382196 122122 382260
rect 118601 381578 118667 381581
rect 64830 381518 70226 381578
rect 115828 381576 118667 381578
rect 115828 381520 118606 381576
rect 118662 381520 118667 381576
rect 115828 381518 118667 381520
rect 61878 380972 61884 381036
rect 61948 381034 61954 381036
rect 62982 381034 62988 381036
rect 61948 380974 62988 381034
rect 61948 380972 61954 380974
rect 62982 380972 62988 380974
rect 63052 381034 63058 381036
rect 64830 381034 64890 381518
rect 118601 381515 118667 381518
rect 63052 380974 64890 381034
rect 63052 380972 63058 380974
rect 118601 380898 118667 380901
rect 115828 380896 118667 380898
rect 67633 380762 67699 380765
rect 70166 380762 70226 380868
rect 115828 380840 118606 380896
rect 118662 380840 118667 380896
rect 115828 380838 118667 380840
rect 118601 380835 118667 380838
rect 67633 380760 70226 380762
rect 67633 380704 67638 380760
rect 67694 380704 70226 380760
rect 67633 380702 70226 380704
rect 67633 380699 67699 380702
rect 49601 380218 49667 380221
rect 55070 380218 55076 380220
rect 49601 380216 55076 380218
rect 49601 380160 49606 380216
rect 49662 380160 55076 380216
rect 49601 380158 55076 380160
rect 49601 380155 49667 380158
rect 55070 380156 55076 380158
rect 55140 380218 55146 380220
rect 64781 380218 64847 380221
rect 55140 380216 64847 380218
rect 55140 380160 64786 380216
rect 64842 380160 64847 380216
rect 122189 380218 122255 380221
rect 129774 380218 129780 380220
rect 122189 380216 129780 380218
rect 55140 380158 64847 380160
rect 55140 380156 55146 380158
rect 64781 380155 64847 380158
rect 67633 379810 67699 379813
rect 70166 379810 70226 380188
rect 122189 380160 122194 380216
rect 122250 380160 129780 380216
rect 122189 380158 129780 380160
rect 122189 380155 122255 380158
rect 129774 380156 129780 380158
rect 129844 380156 129850 380220
rect 67633 379808 70226 379810
rect 67633 379752 67638 379808
rect 67694 379752 70226 379808
rect 67633 379750 70226 379752
rect 67633 379747 67699 379750
rect 61694 379612 61700 379676
rect 61764 379674 61770 379676
rect 66662 379674 66668 379676
rect 61764 379614 66668 379674
rect 61764 379612 61770 379614
rect 66662 379612 66668 379614
rect 66732 379674 66738 379676
rect 66732 379614 70226 379674
rect 66732 379612 66738 379614
rect 70166 379508 70226 379614
rect 117313 379538 117379 379541
rect 118325 379538 118391 379541
rect 115828 379536 118391 379538
rect 115828 379480 117318 379536
rect 117374 379480 118330 379536
rect 118386 379480 118391 379536
rect 115828 379478 118391 379480
rect 117313 379475 117379 379478
rect 118325 379475 118391 379478
rect 123017 378994 123083 378997
rect 123334 378994 123340 378996
rect 123017 378992 123340 378994
rect 123017 378936 123022 378992
rect 123078 378936 123340 378992
rect 123017 378934 123340 378936
rect 123017 378931 123083 378934
rect 123334 378932 123340 378934
rect 123404 378932 123410 378996
rect 118601 378858 118667 378861
rect 115828 378856 118667 378858
rect 115828 378800 118606 378856
rect 118662 378800 118667 378856
rect 115828 378798 118667 378800
rect 118601 378795 118667 378798
rect 580349 378450 580415 378453
rect 583520 378450 584960 378540
rect 580349 378448 584960 378450
rect 580349 378392 580354 378448
rect 580410 378392 584960 378448
rect 580349 378390 584960 378392
rect 580349 378387 580415 378390
rect 64830 378254 70226 378314
rect 583520 378300 584960 378390
rect 64830 378181 64890 378254
rect 64781 378176 64890 378181
rect 64781 378120 64786 378176
rect 64842 378120 64890 378176
rect 70166 378148 70226 378254
rect 118601 378178 118667 378181
rect 115828 378176 118667 378178
rect 64781 378118 64890 378120
rect 115828 378120 118606 378176
rect 118662 378120 118667 378176
rect 115828 378118 118667 378120
rect 64781 378115 64847 378118
rect 118601 378115 118667 378118
rect 59077 378042 59143 378045
rect 60590 378042 60596 378044
rect 59077 378040 60596 378042
rect 59077 377984 59082 378040
rect 59138 377984 60596 378040
rect 59077 377982 60596 377984
rect 59077 377979 59143 377982
rect 60590 377980 60596 377982
rect 60660 377980 60666 378044
rect 53741 377770 53807 377773
rect 69974 377770 69980 377772
rect 53741 377768 69980 377770
rect 53741 377712 53746 377768
rect 53802 377712 69980 377768
rect 53741 377710 69980 377712
rect 53741 377707 53807 377710
rect 69974 377708 69980 377710
rect 70044 377708 70050 377772
rect 67633 377362 67699 377365
rect 70166 377362 70226 377468
rect 67633 377360 70226 377362
rect 67633 377304 67638 377360
rect 67694 377304 70226 377360
rect 67633 377302 70226 377304
rect 67633 377299 67699 377302
rect 64830 376894 70226 376954
rect 60590 376756 60596 376820
rect 60660 376818 60666 376820
rect 64830 376818 64890 376894
rect 60660 376758 64890 376818
rect 70166 376788 70226 376894
rect 117078 376818 117084 376820
rect 115828 376758 117084 376818
rect 60660 376756 60666 376758
rect 117078 376756 117084 376758
rect 117148 376818 117154 376820
rect 118417 376818 118483 376821
rect 117148 376816 118483 376818
rect 117148 376760 118422 376816
rect 118478 376760 118483 376816
rect 117148 376758 118483 376760
rect 117148 376756 117154 376758
rect 118417 376755 118483 376758
rect 117773 376138 117839 376141
rect 115828 376136 117839 376138
rect 115828 376080 117778 376136
rect 117834 376080 117839 376136
rect 115828 376078 117839 376080
rect 117773 376075 117839 376078
rect 69105 376002 69171 376005
rect 69105 376000 70226 376002
rect 69105 375944 69110 376000
rect 69166 375944 70226 376000
rect 69105 375942 70226 375944
rect 69105 375939 69171 375942
rect 70166 375428 70226 375942
rect 118601 375458 118667 375461
rect 115828 375456 118667 375458
rect 115828 375400 118606 375456
rect 118662 375400 118667 375456
rect 115828 375398 118667 375400
rect 118601 375395 118667 375398
rect 69105 374642 69171 374645
rect 70166 374642 70226 374748
rect 69105 374640 70226 374642
rect 69105 374584 69110 374640
rect 69166 374584 70226 374640
rect 69105 374582 70226 374584
rect 146201 374642 146267 374645
rect 262806 374642 262812 374644
rect 146201 374640 262812 374642
rect 146201 374584 146206 374640
rect 146262 374584 262812 374640
rect 146201 374582 262812 374584
rect 69105 374579 69171 374582
rect 146201 374579 146267 374582
rect 262806 374580 262812 374582
rect 262876 374580 262882 374644
rect 67633 374506 67699 374509
rect 67633 374504 70226 374506
rect 67633 374448 67638 374504
rect 67694 374448 70226 374504
rect 67633 374446 70226 374448
rect 67633 374443 67699 374446
rect 70166 374068 70226 374446
rect 118601 374098 118667 374101
rect 115828 374096 118667 374098
rect 115828 374040 118606 374096
rect 118662 374040 118667 374096
rect 115828 374038 118667 374040
rect 118601 374035 118667 374038
rect 65885 373962 65951 373965
rect 66110 373962 66116 373964
rect 65885 373960 66116 373962
rect 65885 373904 65890 373960
rect 65946 373904 66116 373960
rect 65885 373902 66116 373904
rect 65885 373899 65951 373902
rect 66110 373900 66116 373902
rect 66180 373900 66186 373964
rect 118601 373418 118667 373421
rect 115828 373416 118667 373418
rect 115828 373360 118606 373416
rect 118662 373360 118667 373416
rect 115828 373358 118667 373360
rect 118601 373355 118667 373358
rect 151813 373282 151879 373285
rect 287646 373282 287652 373284
rect 151813 373280 287652 373282
rect 151813 373224 151818 373280
rect 151874 373224 287652 373280
rect 151813 373222 287652 373224
rect 151813 373219 151879 373222
rect 287646 373220 287652 373222
rect 287716 373220 287722 373284
rect 66110 372812 66116 372876
rect 66180 372874 66186 372876
rect 66180 372814 70226 372874
rect 66180 372812 66186 372814
rect 70166 372708 70226 372814
rect 117814 372738 117820 372740
rect 115828 372678 117820 372738
rect 117814 372676 117820 372678
rect 117884 372738 117890 372740
rect 123334 372738 123340 372740
rect 117884 372678 123340 372738
rect 117884 372676 117890 372678
rect 123334 372676 123340 372678
rect 123404 372676 123410 372740
rect 67725 371922 67791 371925
rect 70166 371922 70226 372028
rect 67725 371920 70226 371922
rect 67725 371864 67730 371920
rect 67786 371864 70226 371920
rect 67725 371862 70226 371864
rect 67725 371859 67791 371862
rect 67633 371786 67699 371789
rect 67633 371784 70226 371786
rect 67633 371728 67638 371784
rect 67694 371728 70226 371784
rect 67633 371726 70226 371728
rect 67633 371723 67699 371726
rect -960 371378 480 371468
rect 3233 371378 3299 371381
rect -960 371376 3299 371378
rect -960 371320 3238 371376
rect 3294 371320 3299 371376
rect 70166 371348 70226 371726
rect 116209 371378 116275 371381
rect 335854 371378 335860 371380
rect 115828 371376 335860 371378
rect -960 371318 3299 371320
rect 115828 371320 116214 371376
rect 116270 371320 335860 371376
rect 115828 371318 335860 371320
rect -960 371228 480 371318
rect 3233 371315 3299 371318
rect 116209 371315 116275 371318
rect 335854 371316 335860 371318
rect 335924 371316 335930 371380
rect 116209 370698 116275 370701
rect 117865 370698 117931 370701
rect 115828 370696 117931 370698
rect 115828 370640 116214 370696
rect 116270 370640 117870 370696
rect 117926 370640 117931 370696
rect 115828 370638 117931 370640
rect 116209 370635 116275 370638
rect 117865 370635 117931 370638
rect 56317 370562 56383 370565
rect 69054 370562 69060 370564
rect 56317 370560 69060 370562
rect 56317 370504 56322 370560
rect 56378 370504 69060 370560
rect 56317 370502 69060 370504
rect 56317 370499 56383 370502
rect 69054 370500 69060 370502
rect 69124 370500 69130 370564
rect 119470 370500 119476 370564
rect 119540 370562 119546 370564
rect 301497 370562 301563 370565
rect 119540 370560 301563 370562
rect 119540 370504 301502 370560
rect 301558 370504 301563 370560
rect 119540 370502 301563 370504
rect 119540 370500 119546 370502
rect 301497 370499 301563 370502
rect 116025 370426 116091 370429
rect 115798 370424 116091 370426
rect 115798 370368 116030 370424
rect 116086 370368 116091 370424
rect 115798 370366 116091 370368
rect 68369 370154 68435 370157
rect 69197 370154 69263 370157
rect 68369 370152 70226 370154
rect 68369 370096 68374 370152
rect 68430 370096 69202 370152
rect 69258 370096 70226 370152
rect 68369 370094 70226 370096
rect 68369 370091 68435 370094
rect 69197 370091 69263 370094
rect 70166 369988 70226 370094
rect 115798 370018 115858 370366
rect 116025 370363 116091 370366
rect 118049 370018 118115 370021
rect 115798 370016 118115 370018
rect 115798 369988 118054 370016
rect 115828 369960 118054 369988
rect 118110 369960 118115 370016
rect 115828 369958 118115 369960
rect 118049 369955 118115 369958
rect 67357 369746 67423 369749
rect 67357 369744 70226 369746
rect 67357 369688 67362 369744
rect 67418 369688 70226 369744
rect 67357 369686 70226 369688
rect 67357 369683 67423 369686
rect 70166 369308 70226 369686
rect 67633 369066 67699 369069
rect 67633 369064 70226 369066
rect 67633 369008 67638 369064
rect 67694 369008 70226 369064
rect 67633 369006 70226 369008
rect 67633 369003 67699 369006
rect 70166 368628 70226 369006
rect 119286 369004 119292 369068
rect 119356 369066 119362 369068
rect 272517 369066 272583 369069
rect 119356 369064 272583 369066
rect 119356 369008 272522 369064
rect 272578 369008 272583 369064
rect 119356 369006 272583 369008
rect 119356 369004 119362 369006
rect 272517 369003 272583 369006
rect 117313 368658 117379 368661
rect 115828 368656 117379 368658
rect 115828 368600 117318 368656
rect 117374 368600 117379 368656
rect 115828 368598 117379 368600
rect 117313 368595 117379 368598
rect 62982 368324 62988 368388
rect 63052 368386 63058 368388
rect 64137 368386 64203 368389
rect 63052 368384 70226 368386
rect 63052 368328 64142 368384
rect 64198 368328 70226 368384
rect 63052 368326 70226 368328
rect 63052 368324 63058 368326
rect 64137 368323 64203 368326
rect 70166 367268 70226 368326
rect 122046 368324 122052 368388
rect 122116 368386 122122 368388
rect 150525 368386 150591 368389
rect 150985 368386 151051 368389
rect 122116 368384 151051 368386
rect 122116 368328 150530 368384
rect 150586 368328 150990 368384
rect 151046 368328 151051 368384
rect 122116 368326 151051 368328
rect 122116 368324 122122 368326
rect 150525 368323 150591 368326
rect 150985 368323 151051 368326
rect 117313 367978 117379 367981
rect 115828 367976 117379 367978
rect 115828 367920 117318 367976
rect 117374 367920 117379 367976
rect 115828 367918 117379 367920
rect 117313 367915 117379 367918
rect 150985 367706 151051 367709
rect 283557 367706 283623 367709
rect 150985 367704 283623 367706
rect 150985 367648 150990 367704
rect 151046 367648 283562 367704
rect 283618 367648 283623 367704
rect 150985 367646 283623 367648
rect 150985 367643 151051 367646
rect 283557 367643 283623 367646
rect 117405 367298 117471 367301
rect 115828 367296 117471 367298
rect 115828 367240 117410 367296
rect 117466 367240 117471 367296
rect 115828 367238 117471 367240
rect 117405 367235 117471 367238
rect 67633 366482 67699 366485
rect 70166 366482 70226 366588
rect 67633 366480 70226 366482
rect 67633 366424 67638 366480
rect 67694 366424 70226 366480
rect 67633 366422 70226 366424
rect 67633 366419 67699 366422
rect 68001 366074 68067 366077
rect 68870 366074 68876 366076
rect 68001 366072 68876 366074
rect 68001 366016 68006 366072
rect 68062 366016 68876 366072
rect 68001 366014 68876 366016
rect 68001 366011 68067 366014
rect 68870 366012 68876 366014
rect 68940 366074 68946 366076
rect 68940 366014 70226 366074
rect 68940 366012 68946 366014
rect 70166 365908 70226 366014
rect 117313 365938 117379 365941
rect 115828 365936 117379 365938
rect 115828 365880 117318 365936
rect 117374 365880 117379 365936
rect 115828 365878 117379 365880
rect 117313 365875 117379 365878
rect 117313 365258 117379 365261
rect 115828 365256 117379 365258
rect 115828 365200 117318 365256
rect 117374 365200 117379 365256
rect 115828 365198 117379 365200
rect 117313 365195 117379 365198
rect 580257 365122 580323 365125
rect 583520 365122 584960 365212
rect 580257 365120 584960 365122
rect 580257 365064 580262 365120
rect 580318 365064 584960 365120
rect 580257 365062 584960 365064
rect 580257 365059 580323 365062
rect 583520 364972 584960 365062
rect 118918 364850 118924 364852
rect 115798 364790 118924 364850
rect 115798 364548 115858 364790
rect 118918 364788 118924 364790
rect 118988 364850 118994 364852
rect 119061 364850 119127 364853
rect 118988 364848 119127 364850
rect 118988 364792 119066 364848
rect 119122 364792 119127 364848
rect 118988 364790 119127 364792
rect 118988 364788 118994 364790
rect 119061 364787 119127 364790
rect 67633 364442 67699 364445
rect 70166 364442 70226 364548
rect 67633 364440 70226 364442
rect 67633 364384 67638 364440
rect 67694 364384 70226 364440
rect 67633 364382 70226 364384
rect 67633 364379 67699 364382
rect 67725 364306 67791 364309
rect 67725 364304 70226 364306
rect 67725 364248 67730 364304
rect 67786 364248 70226 364304
rect 67725 364246 70226 364248
rect 67725 364243 67791 364246
rect 70166 363868 70226 364246
rect 67633 363626 67699 363629
rect 67633 363624 70226 363626
rect 67633 363568 67638 363624
rect 67694 363568 70226 363624
rect 67633 363566 70226 363568
rect 67633 363563 67699 363566
rect 70166 363188 70226 363566
rect 117681 363218 117747 363221
rect 115828 363216 117747 363218
rect 115828 363160 117686 363216
rect 117742 363160 117747 363216
rect 115828 363158 117747 363160
rect 117681 363155 117747 363158
rect 117313 362538 117379 362541
rect 115828 362536 117379 362538
rect 67449 362402 67515 362405
rect 70166 362402 70226 362508
rect 115828 362480 117318 362536
rect 117374 362480 117379 362536
rect 115828 362478 117379 362480
rect 117313 362475 117379 362478
rect 67449 362400 70226 362402
rect 67449 362344 67454 362400
rect 67510 362344 70226 362400
rect 67449 362342 70226 362344
rect 67449 362339 67515 362342
rect 117313 361858 117379 361861
rect 115828 361856 117379 361858
rect 115828 361800 117318 361856
rect 117374 361800 117379 361856
rect 115828 361798 117379 361800
rect 117313 361795 117379 361798
rect 117313 361178 117379 361181
rect 115828 361176 117379 361178
rect 65926 360980 65932 361044
rect 65996 361042 66002 361044
rect 70166 361042 70226 361148
rect 115828 361120 117318 361176
rect 117374 361120 117379 361176
rect 115828 361118 117379 361120
rect 117313 361115 117379 361118
rect 65996 360982 70226 361042
rect 65996 360980 66002 360982
rect 67633 360906 67699 360909
rect 67633 360904 70226 360906
rect 67633 360848 67638 360904
rect 67694 360848 70226 360904
rect 67633 360846 70226 360848
rect 67633 360843 67699 360846
rect 70166 360468 70226 360846
rect 33777 360090 33843 360093
rect 65374 360090 65380 360092
rect 33777 360088 65380 360090
rect 33777 360032 33782 360088
rect 33838 360032 65380 360088
rect 33777 360030 65380 360032
rect 33777 360027 33843 360030
rect 65374 360028 65380 360030
rect 65444 360090 65450 360092
rect 65926 360090 65932 360092
rect 65444 360030 65932 360090
rect 65444 360028 65450 360030
rect 65926 360028 65932 360030
rect 65996 360028 66002 360092
rect 118877 359818 118943 359821
rect 115828 359816 118943 359818
rect 67633 359274 67699 359277
rect 70166 359274 70226 359788
rect 115828 359760 118882 359816
rect 118938 359760 118943 359816
rect 115828 359758 118943 359760
rect 118877 359755 118943 359758
rect 115289 359546 115355 359549
rect 115289 359544 115490 359546
rect 115289 359488 115294 359544
rect 115350 359488 115490 359544
rect 115289 359486 115490 359488
rect 115289 359483 115355 359486
rect 67633 359272 70226 359274
rect 67633 359216 67638 359272
rect 67694 359216 70226 359272
rect 67633 359214 70226 359216
rect 115430 359274 115490 359486
rect 115430 359214 115858 359274
rect 67633 359211 67699 359214
rect 115430 359108 115490 359214
rect 115798 359138 115858 359214
rect 117865 359138 117931 359141
rect 115798 359136 117931 359138
rect 115798 359108 117870 359136
rect 115828 359080 117870 359108
rect 117926 359080 117931 359136
rect 115828 359078 117931 359080
rect 117865 359075 117931 359078
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect 118601 358458 118667 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect 115828 358456 118667 358458
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 67725 358186 67791 358189
rect 70166 358186 70226 358428
rect 115828 358400 118606 358456
rect 118662 358400 118667 358456
rect 115828 358398 118667 358400
rect 118601 358395 118667 358398
rect 67725 358184 70226 358186
rect 67725 358128 67730 358184
rect 67786 358128 70226 358184
rect 67725 358126 70226 358128
rect 67725 358123 67791 358126
rect 67633 358050 67699 358053
rect 67633 358048 70226 358050
rect 67633 357992 67638 358048
rect 67694 357992 70226 358048
rect 67633 357990 70226 357992
rect 67633 357987 67699 357990
rect 70166 357748 70226 357990
rect 45369 357506 45435 357509
rect 68134 357506 68140 357508
rect 45369 357504 68140 357506
rect 45369 357448 45374 357504
rect 45430 357448 68140 357504
rect 45369 357446 68140 357448
rect 45369 357443 45435 357446
rect 67774 357370 67834 357446
rect 68134 357444 68140 357446
rect 68204 357444 68210 357508
rect 67774 357310 70226 357370
rect 70166 357068 70226 357310
rect 116117 357098 116183 357101
rect 118141 357098 118207 357101
rect 115828 357096 118207 357098
rect 115828 357040 116122 357096
rect 116178 357040 118146 357096
rect 118202 357040 118207 357096
rect 115828 357038 118207 357040
rect 116117 357035 116183 357038
rect 118141 357035 118207 357038
rect 118601 356418 118667 356421
rect 115828 356416 118667 356418
rect 115828 356360 118606 356416
rect 118662 356360 118667 356416
rect 115828 356358 118667 356360
rect 118601 356355 118667 356358
rect 67633 355874 67699 355877
rect 67633 355872 70226 355874
rect 67633 355816 67638 355872
rect 67694 355816 70226 355872
rect 67633 355814 70226 355816
rect 67633 355811 67699 355814
rect 70166 355708 70226 355814
rect 117589 355738 117655 355741
rect 118601 355738 118667 355741
rect 115828 355736 118667 355738
rect 115828 355680 117594 355736
rect 117650 355680 118606 355736
rect 118662 355680 118667 355736
rect 115828 355678 118667 355680
rect 117589 355675 117655 355678
rect 118601 355675 118667 355678
rect 67725 355466 67791 355469
rect 67725 355464 70226 355466
rect 67725 355408 67730 355464
rect 67786 355408 70226 355464
rect 67725 355406 70226 355408
rect 67725 355403 67791 355406
rect 70166 355028 70226 355406
rect 118601 354378 118667 354381
rect 115828 354376 118667 354378
rect 67633 353834 67699 353837
rect 70166 353834 70226 354348
rect 115828 354320 118606 354376
rect 118662 354320 118667 354376
rect 115828 354318 118667 354320
rect 118601 354315 118667 354318
rect 67633 353832 70226 353834
rect 67633 353776 67638 353832
rect 67694 353776 70226 353832
rect 67633 353774 70226 353776
rect 67633 353771 67699 353774
rect 118509 353698 118575 353701
rect 115828 353696 118575 353698
rect 115828 353640 118514 353696
rect 118570 353640 118575 353696
rect 115828 353638 118575 353640
rect 118509 353635 118575 353638
rect 68921 353154 68987 353157
rect 68921 353152 70226 353154
rect 68921 353096 68926 353152
rect 68982 353096 70226 353152
rect 68921 353094 70226 353096
rect 68921 353091 68987 353094
rect 70166 352988 70226 353094
rect 118601 353018 118667 353021
rect 115828 353016 118667 353018
rect 115828 352960 118606 353016
rect 118662 352960 118667 353016
rect 115828 352958 118667 352960
rect 118601 352955 118667 352958
rect 67633 352610 67699 352613
rect 67633 352608 70226 352610
rect 67633 352552 67638 352608
rect 67694 352552 70226 352608
rect 67633 352550 70226 352552
rect 67633 352547 67699 352550
rect 70166 352308 70226 352550
rect 579613 351930 579679 351933
rect 583520 351930 584960 352020
rect 579613 351928 584960 351930
rect 579613 351872 579618 351928
rect 579674 351872 584960 351928
rect 579613 351870 584960 351872
rect 579613 351867 579679 351870
rect 583520 351780 584960 351870
rect 117497 351658 117563 351661
rect 118601 351658 118667 351661
rect 115828 351656 118667 351658
rect 67909 351250 67975 351253
rect 68737 351250 68803 351253
rect 70166 351250 70226 351628
rect 115828 351600 117502 351656
rect 117558 351600 118606 351656
rect 118662 351600 118667 351656
rect 115828 351598 118667 351600
rect 117497 351595 117563 351598
rect 118601 351595 118667 351598
rect 67909 351248 70226 351250
rect 67909 351192 67914 351248
rect 67970 351192 68742 351248
rect 68798 351192 70226 351248
rect 67909 351190 70226 351192
rect 67909 351187 67975 351190
rect 68737 351187 68803 351190
rect 118049 350978 118115 350981
rect 115828 350976 118115 350978
rect 115828 350920 118054 350976
rect 118110 350920 118115 350976
rect 115828 350918 118115 350920
rect 118049 350915 118115 350918
rect 67633 350434 67699 350437
rect 67633 350432 70226 350434
rect 67633 350376 67638 350432
rect 67694 350376 70226 350432
rect 67633 350374 70226 350376
rect 67633 350371 67699 350374
rect 70166 350268 70226 350374
rect 118601 350298 118667 350301
rect 115828 350296 118667 350298
rect 115828 350240 118606 350296
rect 118662 350240 118667 350296
rect 115828 350238 118667 350240
rect 118601 350235 118667 350238
rect 68369 349754 68435 349757
rect 68829 349754 68895 349757
rect 68369 349752 70226 349754
rect 68369 349696 68374 349752
rect 68430 349696 68834 349752
rect 68890 349696 70226 349752
rect 68369 349694 70226 349696
rect 68369 349691 68435 349694
rect 68829 349691 68895 349694
rect 70166 349588 70226 349694
rect 123334 349692 123340 349756
rect 123404 349754 123410 349756
rect 337377 349754 337443 349757
rect 123404 349752 337443 349754
rect 123404 349696 337382 349752
rect 337438 349696 337443 349752
rect 123404 349694 337443 349696
rect 123404 349692 123410 349694
rect 337377 349691 337443 349694
rect 115289 349210 115355 349213
rect 115289 349208 115490 349210
rect 115289 349152 115294 349208
rect 115350 349152 115490 349208
rect 115289 349150 115490 349152
rect 115289 349147 115355 349150
rect 67633 349074 67699 349077
rect 115430 349074 115490 349150
rect 67633 349072 70226 349074
rect 67633 349016 67638 349072
rect 67694 349016 70226 349072
rect 67633 349014 70226 349016
rect 115430 349014 115858 349074
rect 67633 349011 67699 349014
rect 70166 348908 70226 349014
rect 115798 348938 115858 349014
rect 117865 348938 117931 348941
rect 115798 348936 117931 348938
rect 115798 348908 117870 348936
rect 115828 348880 117870 348908
rect 117926 348880 117931 348936
rect 115828 348878 117931 348880
rect 117865 348875 117931 348878
rect 118601 348258 118667 348261
rect 115828 348256 118667 348258
rect 115828 348200 118606 348256
rect 118662 348200 118667 348256
rect 115828 348198 118667 348200
rect 118601 348195 118667 348198
rect 33041 347714 33107 347717
rect 57094 347714 57100 347716
rect 33041 347712 57100 347714
rect 33041 347656 33046 347712
rect 33102 347656 57100 347712
rect 33041 347654 57100 347656
rect 33041 347651 33107 347654
rect 57094 347652 57100 347654
rect 57164 347714 57170 347716
rect 57881 347714 57947 347717
rect 57164 347712 57947 347714
rect 57164 347656 57886 347712
rect 57942 347656 57947 347712
rect 57164 347654 57947 347656
rect 57164 347652 57170 347654
rect 57881 347651 57947 347654
rect 117405 347578 117471 347581
rect 115828 347576 117471 347578
rect 67633 347170 67699 347173
rect 70166 347170 70226 347548
rect 115828 347520 117410 347576
rect 117466 347520 117471 347576
rect 115828 347518 117471 347520
rect 117405 347515 117471 347518
rect 67633 347168 70226 347170
rect 67633 347112 67638 347168
rect 67694 347112 70226 347168
rect 67633 347110 70226 347112
rect 67633 347107 67699 347110
rect 67725 347034 67791 347037
rect 67725 347032 70226 347034
rect 67725 346976 67730 347032
rect 67786 346976 70226 347032
rect 67725 346974 70226 346976
rect 67725 346971 67791 346974
rect 70166 346868 70226 346974
rect 68185 346354 68251 346357
rect 68185 346352 70226 346354
rect 68185 346296 68190 346352
rect 68246 346296 70226 346352
rect 68185 346294 70226 346296
rect 68185 346291 68251 346294
rect 70166 345946 70226 346294
rect 118509 346218 118575 346221
rect 115828 346216 118575 346218
rect 115828 346160 118514 346216
rect 118570 346160 118575 346216
rect 115828 346158 118575 346160
rect 118509 346155 118575 346158
rect 70301 345946 70367 345949
rect 70166 345944 70367 345946
rect 70166 345888 70306 345944
rect 70362 345888 70367 345944
rect 70166 345886 70367 345888
rect 70301 345883 70367 345886
rect 118601 345538 118667 345541
rect 115828 345536 118667 345538
rect -960 345402 480 345492
rect 115828 345480 118606 345536
rect 118662 345480 118667 345536
rect 115828 345478 118667 345480
rect 118601 345475 118667 345478
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 68645 344994 68711 344997
rect 68645 344992 70226 344994
rect 68645 344936 68650 344992
rect 68706 344936 70226 344992
rect 68645 344934 70226 344936
rect 68645 344931 68711 344934
rect 70166 344828 70226 344934
rect 118601 344858 118667 344861
rect 115828 344856 118667 344858
rect 115828 344800 118606 344856
rect 118662 344800 118667 344856
rect 115828 344798 118667 344800
rect 118601 344795 118667 344798
rect 67633 343770 67699 343773
rect 70166 343770 70226 344148
rect 67633 343768 70226 343770
rect 67633 343712 67638 343768
rect 67694 343712 70226 343768
rect 67633 343710 70226 343712
rect 67633 343707 67699 343710
rect 118601 343498 118667 343501
rect 115828 343496 118667 343498
rect 67633 342954 67699 342957
rect 70166 342954 70226 343468
rect 115828 343440 118606 343496
rect 118662 343440 118667 343496
rect 115828 343438 118667 343440
rect 118601 343435 118667 343438
rect 67633 342952 70226 342954
rect 67633 342896 67638 342952
rect 67694 342896 70226 342952
rect 67633 342894 70226 342896
rect 67633 342891 67699 342894
rect 117773 342818 117839 342821
rect 115828 342816 117839 342818
rect 115828 342760 117778 342816
rect 117834 342760 117839 342816
rect 115828 342758 117839 342760
rect 117773 342755 117839 342758
rect 126145 342412 126211 342413
rect 126094 342410 126100 342412
rect 126054 342350 126100 342410
rect 126164 342408 126211 342412
rect 126206 342352 126211 342408
rect 126094 342348 126100 342350
rect 126164 342348 126211 342352
rect 126145 342347 126211 342348
rect 118601 342138 118667 342141
rect 115828 342136 118667 342138
rect 70350 341733 70410 342108
rect 115828 342080 118606 342136
rect 118662 342080 118667 342136
rect 115828 342078 118667 342080
rect 118601 342075 118667 342078
rect 68645 341730 68711 341733
rect 70350 341730 70459 341733
rect 68645 341728 70459 341730
rect 68645 341672 68650 341728
rect 68706 341672 70398 341728
rect 70454 341672 70459 341728
rect 68645 341670 70459 341672
rect 68645 341667 68711 341670
rect 70393 341667 70459 341670
rect 67541 341594 67607 341597
rect 67541 341592 70594 341594
rect 67541 341536 67546 341592
rect 67602 341536 70594 341592
rect 67541 341534 70594 341536
rect 67541 341531 67607 341534
rect 70534 341052 70594 341534
rect 70526 340988 70532 341052
rect 70596 340988 70602 341052
rect 117497 340778 117563 340781
rect 115828 340776 117563 340778
rect 70534 340237 70594 340748
rect 115828 340720 117502 340776
rect 117558 340720 117563 340776
rect 115828 340718 117563 340720
rect 117497 340715 117563 340718
rect 67909 340234 67975 340237
rect 70485 340234 70594 340237
rect 67909 340232 70594 340234
rect 67909 340176 67914 340232
rect 67970 340176 70490 340232
rect 70546 340176 70594 340232
rect 67909 340174 70594 340176
rect 67909 340171 67975 340174
rect 70485 340171 70551 340174
rect 117313 340098 117379 340101
rect 118417 340098 118483 340101
rect 115828 340096 118483 340098
rect 115828 340040 117318 340096
rect 117374 340040 118422 340096
rect 118478 340040 118483 340096
rect 115828 340038 118483 340040
rect 117313 340035 117379 340038
rect 118417 340035 118483 340038
rect 55029 339690 55095 339693
rect 75913 339690 75979 339693
rect 77109 339690 77175 339693
rect 55029 339688 77175 339690
rect 55029 339632 55034 339688
rect 55090 339632 75918 339688
rect 75974 339632 77114 339688
rect 77170 339632 77175 339688
rect 55029 339630 77175 339632
rect 55029 339627 55095 339630
rect 75913 339627 75979 339630
rect 77109 339627 77175 339630
rect 109953 339418 110019 339421
rect 128670 339418 128676 339420
rect 109953 339416 128676 339418
rect 109953 339360 109958 339416
rect 110014 339360 128676 339416
rect 109953 339358 128676 339360
rect 109953 339355 110019 339358
rect 128670 339356 128676 339358
rect 128740 339356 128746 339420
rect 583520 338452 584960 338692
rect 55070 338132 55076 338196
rect 55140 338194 55146 338196
rect 102133 338194 102199 338197
rect 55140 338192 102199 338194
rect 55140 338136 102138 338192
rect 102194 338136 102199 338192
rect 55140 338134 102199 338136
rect 55140 338132 55146 338134
rect 102133 338131 102199 338134
rect 57830 337996 57836 338060
rect 57900 338058 57906 338060
rect 58985 338058 59051 338061
rect 57900 338056 59051 338058
rect 57900 338000 58990 338056
rect 59046 338000 59051 338056
rect 57900 337998 59051 338000
rect 57900 337996 57906 337998
rect 58985 337995 59051 337998
rect 73889 338058 73955 338061
rect 74441 338058 74507 338061
rect 119337 338058 119403 338061
rect 73889 338056 119403 338058
rect 73889 338000 73894 338056
rect 73950 338000 74446 338056
rect 74502 338000 119342 338056
rect 119398 338000 119403 338056
rect 73889 337998 119403 338000
rect 73889 337995 73955 337998
rect 74441 337995 74507 337998
rect 119337 337995 119403 337998
rect 120022 337996 120028 338060
rect 120092 338058 120098 338060
rect 120165 338058 120231 338061
rect 120092 338056 120231 338058
rect 120092 338000 120170 338056
rect 120226 338000 120231 338056
rect 120092 337998 120231 338000
rect 120092 337996 120098 337998
rect 120165 337995 120231 337998
rect 70526 335956 70532 336020
rect 70596 336018 70602 336020
rect 293217 336018 293283 336021
rect 70596 336016 293283 336018
rect 70596 335960 293222 336016
rect 293278 335960 293283 336016
rect 70596 335958 293283 335960
rect 70596 335956 70602 335958
rect 293217 335955 293283 335958
rect 91001 333298 91067 333301
rect 258390 333298 258396 333300
rect 91001 333296 258396 333298
rect 91001 333240 91006 333296
rect 91062 333240 258396 333296
rect 91001 333238 258396 333240
rect 91001 333235 91067 333238
rect 258390 333236 258396 333238
rect 258460 333236 258466 333300
rect -960 332196 480 332436
rect 54886 332012 54892 332076
rect 54956 332074 54962 332076
rect 55029 332074 55095 332077
rect 54956 332072 55095 332074
rect 54956 332016 55034 332072
rect 55090 332016 55095 332072
rect 54956 332014 55095 332016
rect 54956 332012 54962 332014
rect 55029 332011 55095 332014
rect 66069 331802 66135 331805
rect 270534 331802 270540 331804
rect 66069 331800 270540 331802
rect 66069 331744 66074 331800
rect 66130 331744 270540 331800
rect 66069 331742 270540 331744
rect 66069 331739 66135 331742
rect 270534 331740 270540 331742
rect 270604 331740 270610 331804
rect 63309 330578 63375 330581
rect 173014 330578 173020 330580
rect 63309 330576 173020 330578
rect 63309 330520 63314 330576
rect 63370 330520 173020 330576
rect 63309 330518 173020 330520
rect 63309 330515 63375 330518
rect 173014 330516 173020 330518
rect 173084 330516 173090 330580
rect 68870 330380 68876 330444
rect 68940 330442 68946 330444
rect 280889 330442 280955 330445
rect 68940 330440 280955 330442
rect 68940 330384 280894 330440
rect 280950 330384 280955 330440
rect 68940 330382 280955 330384
rect 68940 330380 68946 330382
rect 280889 330379 280955 330382
rect 68737 329082 68803 329085
rect 269062 329082 269068 329084
rect 68737 329080 269068 329082
rect 68737 329024 68742 329080
rect 68798 329024 269068 329080
rect 68737 329022 269068 329024
rect 68737 329019 68803 329022
rect 269062 329020 269068 329022
rect 269132 329020 269138 329084
rect 70894 327660 70900 327724
rect 70964 327722 70970 327724
rect 117313 327722 117379 327725
rect 70964 327720 117379 327722
rect 70964 327664 117318 327720
rect 117374 327664 117379 327720
rect 70964 327662 117379 327664
rect 70964 327660 70970 327662
rect 117313 327659 117379 327662
rect 137093 326498 137159 326501
rect 302182 326498 302188 326500
rect 137093 326496 302188 326498
rect 137093 326440 137098 326496
rect 137154 326440 302188 326496
rect 137093 326438 302188 326440
rect 137093 326435 137159 326438
rect 302182 326436 302188 326438
rect 302252 326436 302258 326500
rect 65374 326300 65380 326364
rect 65444 326362 65450 326364
rect 263542 326362 263548 326364
rect 65444 326302 263548 326362
rect 65444 326300 65450 326302
rect 263542 326300 263548 326302
rect 263612 326300 263618 326364
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect 68829 322146 68895 322149
rect 309726 322146 309732 322148
rect 68829 322144 309732 322146
rect 68829 322088 68834 322144
rect 68890 322088 309732 322144
rect 68829 322086 309732 322088
rect 68829 322083 68895 322086
rect 309726 322084 309732 322086
rect 309796 322084 309802 322148
rect 131665 319426 131731 319429
rect 334014 319426 334020 319428
rect 131665 319424 334020 319426
rect -960 319290 480 319380
rect 131665 319368 131670 319424
rect 131726 319368 334020 319424
rect 131665 319366 334020 319368
rect 131665 319363 131731 319366
rect 334014 319364 334020 319366
rect 334084 319364 334090 319428
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 75269 318066 75335 318069
rect 342294 318066 342300 318068
rect 75269 318064 342300 318066
rect 75269 318008 75274 318064
rect 75330 318008 342300 318064
rect 75269 318006 342300 318008
rect 75269 318003 75335 318006
rect 342294 318004 342300 318006
rect 342364 318004 342370 318068
rect 79409 316706 79475 316709
rect 340822 316706 340828 316708
rect 79409 316704 340828 316706
rect 79409 316648 79414 316704
rect 79470 316648 340828 316704
rect 79409 316646 340828 316648
rect 79409 316643 79475 316646
rect 340822 316644 340828 316646
rect 340892 316644 340898 316708
rect 124397 316026 124463 316029
rect 124806 316026 124812 316028
rect 124397 316024 124812 316026
rect 124397 315968 124402 316024
rect 124458 315968 124812 316024
rect 124397 315966 124812 315968
rect 124397 315963 124463 315966
rect 124806 315964 124812 315966
rect 124876 315964 124882 316028
rect 74441 315346 74507 315349
rect 118734 315346 118740 315348
rect 74441 315344 118740 315346
rect 74441 315288 74446 315344
rect 74502 315288 118740 315344
rect 74441 315286 118740 315288
rect 74441 315283 74507 315286
rect 118734 315284 118740 315286
rect 118804 315284 118810 315348
rect 124806 314740 124812 314804
rect 124876 314802 124882 314804
rect 125726 314802 125732 314804
rect 124876 314742 125732 314802
rect 124876 314740 124882 314742
rect 125726 314740 125732 314742
rect 125796 314740 125802 314804
rect 122557 314260 122623 314261
rect 122557 314256 122604 314260
rect 122668 314258 122674 314260
rect 122557 314200 122562 314256
rect 122557 314196 122604 314200
rect 122668 314198 122714 314258
rect 122668 314196 122674 314198
rect 122557 314195 122623 314196
rect 127249 312490 127315 312493
rect 266854 312490 266860 312492
rect 127249 312488 266860 312490
rect 127249 312432 127254 312488
rect 127310 312432 266860 312488
rect 127249 312430 266860 312432
rect 127249 312427 127315 312430
rect 266854 312428 266860 312430
rect 266924 312428 266930 312492
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 118877 307732 118943 307733
rect 118877 307728 118924 307732
rect 118988 307730 118994 307732
rect 118877 307672 118882 307728
rect 118877 307668 118924 307672
rect 118988 307670 119034 307730
rect 118988 307668 118994 307670
rect 118877 307667 118943 307668
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 70393 302290 70459 302293
rect 322974 302290 322980 302292
rect 70393 302288 322980 302290
rect 70393 302232 70398 302288
rect 70454 302232 322980 302288
rect 70393 302230 322980 302232
rect 70393 302227 70459 302230
rect 322974 302228 322980 302230
rect 323044 302228 323050 302292
rect 42609 302154 42675 302157
rect 65609 302154 65675 302157
rect 66161 302154 66227 302157
rect 42609 302152 66227 302154
rect 42609 302096 42614 302152
rect 42670 302096 65614 302152
rect 65670 302096 66166 302152
rect 66222 302096 66227 302152
rect 42609 302094 66227 302096
rect 42609 302091 42675 302094
rect 65609 302091 65675 302094
rect 66161 302091 66227 302094
rect 71037 301474 71103 301477
rect 122598 301474 122604 301476
rect 71037 301472 122604 301474
rect 71037 301416 71042 301472
rect 71098 301416 122604 301472
rect 71037 301414 122604 301416
rect 71037 301411 71103 301414
rect 122598 301412 122604 301414
rect 122668 301412 122674 301476
rect 73245 300930 73311 300933
rect 330334 300930 330340 300932
rect 73245 300928 330340 300930
rect 73245 300872 73250 300928
rect 73306 300872 330340 300928
rect 73245 300870 330340 300872
rect 73245 300867 73311 300870
rect 330334 300868 330340 300870
rect 330404 300868 330410 300932
rect 68921 299570 68987 299573
rect 326654 299570 326660 299572
rect 68921 299568 326660 299570
rect 68921 299512 68926 299568
rect 68982 299512 326660 299568
rect 68921 299510 326660 299512
rect 68921 299507 68987 299510
rect 326654 299508 326660 299510
rect 326724 299508 326730 299572
rect 66110 298692 66116 298756
rect 66180 298754 66186 298756
rect 298134 298754 298140 298756
rect 66180 298694 298140 298754
rect 66180 298692 66186 298694
rect 298134 298692 298140 298694
rect 298204 298692 298210 298756
rect 580901 298754 580967 298757
rect 583520 298754 584960 298844
rect 580901 298752 584960 298754
rect 580901 298696 580906 298752
rect 580962 298696 584960 298752
rect 580901 298694 584960 298696
rect 580901 298691 580967 298694
rect 583520 298604 584960 298694
rect 101581 297394 101647 297397
rect 131113 297394 131179 297397
rect 101581 297392 132510 297394
rect 101581 297336 101586 297392
rect 101642 297336 131118 297392
rect 131174 297336 132510 297392
rect 101581 297334 132510 297336
rect 101581 297331 101647 297334
rect 131113 297331 131179 297334
rect 132450 296986 132510 297334
rect 133873 296986 133939 296989
rect 132450 296984 133939 296986
rect 132450 296928 133878 296984
rect 133934 296928 133939 296984
rect 132450 296926 133939 296928
rect 133873 296923 133939 296926
rect 113173 296850 113239 296853
rect 342253 296850 342319 296853
rect 113173 296848 342319 296850
rect 113173 296792 113178 296848
rect 113234 296792 342258 296848
rect 342314 296792 342319 296848
rect 113173 296790 342319 296792
rect 113173 296787 113239 296790
rect 342253 296787 342319 296790
rect 59118 295972 59124 296036
rect 59188 296034 59194 296036
rect 96705 296034 96771 296037
rect 59188 296032 96771 296034
rect 59188 295976 96710 296032
rect 96766 295976 96771 296032
rect 59188 295974 96771 295976
rect 59188 295972 59194 295974
rect 96705 295971 96771 295974
rect 119889 295626 119955 295629
rect 121678 295626 121684 295628
rect 119889 295624 121684 295626
rect 119889 295568 119894 295624
rect 119950 295568 121684 295624
rect 119889 295566 121684 295568
rect 119889 295563 119955 295566
rect 121678 295564 121684 295566
rect 121748 295564 121754 295628
rect 100937 295490 101003 295493
rect 255262 295490 255268 295492
rect 100937 295488 255268 295490
rect 100937 295432 100942 295488
rect 100998 295432 255268 295488
rect 100937 295430 255268 295432
rect 100937 295427 101003 295430
rect 255262 295428 255268 295430
rect 255332 295428 255338 295492
rect 111241 295354 111307 295357
rect 340873 295354 340939 295357
rect 111241 295352 340939 295354
rect 111241 295296 111246 295352
rect 111302 295296 340878 295352
rect 340934 295296 340939 295352
rect 111241 295294 340939 295296
rect 111241 295291 111307 295294
rect 340873 295291 340939 295294
rect 58566 294476 58572 294540
rect 58636 294538 58642 294540
rect 91277 294538 91343 294541
rect 58636 294536 91343 294538
rect 58636 294480 91282 294536
rect 91338 294480 91343 294536
rect 58636 294478 91343 294480
rect 58636 294476 58642 294478
rect 91277 294475 91343 294478
rect 95785 294266 95851 294269
rect 178769 294266 178835 294269
rect 95785 294264 178835 294266
rect 95785 294208 95790 294264
rect 95846 294208 178774 294264
rect 178830 294208 178835 294264
rect 95785 294206 178835 294208
rect 95785 294203 95851 294206
rect 178769 294203 178835 294206
rect 75821 294130 75887 294133
rect 188429 294130 188495 294133
rect 75821 294128 188495 294130
rect 75821 294072 75826 294128
rect 75882 294072 188434 294128
rect 188490 294072 188495 294128
rect 75821 294070 188495 294072
rect 75821 294067 75887 294070
rect 188429 294067 188495 294070
rect 108021 293994 108087 293997
rect 313917 293994 313983 293997
rect 108021 293992 313983 293994
rect 108021 293936 108026 293992
rect 108082 293936 313922 293992
rect 313978 293936 313983 293992
rect 108021 293934 313983 293936
rect 108021 293931 108087 293934
rect 313917 293931 313983 293934
rect -960 293178 480 293268
rect 3049 293178 3115 293181
rect -960 293176 3115 293178
rect -960 293120 3054 293176
rect 3110 293120 3115 293176
rect -960 293118 3115 293120
rect -960 293028 480 293118
rect 3049 293115 3115 293118
rect 57237 292906 57303 292909
rect 118325 292906 118391 292909
rect 57237 292904 118391 292906
rect 57237 292848 57242 292904
rect 57298 292848 118330 292904
rect 118386 292848 118391 292904
rect 57237 292846 118391 292848
rect 57237 292843 57303 292846
rect 118325 292843 118391 292846
rect 111885 292770 111951 292773
rect 202229 292770 202295 292773
rect 111885 292768 202295 292770
rect 111885 292712 111890 292768
rect 111946 292712 202234 292768
rect 202290 292712 202295 292768
rect 111885 292710 202295 292712
rect 111885 292707 111951 292710
rect 202229 292707 202295 292710
rect 97073 292634 97139 292637
rect 436093 292634 436159 292637
rect 97073 292632 436159 292634
rect 97073 292576 97078 292632
rect 97134 292576 436098 292632
rect 436154 292576 436159 292632
rect 97073 292574 436159 292576
rect 97073 292571 97139 292574
rect 436093 292571 436159 292574
rect 71129 292362 71195 292365
rect 70718 292360 71195 292362
rect 70718 292304 71134 292360
rect 71190 292304 71195 292360
rect 70718 292302 71195 292304
rect 70718 291788 70778 292302
rect 71129 292299 71195 292302
rect 114553 291954 114619 291957
rect 152457 291954 152523 291957
rect 114553 291952 152523 291954
rect 114553 291896 114558 291952
rect 114614 291896 152462 291952
rect 152518 291896 152523 291952
rect 114553 291894 152523 291896
rect 114553 291891 114619 291894
rect 152457 291891 152523 291894
rect 121545 291818 121611 291821
rect 119876 291816 121611 291818
rect 119876 291760 121550 291816
rect 121606 291760 121611 291816
rect 119876 291758 121611 291760
rect 121545 291755 121611 291758
rect 69982 291214 70226 291274
rect 67725 291138 67791 291141
rect 69982 291138 70042 291214
rect 67725 291136 70042 291138
rect 67725 291080 67730 291136
rect 67786 291080 70042 291136
rect 70166 291108 70226 291214
rect 121545 291138 121611 291141
rect 119876 291136 121611 291138
rect 67725 291078 70042 291080
rect 119876 291080 121550 291136
rect 121606 291080 121611 291136
rect 119876 291078 121611 291080
rect 67725 291075 67791 291078
rect 121545 291075 121611 291078
rect 67633 290866 67699 290869
rect 67633 290864 70226 290866
rect 67633 290808 67638 290864
rect 67694 290808 70226 290864
rect 67633 290806 70226 290808
rect 67633 290803 67699 290806
rect 70166 290428 70226 290806
rect 119846 289914 119906 290428
rect 252502 289914 252508 289916
rect 119846 289854 252508 289914
rect 252502 289852 252508 289854
rect 252572 289852 252578 289916
rect 67633 289234 67699 289237
rect 70166 289234 70226 289748
rect 119294 289508 119354 289748
rect 119286 289444 119292 289508
rect 119356 289506 119362 289508
rect 122373 289506 122439 289509
rect 119356 289504 122439 289506
rect 119356 289448 122378 289504
rect 122434 289448 122439 289504
rect 119356 289446 122439 289448
rect 119356 289444 119362 289446
rect 122373 289443 122439 289446
rect 67633 289232 70226 289234
rect 67633 289176 67638 289232
rect 67694 289176 70226 289232
rect 67633 289174 70226 289176
rect 67633 289171 67699 289174
rect 121729 289098 121795 289101
rect 119876 289096 121795 289098
rect 69841 288826 69907 288829
rect 70350 288826 70410 289068
rect 119876 289040 121734 289096
rect 121790 289040 121795 289096
rect 119876 289038 121795 289040
rect 121729 289035 121795 289038
rect 69841 288824 70410 288826
rect 69841 288768 69846 288824
rect 69902 288768 70410 288824
rect 69841 288766 70410 288768
rect 69841 288763 69907 288766
rect 121821 288418 121887 288421
rect 119876 288416 121887 288418
rect 67817 288146 67883 288149
rect 70350 288146 70410 288388
rect 119876 288360 121826 288416
rect 121882 288360 121887 288416
rect 119876 288358 121887 288360
rect 121821 288355 121887 288358
rect 67817 288144 70410 288146
rect 67817 288088 67822 288144
rect 67878 288088 70410 288144
rect 67817 288086 70410 288088
rect 67817 288083 67883 288086
rect 121545 287738 121611 287741
rect 119876 287736 121611 287738
rect 67817 287466 67883 287469
rect 70166 287466 70226 287708
rect 119876 287680 121550 287736
rect 121606 287680 121611 287736
rect 119876 287678 121611 287680
rect 121545 287675 121611 287678
rect 67817 287464 70226 287466
rect 67817 287408 67822 287464
rect 67878 287408 70226 287464
rect 67817 287406 70226 287408
rect 67817 287403 67883 287406
rect 67541 287058 67607 287061
rect 69982 287058 70226 287070
rect 121545 287058 121611 287061
rect 67541 287056 70226 287058
rect 67541 287000 67546 287056
rect 67602 287010 70226 287056
rect 119876 287056 121611 287058
rect 67602 287000 70042 287010
rect 67541 286998 70042 287000
rect 119876 287000 121550 287056
rect 121606 287000 121611 287056
rect 119876 286998 121611 287000
rect 67541 286995 67607 286998
rect 121545 286995 121611 286998
rect 69105 286786 69171 286789
rect 69105 286784 70226 286786
rect 69105 286728 69110 286784
rect 69166 286728 70226 286784
rect 69105 286726 70226 286728
rect 69105 286723 69171 286726
rect 70166 286348 70226 286726
rect 121545 286378 121611 286381
rect 119876 286376 121611 286378
rect 119876 286320 121550 286376
rect 121606 286320 121611 286376
rect 119876 286318 121611 286320
rect 121545 286315 121611 286318
rect 68921 286106 68987 286109
rect 68921 286104 70226 286106
rect 68921 286048 68926 286104
rect 68982 286048 70226 286104
rect 68921 286046 70226 286048
rect 68921 286043 68987 286046
rect 70166 285668 70226 286046
rect 122741 285698 122807 285701
rect 119876 285696 122807 285698
rect 119876 285640 122746 285696
rect 122802 285640 122807 285696
rect 119876 285638 122807 285640
rect 122741 285635 122807 285638
rect 70526 285364 70532 285428
rect 70596 285364 70602 285428
rect 70534 284988 70594 285364
rect 583520 285276 584960 285516
rect 121545 285018 121611 285021
rect 119876 285016 121611 285018
rect 119876 284960 121550 285016
rect 121606 284960 121611 285016
rect 119876 284958 121611 284960
rect 121545 284955 121611 284958
rect 68277 284474 68343 284477
rect 68277 284472 70226 284474
rect 68277 284416 68282 284472
rect 68338 284416 70226 284472
rect 68277 284414 70226 284416
rect 68277 284411 68343 284414
rect 70166 284308 70226 284414
rect 121637 284340 121703 284341
rect 121637 284338 121684 284340
rect 119876 284336 121684 284338
rect 121748 284338 121754 284340
rect 119876 284280 121642 284336
rect 119876 284278 121684 284280
rect 121637 284276 121684 284278
rect 121748 284278 121830 284338
rect 121748 284276 121754 284278
rect 121637 284275 121703 284276
rect 68921 283794 68987 283797
rect 68921 283792 70226 283794
rect 68921 283736 68926 283792
rect 68982 283736 70226 283792
rect 68921 283734 70226 283736
rect 68921 283731 68987 283734
rect 70166 283628 70226 283734
rect 121545 283658 121611 283661
rect 119876 283656 121611 283658
rect 119876 283600 121550 283656
rect 121606 283600 121611 283656
rect 119876 283598 121611 283600
rect 121545 283595 121611 283598
rect 144177 283522 144243 283525
rect 256734 283522 256740 283524
rect 144177 283520 256740 283522
rect 144177 283464 144182 283520
rect 144238 283464 256740 283520
rect 144177 283462 256740 283464
rect 144177 283459 144243 283462
rect 256734 283460 256740 283462
rect 256804 283460 256810 283524
rect 67633 283386 67699 283389
rect 67633 283384 70226 283386
rect 67633 283328 67638 283384
rect 67694 283328 70226 283384
rect 67633 283326 70226 283328
rect 67633 283323 67699 283326
rect 70166 282948 70226 283326
rect 121545 282978 121611 282981
rect 119876 282976 121611 282978
rect 119876 282920 121550 282976
rect 121606 282920 121611 282976
rect 119876 282918 121611 282920
rect 121545 282915 121611 282918
rect 121637 282298 121703 282301
rect 119876 282296 121703 282298
rect 119876 282240 121642 282296
rect 121698 282240 121703 282296
rect 119876 282238 121703 282240
rect 121637 282235 121703 282238
rect 69013 282162 69079 282165
rect 69013 282160 70226 282162
rect 69013 282104 69018 282160
rect 69074 282104 70226 282160
rect 69013 282102 70226 282104
rect 69013 282099 69079 282102
rect 70166 281588 70226 282102
rect 121545 281618 121611 281621
rect 119876 281616 121611 281618
rect 119876 281560 121550 281616
rect 121606 281560 121611 281616
rect 119876 281558 121611 281560
rect 121545 281555 121611 281558
rect 121637 280938 121703 280941
rect 119876 280936 121703 280938
rect 67725 280530 67791 280533
rect 70166 280530 70226 280908
rect 119876 280880 121642 280936
rect 121698 280880 121703 280936
rect 119876 280878 121703 280880
rect 121637 280875 121703 280878
rect 67725 280528 70226 280530
rect 67725 280472 67730 280528
rect 67786 280472 70226 280528
rect 67725 280470 70226 280472
rect 67725 280467 67791 280470
rect 67633 280394 67699 280397
rect 67633 280392 70226 280394
rect 67633 280336 67638 280392
rect 67694 280336 70226 280392
rect 67633 280334 70226 280336
rect 67633 280331 67699 280334
rect 70166 280228 70226 280334
rect 121545 280258 121611 280261
rect 119876 280256 121611 280258
rect -960 279972 480 280212
rect 119876 280200 121550 280256
rect 121606 280200 121611 280256
rect 119876 280198 121611 280200
rect 121545 280195 121611 280198
rect 68001 279714 68067 279717
rect 69054 279714 69060 279716
rect 68001 279712 69060 279714
rect 68001 279656 68006 279712
rect 68062 279656 69060 279712
rect 68001 279654 69060 279656
rect 68001 279651 68067 279654
rect 69054 279652 69060 279654
rect 69124 279714 69130 279716
rect 69124 279654 70226 279714
rect 69124 279652 69130 279654
rect 70166 279548 70226 279654
rect 121637 279578 121703 279581
rect 119876 279576 121703 279578
rect 119876 279520 121642 279576
rect 121698 279520 121703 279576
rect 119876 279518 121703 279520
rect 121637 279515 121703 279518
rect 67633 279306 67699 279309
rect 67633 279304 70226 279306
rect 67633 279248 67638 279304
rect 67694 279248 70226 279304
rect 67633 279246 70226 279248
rect 67633 279243 67699 279246
rect 70166 278868 70226 279246
rect 121545 278898 121611 278901
rect 119876 278896 121611 278898
rect 119876 278840 121550 278896
rect 121606 278840 121611 278896
rect 119876 278838 121611 278840
rect 121545 278835 121611 278838
rect 67725 277810 67791 277813
rect 70166 277810 70226 278188
rect 67725 277808 70226 277810
rect 67725 277752 67730 277808
rect 67786 277752 70226 277808
rect 67725 277750 70226 277752
rect 119846 277810 119906 278188
rect 327022 277810 327028 277812
rect 119846 277750 327028 277810
rect 67725 277747 67791 277750
rect 327022 277748 327028 277750
rect 327092 277748 327098 277812
rect 67633 277674 67699 277677
rect 67633 277672 70226 277674
rect 67633 277616 67638 277672
rect 67694 277616 70226 277672
rect 67633 277614 70226 277616
rect 67633 277611 67699 277614
rect 70166 277508 70226 277614
rect 121545 277538 121611 277541
rect 119876 277536 121611 277538
rect 119876 277480 121550 277536
rect 121606 277480 121611 277536
rect 119876 277478 121611 277480
rect 121545 277475 121611 277478
rect 121729 276858 121795 276861
rect 119876 276856 121795 276858
rect 67725 276450 67791 276453
rect 70166 276450 70226 276828
rect 119876 276800 121734 276856
rect 121790 276800 121795 276856
rect 119876 276798 121795 276800
rect 121729 276795 121795 276798
rect 67725 276448 70226 276450
rect 67725 276392 67730 276448
rect 67786 276392 70226 276448
rect 67725 276390 70226 276392
rect 67725 276387 67791 276390
rect 67633 276314 67699 276317
rect 67633 276312 70226 276314
rect 67633 276256 67638 276312
rect 67694 276256 70226 276312
rect 67633 276254 70226 276256
rect 67633 276251 67699 276254
rect 70166 276148 70226 276254
rect 121545 276178 121611 276181
rect 119876 276176 121611 276178
rect 119876 276120 121550 276176
rect 121606 276120 121611 276176
rect 119876 276118 121611 276120
rect 121545 276115 121611 276118
rect 121637 275498 121703 275501
rect 119876 275496 121703 275498
rect 67725 275226 67791 275229
rect 70166 275226 70226 275468
rect 119876 275440 121642 275496
rect 121698 275440 121703 275496
rect 119876 275438 121703 275440
rect 121637 275435 121703 275438
rect 67725 275224 70226 275226
rect 67725 275168 67730 275224
rect 67786 275168 70226 275224
rect 67725 275166 70226 275168
rect 67725 275163 67791 275166
rect 67633 274954 67699 274957
rect 67633 274952 70226 274954
rect 67633 274896 67638 274952
rect 67694 274896 70226 274952
rect 67633 274894 70226 274896
rect 67633 274891 67699 274894
rect 70166 274788 70226 274894
rect 121545 274818 121611 274821
rect 119876 274816 121611 274818
rect 119876 274760 121550 274816
rect 121606 274760 121611 274816
rect 119876 274758 121611 274760
rect 121545 274755 121611 274758
rect 68001 274274 68067 274277
rect 69013 274274 69079 274277
rect 68001 274272 70226 274274
rect 68001 274216 68006 274272
rect 68062 274216 69018 274272
rect 69074 274216 70226 274272
rect 68001 274214 70226 274216
rect 68001 274211 68067 274214
rect 69013 274211 69079 274214
rect 70166 274108 70226 274214
rect 121545 274138 121611 274141
rect 119876 274136 121611 274138
rect 119876 274080 121550 274136
rect 121606 274080 121611 274136
rect 119876 274078 121611 274080
rect 121545 274075 121611 274078
rect 67633 273594 67699 273597
rect 67633 273592 70226 273594
rect 67633 273536 67638 273592
rect 67694 273536 70226 273592
rect 67633 273534 70226 273536
rect 67633 273531 67699 273534
rect 70166 273428 70226 273534
rect 121545 273458 121611 273461
rect 119876 273456 121611 273458
rect 119876 273400 121550 273456
rect 121606 273400 121611 273456
rect 119876 273398 121611 273400
rect 121545 273395 121611 273398
rect 121545 272778 121611 272781
rect 119876 272776 121611 272778
rect 67633 272370 67699 272373
rect 70166 272370 70226 272748
rect 119876 272720 121550 272776
rect 121606 272720 121611 272776
rect 119876 272718 121611 272720
rect 121545 272715 121611 272718
rect 67633 272368 70226 272370
rect 67633 272312 67638 272368
rect 67694 272312 70226 272368
rect 67633 272310 70226 272312
rect 67633 272307 67699 272310
rect 68185 272234 68251 272237
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 68185 272232 70226 272234
rect 68185 272176 68190 272232
rect 68246 272176 70226 272232
rect 68185 272174 70226 272176
rect 68185 272171 68251 272174
rect 70166 272068 70226 272174
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 121545 272098 121611 272101
rect 119876 272096 121611 272098
rect 119876 272040 121550 272096
rect 121606 272040 121611 272096
rect 583520 272084 584960 272174
rect 119876 272038 121611 272040
rect 121545 272035 121611 272038
rect 121545 271418 121611 271421
rect 119876 271416 121611 271418
rect 67633 271010 67699 271013
rect 70166 271010 70226 271388
rect 119876 271360 121550 271416
rect 121606 271360 121611 271416
rect 119876 271358 121611 271360
rect 121545 271355 121611 271358
rect 67633 271008 70226 271010
rect 67633 270952 67638 271008
rect 67694 270952 70226 271008
rect 67633 270950 70226 270952
rect 67633 270947 67699 270950
rect 66897 270874 66963 270877
rect 66897 270872 70226 270874
rect 66897 270816 66902 270872
rect 66958 270816 70226 270872
rect 66897 270814 70226 270816
rect 66897 270811 66963 270814
rect 70166 270708 70226 270814
rect 121637 270058 121703 270061
rect 119876 270056 121703 270058
rect 67725 269650 67791 269653
rect 70166 269650 70226 270028
rect 119876 270000 121642 270056
rect 121698 270000 121703 270056
rect 119876 269998 121703 270000
rect 121637 269995 121703 269998
rect 67725 269648 70226 269650
rect 67725 269592 67730 269648
rect 67786 269592 70226 269648
rect 67725 269590 70226 269592
rect 67725 269587 67791 269590
rect 67633 269514 67699 269517
rect 67633 269512 70226 269514
rect 67633 269456 67638 269512
rect 67694 269456 70226 269512
rect 67633 269454 70226 269456
rect 67633 269451 67699 269454
rect 70166 269348 70226 269454
rect 121545 269378 121611 269381
rect 119876 269376 121611 269378
rect 119876 269320 121550 269376
rect 121606 269320 121611 269376
rect 119876 269318 121611 269320
rect 121545 269315 121611 269318
rect 121637 268698 121703 268701
rect 119876 268696 121703 268698
rect 67725 268290 67791 268293
rect 70166 268290 70226 268668
rect 119876 268640 121642 268696
rect 121698 268640 121703 268696
rect 119876 268638 121703 268640
rect 121637 268635 121703 268638
rect 67725 268288 70226 268290
rect 67725 268232 67730 268288
rect 67786 268232 70226 268288
rect 67725 268230 70226 268232
rect 67725 268227 67791 268230
rect 67633 268154 67699 268157
rect 67633 268152 70226 268154
rect 67633 268096 67638 268152
rect 67694 268096 70226 268152
rect 67633 268094 70226 268096
rect 67633 268091 67699 268094
rect 70166 267988 70226 268094
rect 121545 268018 121611 268021
rect 119876 268016 121611 268018
rect 119876 267960 121550 268016
rect 121606 267960 121611 268016
rect 119876 267958 121611 267960
rect 121545 267955 121611 267958
rect 121637 267338 121703 267341
rect 119876 267336 121703 267338
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 67633 267066 67699 267069
rect 70166 267066 70226 267308
rect 119876 267280 121642 267336
rect 121698 267280 121703 267336
rect 119876 267278 121703 267280
rect 121637 267275 121703 267278
rect 67633 267064 70226 267066
rect 67633 267008 67638 267064
rect 67694 267008 70226 267064
rect 67633 267006 70226 267008
rect 67633 267003 67699 267006
rect 121545 266658 121611 266661
rect 119876 266656 121611 266658
rect 67633 266386 67699 266389
rect 70350 266386 70410 266628
rect 119876 266600 121550 266656
rect 121606 266600 121611 266656
rect 119876 266598 121611 266600
rect 121545 266595 121611 266598
rect 67633 266384 70410 266386
rect 67633 266328 67638 266384
rect 67694 266328 70410 266384
rect 67633 266326 70410 266328
rect 67633 266323 67699 266326
rect 121637 265978 121703 265981
rect 119876 265976 121703 265978
rect 67725 265570 67791 265573
rect 70166 265570 70226 265948
rect 119876 265920 121642 265976
rect 121698 265920 121703 265976
rect 119876 265918 121703 265920
rect 121637 265915 121703 265918
rect 67725 265568 70226 265570
rect 67725 265512 67730 265568
rect 67786 265512 70226 265568
rect 67725 265510 70226 265512
rect 67725 265507 67791 265510
rect 67817 265434 67883 265437
rect 67817 265432 70226 265434
rect 67817 265376 67822 265432
rect 67878 265376 70226 265432
rect 67817 265374 70226 265376
rect 67817 265371 67883 265374
rect 70166 265268 70226 265374
rect 121545 265298 121611 265301
rect 119876 265296 121611 265298
rect 119876 265240 121550 265296
rect 121606 265240 121611 265296
rect 119876 265238 121611 265240
rect 121545 265235 121611 265238
rect 67633 264890 67699 264893
rect 67633 264888 70226 264890
rect 67633 264832 67638 264888
rect 67694 264832 70226 264888
rect 67633 264830 70226 264832
rect 67633 264827 67699 264830
rect 70166 264588 70226 264830
rect 121729 264618 121795 264621
rect 119876 264616 121795 264618
rect 119876 264560 121734 264616
rect 121790 264560 121795 264616
rect 119876 264558 121795 264560
rect 121729 264555 121795 264558
rect 121545 263938 121611 263941
rect 119876 263936 121611 263938
rect 67633 263666 67699 263669
rect 70166 263666 70226 263908
rect 119876 263880 121550 263936
rect 121606 263880 121611 263936
rect 119876 263878 121611 263880
rect 121545 263875 121611 263878
rect 67633 263664 70226 263666
rect 67633 263608 67638 263664
rect 67694 263608 70226 263664
rect 67633 263606 70226 263608
rect 67633 263603 67699 263606
rect 121545 263258 121611 263261
rect 119876 263256 121611 263258
rect 67725 262850 67791 262853
rect 70166 262850 70226 263228
rect 119876 263200 121550 263256
rect 121606 263200 121611 263256
rect 119876 263198 121611 263200
rect 121545 263195 121611 263198
rect 67725 262848 70226 262850
rect 67725 262792 67730 262848
rect 67786 262792 70226 262848
rect 67725 262790 70226 262792
rect 67725 262787 67791 262790
rect 121545 262578 121611 262581
rect 119876 262576 121611 262578
rect 67633 262306 67699 262309
rect 70166 262306 70226 262548
rect 119876 262520 121550 262576
rect 121606 262520 121611 262576
rect 119876 262518 121611 262520
rect 121545 262515 121611 262518
rect 67633 262304 70226 262306
rect 67633 262248 67638 262304
rect 67694 262248 70226 262304
rect 67633 262246 70226 262248
rect 67633 262243 67699 262246
rect 121729 261898 121795 261901
rect 119876 261896 121795 261898
rect 67725 261490 67791 261493
rect 70166 261490 70226 261868
rect 119876 261840 121734 261896
rect 121790 261840 121795 261896
rect 119876 261838 121795 261840
rect 121729 261835 121795 261838
rect 67725 261488 70226 261490
rect 67725 261432 67730 261488
rect 67786 261432 70226 261488
rect 67725 261430 70226 261432
rect 67725 261427 67791 261430
rect 121637 261218 121703 261221
rect 119876 261216 121703 261218
rect 67633 260946 67699 260949
rect 70350 260946 70410 261188
rect 119876 261160 121642 261216
rect 121698 261160 121703 261216
rect 119876 261158 121703 261160
rect 121637 261155 121703 261158
rect 67633 260944 70410 260946
rect 67633 260888 67638 260944
rect 67694 260888 70410 260944
rect 67633 260886 70410 260888
rect 67633 260883 67699 260886
rect 67633 260810 67699 260813
rect 67633 260808 70226 260810
rect 67633 260752 67638 260808
rect 67694 260752 70226 260808
rect 67633 260750 70226 260752
rect 67633 260747 67699 260750
rect 70166 260508 70226 260750
rect 121545 260538 121611 260541
rect 119876 260536 121611 260538
rect 119876 260480 121550 260536
rect 121606 260480 121611 260536
rect 119876 260478 121611 260480
rect 121545 260475 121611 260478
rect 121545 259858 121611 259861
rect 119876 259856 121611 259858
rect 67633 259586 67699 259589
rect 70350 259586 70410 259828
rect 119876 259800 121550 259856
rect 121606 259800 121611 259856
rect 119876 259798 121611 259800
rect 121545 259795 121611 259798
rect 67633 259584 70410 259586
rect 67633 259528 67638 259584
rect 67694 259528 70410 259584
rect 67633 259526 70410 259528
rect 67633 259523 67699 259526
rect 121545 259178 121611 259181
rect 119876 259176 121611 259178
rect 67725 258770 67791 258773
rect 70166 258770 70226 259148
rect 119876 259120 121550 259176
rect 121606 259120 121611 259176
rect 119876 259118 121611 259120
rect 121545 259115 121611 259118
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 67725 258768 70226 258770
rect 67725 258712 67730 258768
rect 67786 258712 70226 258768
rect 583520 258756 584960 258846
rect 67725 258710 70226 258712
rect 67725 258707 67791 258710
rect 121637 258498 121703 258501
rect 119876 258496 121703 258498
rect 67633 258226 67699 258229
rect 70350 258226 70410 258468
rect 119876 258440 121642 258496
rect 121698 258440 121703 258496
rect 119876 258438 121703 258440
rect 121637 258435 121703 258438
rect 67633 258224 70410 258226
rect 67633 258168 67638 258224
rect 67694 258168 70410 258224
rect 67633 258166 70410 258168
rect 67633 258163 67699 258166
rect 121637 257818 121703 257821
rect 119876 257816 121703 257818
rect 67909 257274 67975 257277
rect 69238 257274 69244 257276
rect 67909 257272 69244 257274
rect 67909 257216 67914 257272
rect 67970 257216 69244 257272
rect 67909 257214 69244 257216
rect 67909 257211 67975 257214
rect 69238 257212 69244 257214
rect 69308 257274 69314 257276
rect 70166 257274 70226 257788
rect 119876 257760 121642 257816
rect 121698 257760 121703 257816
rect 119876 257758 121703 257760
rect 121637 257755 121703 257758
rect 69308 257214 70226 257274
rect 69308 257212 69314 257214
rect 121545 257138 121611 257141
rect 119876 257136 121611 257138
rect 67633 256866 67699 256869
rect 70350 256866 70410 257108
rect 119876 257080 121550 257136
rect 121606 257080 121611 257136
rect 119876 257078 121611 257080
rect 121545 257075 121611 257078
rect 67633 256864 70410 256866
rect 67633 256808 67638 256864
rect 67694 256808 70410 256864
rect 67633 256806 70410 256808
rect 67633 256803 67699 256806
rect 120165 256458 120231 256461
rect 121637 256458 121703 256461
rect 119876 256456 121703 256458
rect 67633 255914 67699 255917
rect 70166 255914 70226 256428
rect 119876 256400 120170 256456
rect 120226 256400 121642 256456
rect 121698 256400 121703 256456
rect 119876 256398 121703 256400
rect 120165 256395 120231 256398
rect 121637 256395 121703 256398
rect 67633 255912 70226 255914
rect 67633 255856 67638 255912
rect 67694 255856 70226 255912
rect 67633 255854 70226 255856
rect 67633 255851 67699 255854
rect 67725 255370 67791 255373
rect 70166 255370 70226 255748
rect 67725 255368 70226 255370
rect 67725 255312 67730 255368
rect 67786 255312 70226 255368
rect 67725 255310 70226 255312
rect 119846 255370 119906 255748
rect 125726 255370 125732 255372
rect 119846 255310 125732 255370
rect 67725 255307 67791 255310
rect 125726 255308 125732 255310
rect 125796 255308 125802 255372
rect 67633 255234 67699 255237
rect 67633 255232 70226 255234
rect 67633 255176 67638 255232
rect 67694 255176 70226 255232
rect 67633 255174 70226 255176
rect 67633 255171 67699 255174
rect 70166 255068 70226 255174
rect 122281 255098 122347 255101
rect 119876 255096 122347 255098
rect 119876 255040 122286 255096
rect 122342 255040 122347 255096
rect 119876 255038 122347 255040
rect 122281 255035 122347 255038
rect 121545 254418 121611 254421
rect 119876 254416 121611 254418
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 67633 254010 67699 254013
rect 70166 254010 70226 254388
rect 119876 254360 121550 254416
rect 121606 254360 121611 254416
rect 119876 254358 121611 254360
rect 121545 254355 121611 254358
rect 67633 254008 70226 254010
rect 67633 253952 67638 254008
rect 67694 253952 70226 254008
rect 67633 253950 70226 253952
rect 67633 253947 67699 253950
rect 121545 253738 121611 253741
rect 119876 253736 121611 253738
rect 67633 253194 67699 253197
rect 70166 253194 70226 253708
rect 119876 253680 121550 253736
rect 121606 253680 121611 253736
rect 119876 253678 121611 253680
rect 121545 253675 121611 253678
rect 67633 253192 70226 253194
rect 67633 253136 67638 253192
rect 67694 253136 70226 253192
rect 67633 253134 70226 253136
rect 67633 253131 67699 253134
rect 121637 253058 121703 253061
rect 119876 253056 121703 253058
rect 69105 252650 69171 252653
rect 70166 252650 70226 253028
rect 119876 253000 121642 253056
rect 121698 253000 121703 253056
rect 119876 252998 121703 253000
rect 121637 252995 121703 252998
rect 69105 252648 70226 252650
rect 69105 252592 69110 252648
rect 69166 252592 70226 252648
rect 69105 252590 70226 252592
rect 69105 252587 69171 252590
rect 121545 252378 121611 252381
rect 119876 252376 121611 252378
rect 67725 251834 67791 251837
rect 70166 251834 70226 252348
rect 119876 252320 121550 252376
rect 121606 252320 121611 252376
rect 119876 252318 121611 252320
rect 121545 252315 121611 252318
rect 67725 251832 70226 251834
rect 67725 251776 67730 251832
rect 67786 251776 70226 251832
rect 67725 251774 70226 251776
rect 67725 251771 67791 251774
rect 121545 251698 121611 251701
rect 119876 251696 121611 251698
rect 67633 251426 67699 251429
rect 70350 251426 70410 251668
rect 119876 251640 121550 251696
rect 121606 251640 121611 251696
rect 119876 251638 121611 251640
rect 121545 251635 121611 251638
rect 67633 251424 70410 251426
rect 67633 251368 67638 251424
rect 67694 251368 70410 251424
rect 67633 251366 70410 251368
rect 67633 251363 67699 251366
rect 120165 251018 120231 251021
rect 122097 251018 122163 251021
rect 119876 251016 122163 251018
rect 68645 250474 68711 250477
rect 70166 250474 70226 250988
rect 119876 250960 120170 251016
rect 120226 250960 122102 251016
rect 122158 250960 122163 251016
rect 119876 250958 122163 250960
rect 120165 250955 120231 250958
rect 122097 250955 122163 250958
rect 68645 250472 70226 250474
rect 68645 250416 68650 250472
rect 68706 250416 70226 250472
rect 68645 250414 70226 250416
rect 68645 250411 68711 250414
rect 121545 250338 121611 250341
rect 119876 250336 121611 250338
rect 67633 249930 67699 249933
rect 70166 249930 70226 250308
rect 119876 250280 121550 250336
rect 121606 250280 121611 250336
rect 119876 250278 121611 250280
rect 121545 250275 121611 250278
rect 67633 249928 70226 249930
rect 67633 249872 67638 249928
rect 67694 249872 70226 249928
rect 67633 249870 70226 249872
rect 67633 249867 67699 249870
rect 122598 249658 122604 249660
rect 67725 249114 67791 249117
rect 70166 249114 70226 249628
rect 119876 249598 122604 249658
rect 122598 249596 122604 249598
rect 122668 249596 122674 249660
rect 67725 249112 70226 249114
rect 67725 249056 67730 249112
rect 67786 249056 70226 249112
rect 67725 249054 70226 249056
rect 67725 249051 67791 249054
rect 121545 248978 121611 248981
rect 119876 248976 121611 248978
rect 67633 248570 67699 248573
rect 70166 248570 70226 248948
rect 119876 248920 121550 248976
rect 121606 248920 121611 248976
rect 119876 248918 121611 248920
rect 121545 248915 121611 248918
rect 67633 248568 70226 248570
rect 67633 248512 67638 248568
rect 67694 248512 70226 248568
rect 67633 248510 70226 248512
rect 67633 248507 67699 248510
rect 121453 248298 121519 248301
rect 119876 248296 121519 248298
rect 67725 247754 67791 247757
rect 70166 247754 70226 248268
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 121453 248235 121519 248238
rect 122782 248236 122788 248300
rect 122852 248298 122858 248300
rect 124029 248298 124095 248301
rect 122852 248296 124095 248298
rect 122852 248240 124034 248296
rect 124090 248240 124095 248296
rect 122852 248238 124095 248240
rect 122852 248236 122858 248238
rect 124029 248235 124095 248238
rect 67725 247752 70226 247754
rect 67725 247696 67730 247752
rect 67786 247696 70226 247752
rect 67725 247694 70226 247696
rect 67725 247691 67791 247694
rect 120073 247618 120139 247621
rect 121637 247618 121703 247621
rect 119876 247616 121703 247618
rect 67633 247210 67699 247213
rect 70166 247210 70226 247588
rect 119876 247560 120078 247616
rect 120134 247560 121642 247616
rect 121698 247560 121703 247616
rect 119876 247558 121703 247560
rect 120073 247555 120139 247558
rect 121637 247555 121703 247558
rect 67633 247208 70226 247210
rect 67633 247152 67638 247208
rect 67694 247152 70226 247208
rect 67633 247150 70226 247152
rect 67633 247147 67699 247150
rect 121545 246938 121611 246941
rect 119876 246936 121611 246938
rect 67725 246394 67791 246397
rect 70166 246394 70226 246908
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 121545 246875 121611 246878
rect 67725 246392 70226 246394
rect 67725 246336 67730 246392
rect 67786 246336 70226 246392
rect 67725 246334 70226 246336
rect 67725 246331 67791 246334
rect 121453 246258 121519 246261
rect 119876 246256 121519 246258
rect 67633 245850 67699 245853
rect 70166 245850 70226 246228
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 121453 246195 121519 246198
rect 67633 245848 70226 245850
rect 67633 245792 67638 245848
rect 67694 245792 70226 245848
rect 67633 245790 70226 245792
rect 67633 245787 67699 245790
rect 121637 245578 121703 245581
rect 119876 245576 121703 245578
rect 69197 245034 69263 245037
rect 70166 245034 70226 245548
rect 119876 245520 121642 245576
rect 121698 245520 121703 245576
rect 119876 245518 121703 245520
rect 121637 245515 121703 245518
rect 579981 245578 580047 245581
rect 583520 245578 584960 245668
rect 579981 245576 584960 245578
rect 579981 245520 579986 245576
rect 580042 245520 584960 245576
rect 579981 245518 584960 245520
rect 579981 245515 580047 245518
rect 583520 245428 584960 245518
rect 69197 245032 70226 245034
rect 69197 244976 69202 245032
rect 69258 244976 70226 245032
rect 69197 244974 70226 244976
rect 69197 244971 69263 244974
rect 121545 244898 121611 244901
rect 119876 244896 121611 244898
rect 67449 244354 67515 244357
rect 70166 244354 70226 244868
rect 119876 244840 121550 244896
rect 121606 244840 121611 244896
rect 119876 244838 121611 244840
rect 121545 244835 121611 244838
rect 67449 244352 70226 244354
rect 67449 244296 67454 244352
rect 67510 244296 70226 244352
rect 67449 244294 70226 244296
rect 67449 244291 67515 244294
rect 121453 244218 121519 244221
rect 119876 244216 121519 244218
rect 67541 243674 67607 243677
rect 70166 243674 70226 244188
rect 119876 244160 121458 244216
rect 121514 244160 121519 244216
rect 119876 244158 121519 244160
rect 121453 244155 121519 244158
rect 67541 243672 70226 243674
rect 67541 243616 67546 243672
rect 67602 243616 70226 243672
rect 67541 243614 70226 243616
rect 67541 243611 67607 243614
rect 121729 243538 121795 243541
rect 119876 243536 121795 243538
rect 67633 243130 67699 243133
rect 70166 243130 70226 243508
rect 119876 243480 121734 243536
rect 121790 243480 121795 243536
rect 119876 243478 121795 243480
rect 121729 243475 121795 243478
rect 67633 243128 70226 243130
rect 67633 243072 67638 243128
rect 67694 243072 70226 243128
rect 67633 243070 70226 243072
rect 67633 243067 67699 243070
rect 59310 242934 67650 242994
rect 55070 242796 55076 242860
rect 55140 242858 55146 242860
rect 58566 242858 58572 242860
rect 55140 242798 58572 242858
rect 55140 242796 55146 242798
rect 58566 242796 58572 242798
rect 58636 242858 58642 242860
rect 59310 242858 59370 242934
rect 58636 242798 59370 242858
rect 67590 242858 67650 242934
rect 69982 242934 70226 242994
rect 69982 242858 70042 242934
rect 67590 242798 70042 242858
rect 70166 242828 70226 242934
rect 121453 242858 121519 242861
rect 119876 242856 121519 242858
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 58636 242796 58642 242798
rect 121453 242795 121519 242798
rect 67633 241906 67699 241909
rect 70166 241906 70226 242148
rect 67633 241904 70226 241906
rect 67633 241848 67638 241904
rect 67694 241848 70226 241904
rect 67633 241846 70226 241848
rect 67633 241843 67699 241846
rect 119846 241634 119906 242148
rect 129774 241634 129780 241636
rect 119846 241574 129780 241634
rect 129774 241572 129780 241574
rect 129844 241572 129850 241636
rect 121361 241498 121427 241501
rect 119876 241496 121427 241498
rect 119876 241468 121366 241496
rect -960 241090 480 241180
rect 3141 241090 3207 241093
rect -960 241088 3207 241090
rect -960 241032 3146 241088
rect 3202 241032 3207 241088
rect -960 241030 3207 241032
rect -960 240940 480 241030
rect 3141 241027 3207 241030
rect 70166 240954 70226 241468
rect 119846 241440 121366 241468
rect 121422 241440 121427 241496
rect 119846 241438 121427 241440
rect 119286 241164 119292 241228
rect 119356 241226 119362 241228
rect 119846 241226 119906 241438
rect 121361 241435 121427 241438
rect 119356 241166 119906 241226
rect 119356 241164 119362 241166
rect 64830 240894 70226 240954
rect 53598 240212 53604 240276
rect 53668 240274 53674 240276
rect 64830 240274 64890 240894
rect 121453 240818 121519 240821
rect 119876 240816 121519 240818
rect 70534 240276 70594 240788
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 121453 240755 121519 240758
rect 53668 240214 64890 240274
rect 53668 240212 53674 240214
rect 70526 240212 70532 240276
rect 70596 240212 70602 240276
rect 121453 240138 121519 240141
rect 119876 240136 121519 240138
rect 119876 240080 121458 240136
rect 121514 240080 121519 240136
rect 119876 240078 121519 240080
rect 121453 240075 121519 240078
rect 68645 239458 68711 239461
rect 321502 239458 321508 239460
rect 68645 239456 321508 239458
rect 68645 239400 68650 239456
rect 68706 239400 321508 239456
rect 68645 239398 321508 239400
rect 68645 239395 68711 239398
rect 321502 239396 321508 239398
rect 321572 239396 321578 239460
rect 59118 238580 59124 238644
rect 59188 238642 59194 238644
rect 72601 238642 72667 238645
rect 59188 238640 72667 238642
rect 59188 238584 72606 238640
rect 72662 238584 72667 238640
rect 59188 238582 72667 238584
rect 59188 238580 59194 238582
rect 72601 238579 72667 238582
rect 113817 238642 113883 238645
rect 128445 238642 128511 238645
rect 113817 238640 128511 238642
rect 113817 238584 113822 238640
rect 113878 238584 128450 238640
rect 128506 238584 128511 238640
rect 113817 238582 128511 238584
rect 113817 238579 113883 238582
rect 128445 238579 128511 238582
rect 117037 238506 117103 238509
rect 127617 238506 127683 238509
rect 117037 238504 127683 238506
rect 117037 238448 117042 238504
rect 117098 238448 127622 238504
rect 127678 238448 127683 238504
rect 117037 238446 127683 238448
rect 117037 238443 117103 238446
rect 127617 238443 127683 238446
rect 70526 237900 70532 237964
rect 70596 237962 70602 237964
rect 90357 237962 90423 237965
rect 70596 237960 90423 237962
rect 70596 237904 90362 237960
rect 90418 237904 90423 237960
rect 70596 237902 90423 237904
rect 70596 237900 70602 237902
rect 90357 237899 90423 237902
rect 60549 236602 60615 236605
rect 334198 236602 334204 236604
rect 60549 236600 334204 236602
rect 60549 236544 60554 236600
rect 60610 236544 334204 236600
rect 60549 236542 334204 236544
rect 60549 236539 60615 236542
rect 334198 236540 334204 236542
rect 334268 236540 334274 236604
rect 57094 235860 57100 235924
rect 57164 235922 57170 235924
rect 119337 235922 119403 235925
rect 57164 235920 119403 235922
rect 57164 235864 119342 235920
rect 119398 235864 119403 235920
rect 57164 235862 119403 235864
rect 57164 235860 57170 235862
rect 119337 235859 119403 235862
rect 68921 232658 68987 232661
rect 173198 232658 173204 232660
rect 68921 232656 173204 232658
rect 68921 232600 68926 232656
rect 68982 232600 173204 232656
rect 68921 232598 173204 232600
rect 68921 232595 68987 232598
rect 173198 232596 173204 232598
rect 173268 232596 173274 232660
rect 69054 232460 69060 232524
rect 69124 232522 69130 232524
rect 455413 232522 455479 232525
rect 69124 232520 455479 232522
rect 69124 232464 455418 232520
rect 455474 232464 455479 232520
rect 69124 232462 455479 232464
rect 69124 232460 69130 232462
rect 455413 232459 455479 232462
rect 580257 232386 580323 232389
rect 583520 232386 584960 232476
rect 580257 232384 584960 232386
rect 580257 232328 580262 232384
rect 580318 232328 584960 232384
rect 580257 232326 584960 232328
rect 580257 232323 580323 232326
rect 583520 232236 584960 232326
rect 80145 229802 80211 229805
rect 320214 229802 320220 229804
rect 80145 229800 320220 229802
rect 80145 229744 80150 229800
rect 80206 229744 320220 229800
rect 80145 229742 320220 229744
rect 80145 229739 80211 229742
rect 320214 229740 320220 229742
rect 320284 229740 320290 229804
rect -960 227884 480 228124
rect 114645 226266 114711 226269
rect 136633 226266 136699 226269
rect 114645 226264 136699 226266
rect 114645 226208 114650 226264
rect 114706 226208 136638 226264
rect 136694 226208 136699 226264
rect 114645 226206 136699 226208
rect 114645 226203 114711 226206
rect 136633 226203 136699 226206
rect 136633 225722 136699 225725
rect 338614 225722 338620 225724
rect 136633 225720 338620 225722
rect 136633 225664 136638 225720
rect 136694 225664 338620 225720
rect 136633 225662 338620 225664
rect 136633 225659 136699 225662
rect 338614 225660 338620 225662
rect 338684 225660 338690 225724
rect 69238 225524 69244 225588
rect 69308 225586 69314 225588
rect 462313 225586 462379 225589
rect 69308 225584 462379 225586
rect 69308 225528 462318 225584
rect 462374 225528 462379 225584
rect 69308 225526 462379 225528
rect 69308 225524 69314 225526
rect 462313 225523 462379 225526
rect 84285 220146 84351 220149
rect 328494 220146 328500 220148
rect 84285 220144 328500 220146
rect 84285 220088 84290 220144
rect 84346 220088 328500 220144
rect 84285 220086 328500 220088
rect 84285 220083 84351 220086
rect 328494 220084 328500 220086
rect 328564 220084 328570 220148
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3233 201922 3299 201925
rect -960 201920 3299 201922
rect -960 201864 3238 201920
rect 3294 201864 3299 201920
rect -960 201862 3299 201864
rect -960 201772 480 201862
rect 3233 201859 3299 201862
rect 106917 197978 106983 197981
rect 494094 197978 494100 197980
rect 106917 197976 494100 197978
rect 106917 197920 106922 197976
rect 106978 197920 494100 197976
rect 106917 197918 494100 197920
rect 106917 197915 106983 197918
rect 494094 197916 494100 197918
rect 494164 197916 494170 197980
rect 147029 193898 147095 193901
rect 263726 193898 263732 193900
rect 147029 193896 263732 193898
rect 147029 193840 147034 193896
rect 147090 193840 263732 193896
rect 147029 193838 263732 193840
rect 147029 193835 147095 193838
rect 263726 193836 263732 193838
rect 263796 193836 263802 193900
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 58566 188260 58572 188324
rect 58636 188322 58642 188324
rect 503805 188322 503871 188325
rect 58636 188320 503871 188322
rect 58636 188264 503810 188320
rect 503866 188264 503871 188320
rect 58636 188262 503871 188264
rect 58636 188260 58642 188262
rect 503805 188259 503871 188262
rect 304257 184242 304323 184245
rect 339534 184242 339540 184244
rect 304257 184240 339540 184242
rect 304257 184184 304262 184240
rect 304318 184184 339540 184240
rect 304257 184182 339540 184184
rect 304257 184179 304323 184182
rect 339534 184180 339540 184182
rect 339604 184180 339610 184244
rect 1301 181386 1367 181389
rect 118734 181386 118740 181388
rect 1301 181384 118740 181386
rect 1301 181328 1306 181384
rect 1362 181328 118740 181384
rect 1301 181326 118740 181328
rect 1301 181323 1367 181326
rect 118734 181324 118740 181326
rect 118804 181324 118810 181388
rect 242157 181386 242223 181389
rect 260046 181386 260052 181388
rect 242157 181384 260052 181386
rect 242157 181328 242162 181384
rect 242218 181328 260052 181384
rect 242157 181326 260052 181328
rect 242157 181323 242223 181326
rect 260046 181324 260052 181326
rect 260116 181324 260122 181388
rect 220077 180162 220143 180165
rect 258390 180162 258396 180164
rect 220077 180160 258396 180162
rect 220077 180104 220082 180160
rect 220138 180104 258396 180160
rect 220077 180102 258396 180104
rect 220077 180099 220143 180102
rect 258390 180100 258396 180102
rect 258460 180100 258466 180164
rect 224217 180026 224283 180029
rect 266302 180026 266308 180028
rect 224217 180024 266308 180026
rect 224217 179968 224222 180024
rect 224278 179968 266308 180024
rect 224217 179966 266308 179968
rect 224217 179963 224283 179966
rect 266302 179964 266308 179966
rect 266372 179964 266378 180028
rect 121453 179482 121519 179485
rect 214414 179482 214420 179484
rect 121453 179480 214420 179482
rect 121453 179424 121458 179480
rect 121514 179424 214420 179480
rect 121453 179422 214420 179424
rect 121453 179419 121519 179422
rect 214414 179420 214420 179422
rect 214484 179420 214490 179484
rect 491293 179346 491359 179349
rect 491293 179344 493794 179346
rect 491293 179288 491298 179344
rect 491354 179288 493794 179344
rect 491293 179286 493794 179288
rect 491293 179283 491359 179286
rect 493734 178908 493794 179286
rect 580257 179210 580323 179213
rect 583520 179210 584960 179300
rect 580257 179208 584960 179210
rect 580257 179152 580262 179208
rect 580318 179152 584960 179208
rect 580257 179150 584960 179152
rect 580257 179147 580323 179150
rect 583520 179060 584960 179150
rect 247677 178666 247743 178669
rect 255446 178666 255452 178668
rect 247677 178664 255452 178666
rect 247677 178608 247682 178664
rect 247738 178608 255452 178664
rect 247677 178606 255452 178608
rect 247677 178603 247743 178606
rect 255446 178604 255452 178606
rect 255516 178604 255522 178668
rect 318057 178666 318123 178669
rect 326061 178666 326127 178669
rect 318057 178664 326127 178666
rect 318057 178608 318062 178664
rect 318118 178608 326066 178664
rect 326122 178608 326127 178664
rect 318057 178606 326127 178608
rect 318057 178603 318123 178606
rect 326061 178603 326127 178606
rect 416773 178666 416839 178669
rect 416773 178664 420164 178666
rect 416773 178608 416778 178664
rect 416834 178608 420164 178664
rect 416773 178606 420164 178608
rect 416773 178603 416839 178606
rect 166206 178122 166212 178124
rect 113130 178062 166212 178122
rect 112110 177924 112116 177988
rect 112180 177986 112186 177988
rect 113130 177986 113190 178062
rect 166206 178060 166212 178062
rect 166276 178060 166282 178124
rect 112180 177926 113190 177986
rect 112180 177924 112186 177926
rect 496997 177850 497063 177853
rect 494316 177848 497063 177850
rect 494316 177792 497002 177848
rect 497058 177792 497063 177848
rect 494316 177790 497063 177792
rect 496997 177787 497063 177790
rect 97073 177716 97139 177717
rect 97022 177714 97028 177716
rect 96982 177654 97028 177714
rect 97092 177712 97139 177716
rect 97134 177656 97139 177712
rect 97022 177652 97028 177654
rect 97092 177652 97139 177656
rect 100702 177652 100708 177716
rect 100772 177714 100778 177716
rect 102041 177714 102107 177717
rect 100772 177712 102107 177714
rect 100772 177656 102046 177712
rect 102102 177656 102107 177712
rect 100772 177654 102107 177656
rect 100772 177652 100778 177654
rect 97073 177651 97139 177652
rect 102041 177651 102107 177654
rect 105670 177652 105676 177716
rect 105740 177714 105746 177716
rect 106181 177714 106247 177717
rect 110689 177716 110755 177717
rect 114369 177716 114435 177717
rect 110638 177714 110644 177716
rect 105740 177712 106247 177714
rect 105740 177656 106186 177712
rect 106242 177656 106247 177712
rect 105740 177654 106247 177656
rect 110598 177654 110644 177714
rect 110708 177712 110755 177716
rect 114318 177714 114324 177716
rect 110750 177656 110755 177712
rect 105740 177652 105746 177654
rect 106181 177651 106247 177654
rect 110638 177652 110644 177654
rect 110708 177652 110755 177656
rect 114278 177654 114324 177714
rect 114388 177712 114435 177716
rect 114430 177656 114435 177712
rect 114318 177652 114324 177654
rect 114388 177652 114435 177656
rect 118366 177652 118372 177716
rect 118436 177714 118442 177716
rect 118509 177714 118575 177717
rect 118436 177712 118575 177714
rect 118436 177656 118514 177712
rect 118570 177656 118575 177712
rect 118436 177654 118575 177656
rect 118436 177652 118442 177654
rect 110689 177651 110755 177652
rect 114369 177651 114435 177652
rect 118509 177651 118575 177654
rect 120758 177652 120764 177716
rect 120828 177714 120834 177716
rect 121361 177714 121427 177717
rect 120828 177712 121427 177714
rect 120828 177656 121366 177712
rect 121422 177656 121427 177712
rect 120828 177654 121427 177656
rect 120828 177652 120834 177654
rect 121361 177651 121427 177654
rect 125726 177652 125732 177716
rect 125796 177714 125802 177716
rect 126881 177714 126947 177717
rect 130745 177716 130811 177717
rect 132401 177716 132467 177717
rect 130694 177714 130700 177716
rect 125796 177712 126947 177714
rect 125796 177656 126886 177712
rect 126942 177656 126947 177712
rect 125796 177654 126947 177656
rect 130654 177654 130700 177714
rect 130764 177712 130811 177716
rect 132350 177714 132356 177716
rect 130806 177656 130811 177712
rect 125796 177652 125802 177654
rect 126881 177651 126947 177654
rect 130694 177652 130700 177654
rect 130764 177652 130811 177656
rect 132310 177654 132356 177714
rect 132420 177712 132467 177716
rect 132462 177656 132467 177712
rect 132350 177652 132356 177654
rect 132420 177652 132467 177656
rect 130745 177651 130811 177652
rect 132401 177651 132467 177652
rect 238017 177578 238083 177581
rect 249374 177578 249380 177580
rect 238017 177576 249380 177578
rect 238017 177520 238022 177576
rect 238078 177520 249380 177576
rect 238017 177518 249380 177520
rect 238017 177515 238083 177518
rect 249374 177516 249380 177518
rect 249444 177516 249450 177580
rect 228357 177442 228423 177445
rect 289169 177442 289235 177445
rect 228357 177440 289235 177442
rect 228357 177384 228362 177440
rect 228418 177384 289174 177440
rect 289230 177384 289235 177440
rect 228357 177382 289235 177384
rect 228357 177379 228423 177382
rect 289169 177379 289235 177382
rect 312629 177442 312695 177445
rect 331438 177442 331444 177444
rect 312629 177440 331444 177442
rect 312629 177384 312634 177440
rect 312690 177384 331444 177440
rect 312629 177382 331444 177384
rect 312629 177379 312695 177382
rect 331438 177380 331444 177382
rect 331508 177380 331514 177444
rect 162117 177306 162183 177309
rect 184289 177306 184355 177309
rect 162117 177304 184355 177306
rect 162117 177248 162122 177304
rect 162178 177248 184294 177304
rect 184350 177248 184355 177304
rect 162117 177246 184355 177248
rect 162117 177243 162183 177246
rect 184289 177243 184355 177246
rect 222837 177306 222903 177309
rect 417509 177306 417575 177309
rect 222837 177304 417575 177306
rect 222837 177248 222842 177304
rect 222898 177248 417514 177304
rect 417570 177248 417575 177304
rect 222837 177246 417575 177248
rect 222837 177243 222903 177246
rect 417509 177243 417575 177246
rect 123150 177108 123156 177172
rect 123220 177170 123226 177172
rect 124121 177170 124187 177173
rect 123220 177168 124187 177170
rect 123220 177112 124126 177168
rect 124182 177112 124187 177168
rect 123220 177110 124187 177112
rect 123220 177108 123226 177110
rect 124121 177107 124187 177110
rect 108113 177036 108179 177037
rect 108062 177034 108068 177036
rect 108022 176974 108068 177034
rect 108132 177032 108179 177036
rect 108174 176976 108179 177032
rect 108062 176972 108068 176974
rect 108132 176972 108179 176976
rect 113214 176972 113220 177036
rect 113284 177034 113290 177036
rect 114001 177034 114067 177037
rect 115841 177036 115907 177037
rect 115790 177034 115796 177036
rect 113284 177032 114067 177034
rect 113284 176976 114006 177032
rect 114062 176976 114067 177032
rect 113284 176974 114067 176976
rect 115750 176974 115796 177034
rect 115860 177032 115907 177036
rect 115902 176976 115907 177032
rect 113284 176972 113290 176974
rect 108113 176971 108179 176972
rect 114001 176971 114067 176974
rect 115790 176972 115796 176974
rect 115860 176972 115907 176976
rect 115841 176971 115907 176972
rect 416773 177034 416839 177037
rect 416773 177032 420164 177034
rect 416773 176976 416778 177032
rect 416834 176976 420164 177032
rect 416773 176974 420164 176976
rect 416773 176971 416839 176974
rect 101990 176836 101996 176900
rect 102060 176898 102066 176900
rect 168230 176898 168236 176900
rect 102060 176838 168236 176898
rect 102060 176836 102066 176838
rect 168230 176836 168236 176838
rect 168300 176836 168306 176900
rect 100661 176762 100727 176765
rect 103329 176762 103395 176765
rect 107009 176764 107075 176765
rect 106958 176762 106964 176764
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 103286 176760 103395 176762
rect 103286 176704 103334 176760
rect 103390 176704 103395 176760
rect 103286 176699 103395 176704
rect 106918 176702 106964 176762
rect 107028 176760 107075 176764
rect 107070 176704 107075 176760
rect 106958 176700 106964 176702
rect 107028 176700 107075 176704
rect 109534 176700 109540 176764
rect 109604 176762 109610 176764
rect 109953 176762 110019 176765
rect 119521 176764 119587 176765
rect 119470 176762 119476 176764
rect 109604 176760 110019 176762
rect 109604 176704 109958 176760
rect 110014 176704 110019 176760
rect 109604 176702 110019 176704
rect 119430 176702 119476 176762
rect 119540 176760 119587 176764
rect 119582 176704 119587 176760
rect 109604 176700 109610 176702
rect 107009 176699 107075 176700
rect 109953 176699 110019 176702
rect 119470 176700 119476 176702
rect 119540 176700 119587 176704
rect 121862 176700 121868 176764
rect 121932 176762 121938 176764
rect 122097 176762 122163 176765
rect 124489 176764 124555 176765
rect 124438 176762 124444 176764
rect 121932 176760 122163 176762
rect 121932 176704 122102 176760
rect 122158 176704 122163 176760
rect 121932 176702 122163 176704
rect 124398 176702 124444 176762
rect 124508 176760 124555 176764
rect 124550 176704 124555 176760
rect 121932 176700 121938 176702
rect 119521 176699 119587 176700
rect 122097 176699 122163 176702
rect 124438 176700 124444 176702
rect 124508 176700 124555 176704
rect 127014 176700 127020 176764
rect 127084 176762 127090 176764
rect 127893 176762 127959 176765
rect 133137 176764 133203 176765
rect 134425 176764 134491 176765
rect 136081 176764 136147 176765
rect 133086 176762 133092 176764
rect 127084 176760 127959 176762
rect 127084 176704 127898 176760
rect 127954 176704 127959 176760
rect 127084 176702 127959 176704
rect 133046 176702 133092 176762
rect 133156 176760 133203 176764
rect 134374 176762 134380 176764
rect 133198 176704 133203 176760
rect 127084 176700 127090 176702
rect 124489 176699 124555 176700
rect 127893 176699 127959 176702
rect 133086 176700 133092 176702
rect 133156 176700 133203 176704
rect 134334 176702 134380 176762
rect 134444 176760 134491 176764
rect 136030 176762 136036 176764
rect 134486 176704 134491 176760
rect 134374 176700 134380 176702
rect 134444 176700 134491 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 269614 176700 269620 176764
rect 269684 176762 269690 176764
rect 316033 176762 316099 176765
rect 496997 176762 497063 176765
rect 269684 176760 316099 176762
rect 269684 176704 316038 176760
rect 316094 176704 316099 176760
rect 269684 176702 316099 176704
rect 494316 176760 497063 176762
rect 494316 176704 497002 176760
rect 497058 176704 497063 176760
rect 494316 176702 497063 176704
rect 269684 176700 269690 176702
rect 133137 176699 133203 176700
rect 134425 176699 134491 176700
rect 136081 176699 136147 176700
rect 316033 176699 316099 176702
rect 496997 176699 497063 176702
rect 103286 176492 103346 176699
rect 246481 176626 246547 176629
rect 249742 176626 249748 176628
rect 246481 176624 249748 176626
rect 246481 176568 246486 176624
rect 246542 176568 249748 176624
rect 246481 176566 249748 176568
rect 246481 176563 246547 176566
rect 249742 176564 249748 176566
rect 249812 176564 249818 176628
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 213913 176218 213979 176221
rect 213913 176216 217242 176218
rect 213913 176160 213918 176216
rect 213974 176160 217242 176216
rect 213913 176158 217242 176160
rect 213913 176155 213979 176158
rect -960 175796 480 176036
rect 217182 175644 217242 176158
rect 228449 175946 228515 175949
rect 249190 175946 249196 175948
rect 228449 175944 249196 175946
rect 228449 175888 228454 175944
rect 228510 175888 249196 175944
rect 228449 175886 249196 175888
rect 228449 175883 228515 175886
rect 249190 175884 249196 175886
rect 249260 175884 249266 175948
rect 318241 175946 318307 175949
rect 335537 175946 335603 175949
rect 318241 175944 335603 175946
rect 318241 175888 318246 175944
rect 318302 175888 335542 175944
rect 335598 175888 335603 175944
rect 318241 175886 335603 175888
rect 318241 175883 318307 175886
rect 335537 175883 335603 175886
rect 304349 175810 304415 175813
rect 304349 175808 321386 175810
rect 304349 175752 304354 175808
rect 304410 175752 321386 175808
rect 304349 175750 321386 175752
rect 304349 175747 304415 175750
rect 249333 175674 249399 175677
rect 248860 175672 249399 175674
rect 248860 175616 249338 175672
rect 249394 175616 249399 175672
rect 248860 175614 249399 175616
rect 249333 175611 249399 175614
rect 296670 175614 310132 175674
rect 104617 175540 104683 175541
rect 116945 175540 117011 175541
rect 128169 175540 128235 175541
rect 129457 175540 129523 175541
rect 148225 175540 148291 175541
rect 158897 175540 158963 175541
rect 98310 175476 98316 175540
rect 98380 175538 98386 175540
rect 104566 175538 104572 175540
rect 98380 175478 103530 175538
rect 104526 175478 104572 175538
rect 104636 175536 104683 175540
rect 116894 175538 116900 175540
rect 104678 175480 104683 175536
rect 98380 175476 98386 175478
rect 103470 175402 103530 175478
rect 104566 175476 104572 175478
rect 104636 175476 104683 175480
rect 116854 175478 116900 175538
rect 116964 175536 117011 175540
rect 128118 175538 128124 175540
rect 117006 175480 117011 175536
rect 116894 175476 116900 175478
rect 116964 175476 117011 175480
rect 128078 175478 128124 175538
rect 128188 175536 128235 175540
rect 129406 175538 129412 175540
rect 128230 175480 128235 175536
rect 128118 175476 128124 175478
rect 128188 175476 128235 175480
rect 129366 175478 129412 175538
rect 129476 175536 129523 175540
rect 148174 175538 148180 175540
rect 129518 175480 129523 175536
rect 129406 175476 129412 175478
rect 129476 175476 129523 175480
rect 148134 175478 148180 175538
rect 148244 175536 148291 175540
rect 158846 175538 158852 175540
rect 148286 175480 148291 175536
rect 148174 175476 148180 175478
rect 148244 175476 148291 175480
rect 158806 175478 158852 175538
rect 158916 175536 158963 175540
rect 158958 175480 158963 175536
rect 158846 175476 158852 175478
rect 158916 175476 158963 175480
rect 104617 175475 104683 175476
rect 116945 175475 117011 175476
rect 128169 175475 128235 175476
rect 129457 175475 129523 175476
rect 148225 175475 148291 175476
rect 158897 175475 158963 175476
rect 213269 175402 213335 175405
rect 103470 175400 213335 175402
rect 103470 175344 213274 175400
rect 213330 175344 213335 175400
rect 103470 175342 213335 175344
rect 213269 175339 213335 175342
rect 262070 175340 262076 175404
rect 262140 175402 262146 175404
rect 296670 175402 296730 175614
rect 321326 175508 321386 175750
rect 498101 175674 498167 175677
rect 494316 175672 498167 175674
rect 494316 175616 498106 175672
rect 498162 175616 498167 175672
rect 494316 175614 498167 175616
rect 498101 175611 498167 175614
rect 262140 175342 296730 175402
rect 262140 175340 262146 175342
rect 249149 175266 249215 175269
rect 248952 175264 249215 175266
rect 248952 175208 249154 175264
rect 249210 175208 249215 175264
rect 248952 175206 249215 175208
rect 249149 175203 249215 175206
rect 307385 175266 307451 175269
rect 321461 175266 321527 175269
rect 416773 175266 416839 175269
rect 307385 175264 310040 175266
rect 307385 175208 307390 175264
rect 307446 175208 310040 175264
rect 307385 175206 310040 175208
rect 321461 175264 321570 175266
rect 321461 175208 321466 175264
rect 321522 175208 321570 175264
rect 307385 175203 307451 175206
rect 321461 175203 321570 175208
rect 416773 175264 420164 175266
rect 416773 175208 416778 175264
rect 416834 175208 420164 175264
rect 416773 175206 420164 175208
rect 416773 175203 416839 175206
rect 213913 175130 213979 175133
rect 213913 175128 217242 175130
rect 213913 175072 213918 175128
rect 213974 175072 217242 175128
rect 213913 175070 217242 175072
rect 213913 175067 213979 175070
rect 217182 174964 217242 175070
rect 307477 174858 307543 174861
rect 307477 174856 310040 174858
rect 307477 174800 307482 174856
rect 307538 174800 310040 174856
rect 307477 174798 310040 174800
rect 307477 174795 307543 174798
rect 214005 174722 214071 174725
rect 214005 174720 217242 174722
rect 214005 174664 214010 174720
rect 214066 174664 217242 174720
rect 249149 174706 249215 174709
rect 214005 174662 217242 174664
rect 214005 174659 214071 174662
rect 217182 174284 217242 174662
rect 248860 174704 249215 174706
rect 248860 174648 249154 174704
rect 249210 174648 249215 174704
rect 321510 174692 321570 175203
rect 248860 174646 249215 174648
rect 249149 174643 249215 174646
rect 335854 174524 335860 174588
rect 335924 174586 335930 174588
rect 348417 174586 348483 174589
rect 335924 174584 348483 174586
rect 335924 174528 348422 174584
rect 348478 174528 348483 174584
rect 335924 174526 348483 174528
rect 335924 174524 335930 174526
rect 348417 174523 348483 174526
rect 307661 174450 307727 174453
rect 496997 174450 497063 174453
rect 307661 174448 310040 174450
rect 307661 174392 307666 174448
rect 307722 174392 310040 174448
rect 307661 174390 310040 174392
rect 494316 174448 497063 174450
rect 494316 174392 497002 174448
rect 497058 174392 497063 174448
rect 494316 174390 497063 174392
rect 307661 174387 307727 174390
rect 496997 174387 497063 174390
rect 249190 174314 249196 174316
rect 248952 174254 249196 174314
rect 249190 174252 249196 174254
rect 249260 174252 249266 174316
rect 164877 174042 164943 174045
rect 165613 174042 165679 174045
rect 164877 174040 165679 174042
rect 164877 173984 164882 174040
rect 164938 173984 165618 174040
rect 165674 173984 165679 174040
rect 164877 173982 165679 173984
rect 164877 173979 164943 173982
rect 165613 173979 165679 173982
rect 305729 174042 305795 174045
rect 307385 174042 307451 174045
rect 305729 174040 307451 174042
rect 305729 173984 305734 174040
rect 305790 173984 307390 174040
rect 307446 173984 307451 174040
rect 305729 173982 307451 173984
rect 305729 173979 305795 173982
rect 307385 173979 307451 173982
rect 307569 174042 307635 174045
rect 324313 174042 324379 174045
rect 307569 174040 310040 174042
rect 307569 173984 307574 174040
rect 307630 173984 310040 174040
rect 307569 173982 310040 173984
rect 321908 174040 324379 174042
rect 321908 173984 324318 174040
rect 324374 173984 324379 174040
rect 321908 173982 324379 173984
rect 307569 173979 307635 173982
rect 324313 173979 324379 173982
rect 213913 173770 213979 173773
rect 249374 173770 249380 173772
rect 213913 173768 217242 173770
rect 213913 173712 213918 173768
rect 213974 173712 217242 173768
rect 213913 173710 217242 173712
rect 248952 173710 249380 173770
rect 213913 173707 213979 173710
rect 217182 173604 217242 173710
rect 249374 173708 249380 173710
rect 249444 173708 249450 173772
rect 307569 173634 307635 173637
rect 307569 173632 310040 173634
rect 307569 173576 307574 173632
rect 307630 173576 310040 173632
rect 307569 173574 310040 173576
rect 307569 173571 307635 173574
rect 214005 173362 214071 173365
rect 249241 173362 249307 173365
rect 214005 173360 217242 173362
rect 214005 173304 214010 173360
rect 214066 173304 217242 173360
rect 214005 173302 217242 173304
rect 248952 173360 249307 173362
rect 248952 173304 249246 173360
rect 249302 173304 249307 173360
rect 248952 173302 249307 173304
rect 214005 173299 214071 173302
rect 217182 172924 217242 173302
rect 249241 173299 249307 173302
rect 307477 173226 307543 173229
rect 324313 173226 324379 173229
rect 307477 173224 310040 173226
rect 307477 173168 307482 173224
rect 307538 173168 310040 173224
rect 307477 173166 310040 173168
rect 321908 173224 324379 173226
rect 321908 173168 324318 173224
rect 324374 173168 324379 173224
rect 321908 173166 324379 173168
rect 307477 173163 307543 173166
rect 324313 173163 324379 173166
rect 249425 172818 249491 172821
rect 248952 172816 249491 172818
rect 248952 172760 249430 172816
rect 249486 172760 249491 172816
rect 248952 172758 249491 172760
rect 249425 172755 249491 172758
rect 307661 172682 307727 172685
rect 321277 172682 321343 172685
rect 307661 172680 310040 172682
rect 307661 172624 307666 172680
rect 307722 172624 310040 172680
rect 307661 172622 310040 172624
rect 321277 172680 321386 172682
rect 321277 172624 321282 172680
rect 321338 172624 321386 172680
rect 307661 172619 307727 172622
rect 321277 172619 321386 172624
rect 214097 172410 214163 172413
rect 252461 172410 252527 172413
rect 214097 172408 217242 172410
rect 214097 172352 214102 172408
rect 214158 172352 217242 172408
rect 214097 172350 217242 172352
rect 248952 172408 252527 172410
rect 248952 172352 252466 172408
rect 252522 172352 252527 172408
rect 321326 172380 321386 172619
rect 336038 172484 336044 172548
rect 336108 172546 336114 172548
rect 420134 172546 420194 173604
rect 496854 173362 496860 173364
rect 494316 173302 496860 173362
rect 496854 173300 496860 173302
rect 496924 173300 496930 173364
rect 336108 172486 420194 172546
rect 336108 172484 336114 172486
rect 248952 172350 252527 172352
rect 214097 172347 214163 172350
rect 217182 172244 217242 172350
rect 252461 172347 252527 172350
rect 306557 172274 306623 172277
rect 306557 172272 310040 172274
rect 306557 172216 306562 172272
rect 306618 172216 310040 172272
rect 306557 172214 310040 172216
rect 306557 172211 306623 172214
rect 213913 172002 213979 172005
rect 213913 172000 217242 172002
rect 213913 171944 213918 172000
rect 213974 171944 217242 172000
rect 213913 171942 217242 171944
rect 213913 171939 213979 171942
rect 167637 171594 167703 171597
rect 164694 171592 167703 171594
rect 164694 171536 167642 171592
rect 167698 171536 167703 171592
rect 217182 171564 217242 171942
rect 252369 171866 252435 171869
rect 248952 171864 252435 171866
rect 248952 171808 252374 171864
rect 252430 171808 252435 171864
rect 248952 171806 252435 171808
rect 252369 171803 252435 171806
rect 307661 171866 307727 171869
rect 416773 171866 416839 171869
rect 307661 171864 310040 171866
rect 307661 171808 307666 171864
rect 307722 171808 310040 171864
rect 307661 171806 310040 171808
rect 416773 171864 420164 171866
rect 416773 171808 416778 171864
rect 416834 171808 420164 171864
rect 416773 171806 420164 171808
rect 307661 171803 307727 171806
rect 416773 171803 416839 171806
rect 494286 171730 494346 172244
rect 494421 171730 494487 171733
rect 494286 171728 494487 171730
rect 164694 171534 167703 171536
rect 167637 171531 167703 171534
rect 250069 171458 250135 171461
rect 248952 171456 250135 171458
rect 248952 171400 250074 171456
rect 250130 171400 250135 171456
rect 248952 171398 250135 171400
rect 250069 171395 250135 171398
rect 307293 171458 307359 171461
rect 307293 171456 310040 171458
rect 307293 171400 307298 171456
rect 307354 171400 310040 171456
rect 307293 171398 310040 171400
rect 307293 171395 307359 171398
rect 321878 171322 321938 171700
rect 494286 171672 494426 171728
rect 494482 171672 494487 171728
rect 494286 171670 494487 171672
rect 494421 171667 494487 171670
rect 326061 171322 326127 171325
rect 321878 171320 326127 171322
rect 321878 171264 326066 171320
rect 326122 171264 326127 171320
rect 321878 171262 326127 171264
rect 326061 171259 326127 171262
rect 216998 171126 217242 171186
rect 213913 171050 213979 171053
rect 216998 171050 217058 171126
rect 213913 171048 217058 171050
rect 213913 170992 213918 171048
rect 213974 170992 217058 171048
rect 217182 171020 217242 171126
rect 494102 171053 494162 171156
rect 307293 171050 307359 171053
rect 307293 171048 310040 171050
rect 213913 170990 217058 170992
rect 307293 170992 307298 171048
rect 307354 170992 310040 171048
rect 307293 170990 310040 170992
rect 494102 171048 494211 171053
rect 494102 170992 494150 171048
rect 494206 170992 494211 171048
rect 494102 170990 494211 170992
rect 213913 170987 213979 170990
rect 307293 170987 307359 170990
rect 494145 170987 494211 170990
rect 252461 170914 252527 170917
rect 324313 170914 324379 170917
rect 248952 170912 252527 170914
rect 248952 170856 252466 170912
rect 252522 170856 252527 170912
rect 248952 170854 252527 170856
rect 321908 170912 324379 170914
rect 321908 170856 324318 170912
rect 324374 170856 324379 170912
rect 321908 170854 324379 170856
rect 252461 170851 252527 170854
rect 324313 170851 324379 170854
rect 214741 170778 214807 170781
rect 214741 170776 217242 170778
rect 214741 170720 214746 170776
rect 214802 170720 217242 170776
rect 214741 170718 217242 170720
rect 214741 170715 214807 170718
rect 217182 170340 217242 170718
rect 307569 170642 307635 170645
rect 321829 170642 321895 170645
rect 307569 170640 310040 170642
rect 307569 170584 307574 170640
rect 307630 170584 310040 170640
rect 307569 170582 310040 170584
rect 321829 170640 321938 170642
rect 321829 170584 321834 170640
rect 321890 170584 321938 170640
rect 307569 170579 307635 170582
rect 321829 170579 321938 170584
rect 252369 170506 252435 170509
rect 248952 170504 252435 170506
rect 248952 170448 252374 170504
rect 252430 170448 252435 170504
rect 248952 170446 252435 170448
rect 252369 170443 252435 170446
rect 307109 170234 307175 170237
rect 307109 170232 310040 170234
rect 307109 170176 307114 170232
rect 307170 170176 310040 170232
rect 307109 170174 310040 170176
rect 307109 170171 307175 170174
rect 252461 170098 252527 170101
rect 248952 170096 252527 170098
rect 248952 170040 252466 170096
rect 252522 170040 252527 170096
rect 321878 170068 321938 170579
rect 416773 170234 416839 170237
rect 416773 170232 420164 170234
rect 416773 170176 416778 170232
rect 416834 170176 420164 170232
rect 416773 170174 420164 170176
rect 416773 170171 416839 170174
rect 248952 170038 252527 170040
rect 252461 170035 252527 170038
rect 496997 169962 497063 169965
rect 494316 169960 497063 169962
rect 494316 169904 497002 169960
rect 497058 169904 497063 169960
rect 494316 169902 497063 169904
rect 496997 169899 497063 169902
rect 307661 169826 307727 169829
rect 216998 169766 217242 169826
rect 213913 169690 213979 169693
rect 216998 169690 217058 169766
rect 213913 169688 217058 169690
rect 213913 169632 213918 169688
rect 213974 169632 217058 169688
rect 217182 169660 217242 169766
rect 307661 169824 310040 169826
rect 307661 169768 307666 169824
rect 307722 169768 310040 169824
rect 307661 169766 310040 169768
rect 307661 169763 307727 169766
rect 213913 169630 217058 169632
rect 213913 169627 213979 169630
rect 252829 169554 252895 169557
rect 248952 169552 252895 169554
rect 248952 169496 252834 169552
rect 252890 169496 252895 169552
rect 248952 169494 252895 169496
rect 252829 169491 252895 169494
rect 321318 169492 321324 169556
rect 321388 169492 321394 169556
rect 214005 169418 214071 169421
rect 214005 169416 217242 169418
rect 214005 169360 214010 169416
rect 214066 169360 217242 169416
rect 321326 169388 321386 169492
rect 214005 169358 217242 169360
rect 214005 169355 214071 169358
rect 217182 168980 217242 169358
rect 307477 169282 307543 169285
rect 307477 169280 310040 169282
rect 307477 169224 307482 169280
rect 307538 169224 310040 169280
rect 307477 169222 310040 169224
rect 307477 169219 307543 169222
rect 252461 169146 252527 169149
rect 248952 169144 252527 169146
rect 248952 169088 252466 169144
rect 252522 169088 252527 169144
rect 248952 169086 252527 169088
rect 252461 169083 252527 169086
rect 307661 168874 307727 168877
rect 495525 168874 495591 168877
rect 307661 168872 310040 168874
rect 307661 168816 307666 168872
rect 307722 168816 310040 168872
rect 307661 168814 310040 168816
rect 494316 168872 495591 168874
rect 494316 168816 495530 168872
rect 495586 168816 495591 168872
rect 494316 168814 495591 168816
rect 307661 168811 307727 168814
rect 495525 168811 495591 168814
rect 252369 168602 252435 168605
rect 324497 168602 324563 168605
rect 248952 168600 252435 168602
rect 248952 168544 252374 168600
rect 252430 168544 252435 168600
rect 248952 168542 252435 168544
rect 321908 168600 324563 168602
rect 321908 168544 324502 168600
rect 324558 168544 324563 168600
rect 321908 168542 324563 168544
rect 252369 168539 252435 168542
rect 324497 168539 324563 168542
rect 307569 168466 307635 168469
rect 307569 168464 310040 168466
rect 307569 168408 307574 168464
rect 307630 168408 310040 168464
rect 307569 168406 310040 168408
rect 307569 168403 307635 168406
rect 335854 168404 335860 168468
rect 335924 168466 335930 168468
rect 335924 168406 420164 168466
rect 335924 168404 335930 168406
rect 213913 168058 213979 168061
rect 217182 168058 217242 168300
rect 249793 168194 249859 168197
rect 248952 168192 249859 168194
rect 248952 168136 249798 168192
rect 249854 168136 249859 168192
rect 248952 168134 249859 168136
rect 249793 168131 249859 168134
rect 213913 168056 217242 168058
rect 213913 168000 213918 168056
rect 213974 168000 217242 168056
rect 213913 167998 217242 168000
rect 307477 168058 307543 168061
rect 307477 168056 310040 168058
rect 307477 168000 307482 168056
rect 307538 168000 310040 168056
rect 307477 167998 310040 168000
rect 213913 167995 213979 167998
rect 307477 167995 307543 167998
rect 214005 167922 214071 167925
rect 214005 167920 217242 167922
rect 214005 167864 214010 167920
rect 214066 167864 217242 167920
rect 214005 167862 217242 167864
rect 214005 167859 214071 167862
rect 217182 167620 217242 167862
rect 324405 167786 324471 167789
rect 496997 167786 497063 167789
rect 321908 167784 324471 167786
rect 321908 167728 324410 167784
rect 324466 167728 324471 167784
rect 321908 167726 324471 167728
rect 494316 167784 497063 167786
rect 494316 167728 497002 167784
rect 497058 167728 497063 167784
rect 494316 167726 497063 167728
rect 324405 167723 324471 167726
rect 496997 167723 497063 167726
rect 252369 167650 252435 167653
rect 248952 167648 252435 167650
rect 248952 167592 252374 167648
rect 252430 167592 252435 167648
rect 248952 167590 252435 167592
rect 252369 167587 252435 167590
rect 307661 167650 307727 167653
rect 307661 167648 310040 167650
rect 307661 167592 307666 167648
rect 307722 167592 310040 167648
rect 307661 167590 310040 167592
rect 307661 167587 307727 167590
rect 252461 167242 252527 167245
rect 248952 167240 252527 167242
rect 248952 167184 252466 167240
rect 252522 167184 252527 167240
rect 248952 167182 252527 167184
rect 252461 167179 252527 167182
rect 307569 167242 307635 167245
rect 307569 167240 310040 167242
rect 307569 167184 307574 167240
rect 307630 167184 310040 167240
rect 307569 167182 310040 167184
rect 307569 167179 307635 167182
rect 324313 167106 324379 167109
rect 321908 167104 324379 167106
rect 321908 167048 324318 167104
rect 324374 167048 324379 167104
rect 321908 167046 324379 167048
rect 324313 167043 324379 167046
rect 214649 166970 214715 166973
rect 216998 166970 217242 167010
rect 214649 166968 217242 166970
rect 214649 166912 214654 166968
rect 214710 166950 217242 166968
rect 214710 166912 217058 166950
rect 217182 166940 217242 166950
rect 214649 166910 217058 166912
rect 214649 166907 214715 166910
rect 306741 166834 306807 166837
rect 306741 166832 310040 166834
rect 306741 166776 306746 166832
rect 306802 166776 310040 166832
rect 306741 166774 310040 166776
rect 306741 166771 306807 166774
rect 213913 166698 213979 166701
rect 252461 166698 252527 166701
rect 213913 166696 217242 166698
rect 213913 166640 213918 166696
rect 213974 166640 217242 166696
rect 213913 166638 217242 166640
rect 248952 166696 252527 166698
rect 248952 166640 252466 166696
rect 252522 166640 252527 166696
rect 248952 166638 252527 166640
rect 213913 166635 213979 166638
rect 217182 166396 217242 166638
rect 252461 166635 252527 166638
rect 307477 166426 307543 166429
rect 307477 166424 310040 166426
rect 307477 166368 307482 166424
rect 307538 166368 310040 166424
rect 307477 166366 310040 166368
rect 307477 166363 307543 166366
rect 255446 166290 255452 166292
rect 248952 166230 255452 166290
rect 255446 166228 255452 166230
rect 255516 166228 255522 166292
rect 324313 166290 324379 166293
rect 321908 166288 324379 166290
rect 321908 166232 324318 166288
rect 324374 166232 324379 166288
rect 321908 166230 324379 166232
rect 324313 166227 324379 166230
rect 213361 166154 213427 166157
rect 213361 166152 217242 166154
rect 213361 166096 213366 166152
rect 213422 166096 217242 166152
rect 213361 166094 217242 166096
rect 213361 166091 213427 166094
rect 217182 165716 217242 166094
rect 307661 165882 307727 165885
rect 307661 165880 310040 165882
rect 307661 165824 307666 165880
rect 307722 165824 310040 165880
rect 307661 165822 310040 165824
rect 307661 165819 307727 165822
rect 252461 165746 252527 165749
rect 248952 165744 252527 165746
rect 248952 165688 252466 165744
rect 252522 165688 252527 165744
rect 248952 165686 252527 165688
rect 252461 165683 252527 165686
rect 338798 165684 338804 165748
rect 338868 165746 338874 165748
rect 420134 165746 420194 166804
rect 496997 166698 497063 166701
rect 494316 166696 497063 166698
rect 494316 166640 497002 166696
rect 497058 166640 497063 166696
rect 494316 166638 497063 166640
rect 496997 166635 497063 166638
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 338868 165686 420194 165746
rect 583520 165732 584960 165822
rect 338868 165684 338874 165686
rect 307385 165474 307451 165477
rect 324313 165474 324379 165477
rect 496997 165474 497063 165477
rect 307385 165472 310040 165474
rect 307385 165416 307390 165472
rect 307446 165416 310040 165472
rect 307385 165414 310040 165416
rect 321908 165472 324379 165474
rect 321908 165416 324318 165472
rect 324374 165416 324379 165472
rect 321908 165414 324379 165416
rect 494316 165472 497063 165474
rect 494316 165416 497002 165472
rect 497058 165416 497063 165472
rect 494316 165414 497063 165416
rect 307385 165411 307451 165414
rect 324313 165411 324379 165414
rect 496997 165411 497063 165414
rect 213913 165338 213979 165341
rect 252461 165338 252527 165341
rect 213913 165336 217242 165338
rect 213913 165280 213918 165336
rect 213974 165280 217242 165336
rect 213913 165278 217242 165280
rect 248952 165336 252527 165338
rect 248952 165280 252466 165336
rect 252522 165280 252527 165336
rect 248952 165278 252527 165280
rect 213913 165275 213979 165278
rect 217182 165036 217242 165278
rect 252461 165275 252527 165278
rect 307201 165066 307267 165069
rect 416773 165066 416839 165069
rect 307201 165064 310040 165066
rect 307201 165008 307206 165064
rect 307262 165008 310040 165064
rect 307201 165006 310040 165008
rect 416773 165064 420164 165066
rect 416773 165008 416778 165064
rect 416834 165008 420164 165064
rect 416773 165006 420164 165008
rect 307201 165003 307267 165006
rect 416773 165003 416839 165006
rect 214005 164794 214071 164797
rect 252277 164794 252343 164797
rect 324405 164794 324471 164797
rect 214005 164792 217242 164794
rect 214005 164736 214010 164792
rect 214066 164736 217242 164792
rect 214005 164734 217242 164736
rect 248952 164792 252343 164794
rect 248952 164736 252282 164792
rect 252338 164736 252343 164792
rect 248952 164734 252343 164736
rect 321908 164792 324471 164794
rect 321908 164736 324410 164792
rect 324466 164736 324471 164792
rect 321908 164734 324471 164736
rect 214005 164731 214071 164734
rect 217182 164356 217242 164734
rect 252277 164731 252343 164734
rect 324405 164731 324471 164734
rect 307569 164658 307635 164661
rect 307569 164656 310040 164658
rect 307569 164600 307574 164656
rect 307630 164600 310040 164656
rect 307569 164598 310040 164600
rect 307569 164595 307635 164598
rect 252369 164386 252435 164389
rect 497089 164386 497155 164389
rect 248952 164384 252435 164386
rect 248952 164328 252374 164384
rect 252430 164328 252435 164384
rect 248952 164326 252435 164328
rect 494316 164384 497155 164386
rect 494316 164328 497094 164384
rect 497150 164328 497155 164384
rect 494316 164326 497155 164328
rect 252369 164323 252435 164326
rect 497089 164323 497155 164326
rect 307661 164250 307727 164253
rect 307661 164248 310040 164250
rect 307661 164192 307666 164248
rect 307722 164192 310040 164248
rect 307661 164190 310040 164192
rect 307661 164187 307727 164190
rect 213913 163978 213979 163981
rect 252461 163978 252527 163981
rect 324313 163978 324379 163981
rect 213913 163976 217242 163978
rect 213913 163920 213918 163976
rect 213974 163920 217242 163976
rect 213913 163918 217242 163920
rect 248952 163976 252527 163978
rect 248952 163920 252466 163976
rect 252522 163920 252527 163976
rect 248952 163918 252527 163920
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 213913 163915 213979 163918
rect 217182 163676 217242 163918
rect 252461 163915 252527 163918
rect 324313 163915 324379 163918
rect 307569 163842 307635 163845
rect 307569 163840 310040 163842
rect 307569 163784 307574 163840
rect 307630 163784 310040 163840
rect 307569 163782 310040 163784
rect 307569 163779 307635 163782
rect 252369 163434 252435 163437
rect 248952 163432 252435 163434
rect 248952 163376 252374 163432
rect 252430 163376 252435 163432
rect 248952 163374 252435 163376
rect 252369 163371 252435 163374
rect 307661 163434 307727 163437
rect 307661 163432 310040 163434
rect 307661 163376 307666 163432
rect 307722 163376 310040 163432
rect 307661 163374 310040 163376
rect 307661 163371 307727 163374
rect 324405 163162 324471 163165
rect 200070 163102 217242 163162
rect 321908 163160 324471 163162
rect 321908 163104 324410 163160
rect 324466 163104 324471 163160
rect 321908 163102 324471 163104
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 166206 162828 166212 162892
rect 166276 162890 166282 162892
rect 200070 162890 200130 163102
rect 217182 162996 217242 163102
rect 324405 163099 324471 163102
rect 252277 163026 252343 163029
rect 248952 163024 252343 163026
rect 248952 162968 252282 163024
rect 252338 162968 252343 163024
rect 248952 162966 252343 162968
rect 252277 162963 252343 162966
rect 307109 163026 307175 163029
rect 307109 163024 310040 163026
rect 307109 162968 307114 163024
rect 307170 162968 310040 163024
rect 307109 162966 310040 162968
rect 307109 162963 307175 162966
rect 166276 162830 200130 162890
rect 166276 162828 166282 162830
rect 345606 162828 345612 162892
rect 345676 162890 345682 162892
rect 420134 162890 420194 163404
rect 496997 163298 497063 163301
rect 494316 163296 497063 163298
rect 494316 163240 497002 163296
rect 497058 163240 497063 163296
rect 494316 163238 497063 163240
rect 496997 163235 497063 163238
rect 345676 162830 420194 162890
rect 345676 162828 345682 162830
rect 213913 162618 213979 162621
rect 213913 162616 217242 162618
rect 213913 162560 213918 162616
rect 213974 162560 217242 162616
rect 213913 162558 217242 162560
rect 213913 162555 213979 162558
rect 217182 162316 217242 162558
rect 252553 162482 252619 162485
rect 248952 162480 252619 162482
rect 248952 162424 252558 162480
rect 252614 162424 252619 162480
rect 248952 162422 252619 162424
rect 252553 162419 252619 162422
rect 307569 162482 307635 162485
rect 324313 162482 324379 162485
rect 307569 162480 310040 162482
rect 307569 162424 307574 162480
rect 307630 162424 310040 162480
rect 307569 162422 310040 162424
rect 321908 162480 324379 162482
rect 321908 162424 324318 162480
rect 324374 162424 324379 162480
rect 321908 162422 324379 162424
rect 307569 162419 307635 162422
rect 324313 162419 324379 162422
rect 496997 162210 497063 162213
rect 494316 162208 497063 162210
rect 494316 162152 497002 162208
rect 497058 162152 497063 162208
rect 494316 162150 497063 162152
rect 496997 162147 497063 162150
rect 214414 162012 214420 162076
rect 214484 162074 214490 162076
rect 252461 162074 252527 162077
rect 214484 162014 217242 162074
rect 248952 162072 252527 162074
rect 248952 162016 252466 162072
rect 252522 162016 252527 162072
rect 248952 162014 252527 162016
rect 214484 162012 214490 162014
rect 217182 161772 217242 162014
rect 252461 162011 252527 162014
rect 307661 162074 307727 162077
rect 307661 162072 310040 162074
rect 307661 162016 307666 162072
rect 307722 162016 310040 162072
rect 307661 162014 310040 162016
rect 307661 162011 307727 162014
rect 416773 161802 416839 161805
rect 416773 161800 420164 161802
rect 416773 161744 416778 161800
rect 416834 161744 420164 161800
rect 416773 161742 420164 161744
rect 416773 161739 416839 161742
rect 307293 161666 307359 161669
rect 324405 161666 324471 161669
rect 307293 161664 310040 161666
rect 307293 161608 307298 161664
rect 307354 161608 310040 161664
rect 307293 161606 310040 161608
rect 321908 161664 324471 161666
rect 321908 161608 324410 161664
rect 324466 161608 324471 161664
rect 321908 161606 324471 161608
rect 307293 161603 307359 161606
rect 324405 161603 324471 161606
rect 252369 161530 252435 161533
rect 248952 161528 252435 161530
rect 248952 161472 252374 161528
rect 252430 161472 252435 161528
rect 248952 161470 252435 161472
rect 252369 161467 252435 161470
rect 213913 161394 213979 161397
rect 213913 161392 217242 161394
rect 213913 161336 213918 161392
rect 213974 161336 217242 161392
rect 213913 161334 217242 161336
rect 213913 161331 213979 161334
rect 217182 161092 217242 161334
rect 307569 161258 307635 161261
rect 307569 161256 310040 161258
rect 307569 161200 307574 161256
rect 307630 161200 310040 161256
rect 307569 161198 310040 161200
rect 307569 161195 307635 161198
rect 248860 161018 249442 161078
rect 214557 160850 214623 160853
rect 249382 160850 249442 161018
rect 496997 160986 497063 160989
rect 494316 160984 497063 160986
rect 494316 160928 497002 160984
rect 497058 160928 497063 160984
rect 494316 160926 497063 160928
rect 496997 160923 497063 160926
rect 263726 160850 263732 160852
rect 214557 160848 217242 160850
rect 214557 160792 214562 160848
rect 214618 160792 217242 160848
rect 214557 160790 217242 160792
rect 249382 160790 263732 160850
rect 214557 160787 214623 160790
rect 168230 160652 168236 160716
rect 168300 160714 168306 160716
rect 214097 160714 214163 160717
rect 168300 160712 214163 160714
rect 168300 160656 214102 160712
rect 214158 160656 214163 160712
rect 168300 160654 214163 160656
rect 168300 160652 168306 160654
rect 214097 160651 214163 160654
rect 217182 160412 217242 160790
rect 263726 160788 263732 160790
rect 263796 160788 263802 160852
rect 307293 160850 307359 160853
rect 324313 160850 324379 160853
rect 307293 160848 310040 160850
rect 307293 160792 307298 160848
rect 307354 160792 310040 160848
rect 307293 160790 310040 160792
rect 321908 160848 324379 160850
rect 321908 160792 324318 160848
rect 324374 160792 324379 160848
rect 321908 160790 324379 160792
rect 307293 160787 307359 160790
rect 324313 160787 324379 160790
rect 249977 160578 250043 160581
rect 248952 160576 250043 160578
rect 248952 160520 249982 160576
rect 250038 160520 250043 160576
rect 248952 160518 250043 160520
rect 249977 160515 250043 160518
rect 307661 160442 307727 160445
rect 307661 160440 310040 160442
rect 307661 160384 307666 160440
rect 307722 160384 310040 160440
rect 307661 160382 310040 160384
rect 307661 160379 307727 160382
rect 252461 160306 252527 160309
rect 249198 160304 252527 160306
rect 249198 160248 252466 160304
rect 252522 160248 252527 160304
rect 249198 160246 252527 160248
rect 249198 160170 249258 160246
rect 252461 160243 252527 160246
rect 322933 160170 322999 160173
rect 248952 160110 249258 160170
rect 321908 160168 322999 160170
rect 321908 160112 322938 160168
rect 322994 160112 322999 160168
rect 321908 160110 322999 160112
rect 322933 160107 322999 160110
rect 307661 160034 307727 160037
rect 416773 160034 416839 160037
rect 307661 160032 310040 160034
rect 307661 159976 307666 160032
rect 307722 159976 310040 160032
rect 307661 159974 310040 159976
rect 416773 160032 420164 160034
rect 416773 159976 416778 160032
rect 416834 159976 420164 160032
rect 416773 159974 420164 159976
rect 307661 159971 307727 159974
rect 416773 159971 416839 159974
rect 213913 159898 213979 159901
rect 496997 159898 497063 159901
rect 213913 159896 217242 159898
rect 213913 159840 213918 159896
rect 213974 159840 217242 159896
rect 213913 159838 217242 159840
rect 494316 159896 497063 159898
rect 494316 159840 497002 159896
rect 497058 159840 497063 159896
rect 494316 159838 497063 159840
rect 213913 159835 213979 159838
rect 217182 159732 217242 159838
rect 496997 159835 497063 159838
rect 251725 159626 251791 159629
rect 248952 159624 251791 159626
rect 248952 159568 251730 159624
rect 251786 159568 251791 159624
rect 248952 159566 251791 159568
rect 251725 159563 251791 159566
rect 307109 159626 307175 159629
rect 307109 159624 310040 159626
rect 307109 159568 307114 159624
rect 307170 159568 310040 159624
rect 307109 159566 310040 159568
rect 307109 159563 307175 159566
rect 214005 159490 214071 159493
rect 214005 159488 217242 159490
rect 214005 159432 214010 159488
rect 214066 159432 217242 159488
rect 214005 159430 217242 159432
rect 214005 159427 214071 159430
rect 217182 159052 217242 159430
rect 324313 159354 324379 159357
rect 321908 159352 324379 159354
rect 321908 159296 324318 159352
rect 324374 159296 324379 159352
rect 321908 159294 324379 159296
rect 324313 159291 324379 159294
rect 252502 159218 252508 159220
rect 248952 159158 252508 159218
rect 252502 159156 252508 159158
rect 252572 159156 252578 159220
rect 306741 159082 306807 159085
rect 306741 159080 310040 159082
rect 306741 159024 306746 159080
rect 306802 159024 310040 159080
rect 306741 159022 310040 159024
rect 306741 159019 306807 159022
rect 252461 158810 252527 158813
rect 497089 158810 497155 158813
rect 248952 158808 252527 158810
rect 248952 158752 252466 158808
rect 252522 158752 252527 158808
rect 248952 158750 252527 158752
rect 494316 158808 497155 158810
rect 494316 158752 497094 158808
rect 497150 158752 497155 158808
rect 494316 158750 497155 158752
rect 252461 158747 252527 158750
rect 497089 158747 497155 158750
rect 213913 158674 213979 158677
rect 307569 158674 307635 158677
rect 213913 158672 217242 158674
rect 213913 158616 213918 158672
rect 213974 158616 217242 158672
rect 213913 158614 217242 158616
rect 213913 158611 213979 158614
rect 217182 158372 217242 158614
rect 307569 158672 310040 158674
rect 307569 158616 307574 158672
rect 307630 158616 310040 158672
rect 307569 158614 310040 158616
rect 307569 158611 307635 158614
rect 324313 158538 324379 158541
rect 321908 158536 324379 158538
rect 321908 158480 324318 158536
rect 324374 158480 324379 158536
rect 321908 158478 324379 158480
rect 324313 158475 324379 158478
rect 416773 158402 416839 158405
rect 416773 158400 420164 158402
rect 416773 158344 416778 158400
rect 416834 158344 420164 158400
rect 416773 158342 420164 158344
rect 416773 158339 416839 158342
rect 252461 158266 252527 158269
rect 248952 158264 252527 158266
rect 248952 158208 252466 158264
rect 252522 158208 252527 158264
rect 248952 158206 252527 158208
rect 252461 158203 252527 158206
rect 306557 158266 306623 158269
rect 306557 158264 310040 158266
rect 306557 158208 306562 158264
rect 306618 158208 310040 158264
rect 306557 158206 310040 158208
rect 306557 158203 306623 158206
rect 214097 158130 214163 158133
rect 214097 158128 217242 158130
rect 214097 158072 214102 158128
rect 214158 158072 217242 158128
rect 214097 158070 217242 158072
rect 214097 158067 214163 158070
rect 217182 157692 217242 158070
rect 251265 157858 251331 157861
rect 248952 157856 251331 157858
rect 248952 157800 251270 157856
rect 251326 157800 251331 157856
rect 248952 157798 251331 157800
rect 251265 157795 251331 157798
rect 307385 157858 307451 157861
rect 324405 157858 324471 157861
rect 307385 157856 310040 157858
rect 307385 157800 307390 157856
rect 307446 157800 310040 157856
rect 307385 157798 310040 157800
rect 321908 157856 324471 157858
rect 321908 157800 324410 157856
rect 324466 157800 324471 157856
rect 321908 157798 324471 157800
rect 307385 157795 307451 157798
rect 324405 157795 324471 157798
rect 496997 157722 497063 157725
rect 494316 157720 497063 157722
rect 494316 157664 497002 157720
rect 497058 157664 497063 157720
rect 494316 157662 497063 157664
rect 496997 157659 497063 157662
rect 307661 157450 307727 157453
rect 307661 157448 310040 157450
rect 307661 157392 307666 157448
rect 307722 157392 310040 157448
rect 307661 157390 310040 157392
rect 307661 157387 307727 157390
rect 213913 157314 213979 157317
rect 255262 157314 255268 157316
rect 213913 157312 217242 157314
rect 213913 157256 213918 157312
rect 213974 157256 217242 157312
rect 213913 157254 217242 157256
rect 248952 157254 255268 157314
rect 213913 157251 213979 157254
rect 217182 157148 217242 157254
rect 255262 157252 255268 157254
rect 255332 157252 255338 157316
rect 307477 157042 307543 157045
rect 324313 157042 324379 157045
rect 307477 157040 310040 157042
rect 307477 156984 307482 157040
rect 307538 156984 310040 157040
rect 307477 156982 310040 156984
rect 321908 157040 324379 157042
rect 321908 156984 324318 157040
rect 324374 156984 324379 157040
rect 321908 156982 324379 156984
rect 307477 156979 307543 156982
rect 324313 156979 324379 156982
rect 214005 156906 214071 156909
rect 252461 156906 252527 156909
rect 214005 156904 217242 156906
rect 214005 156848 214010 156904
rect 214066 156848 217242 156904
rect 214005 156846 217242 156848
rect 248952 156904 252527 156906
rect 248952 156848 252466 156904
rect 252522 156848 252527 156904
rect 248952 156846 252527 156848
rect 214005 156843 214071 156846
rect 217182 156468 217242 156846
rect 252461 156843 252527 156846
rect 307569 156634 307635 156637
rect 416773 156634 416839 156637
rect 307569 156632 310040 156634
rect 307569 156576 307574 156632
rect 307630 156576 310040 156632
rect 307569 156574 310040 156576
rect 416773 156632 420164 156634
rect 416773 156576 416778 156632
rect 416834 156576 420164 156632
rect 416773 156574 420164 156576
rect 307569 156571 307635 156574
rect 416773 156571 416839 156574
rect 496997 156498 497063 156501
rect 494316 156496 497063 156498
rect 494316 156440 497002 156496
rect 497058 156440 497063 156496
rect 494316 156438 497063 156440
rect 496997 156435 497063 156438
rect 251357 156362 251423 156365
rect 324313 156362 324379 156365
rect 248952 156360 251423 156362
rect 248952 156304 251362 156360
rect 251418 156304 251423 156360
rect 248952 156302 251423 156304
rect 321908 156360 324379 156362
rect 321908 156304 324318 156360
rect 324374 156304 324379 156360
rect 321908 156302 324379 156304
rect 251357 156299 251423 156302
rect 324313 156299 324379 156302
rect 307661 156226 307727 156229
rect 307661 156224 310040 156226
rect 307661 156168 307666 156224
rect 307722 156168 310040 156224
rect 307661 156166 310040 156168
rect 307661 156163 307727 156166
rect 213269 155954 213335 155957
rect 252645 155954 252711 155957
rect 213269 155952 217242 155954
rect 213269 155896 213274 155952
rect 213330 155896 217242 155952
rect 213269 155894 217242 155896
rect 248952 155952 252711 155954
rect 248952 155896 252650 155952
rect 252706 155896 252711 155952
rect 248952 155894 252711 155896
rect 213269 155891 213335 155894
rect 217182 155788 217242 155894
rect 252645 155891 252711 155894
rect 306557 155682 306623 155685
rect 306557 155680 310040 155682
rect 306557 155624 306562 155680
rect 306618 155624 310040 155680
rect 306557 155622 310040 155624
rect 306557 155619 306623 155622
rect 213913 155546 213979 155549
rect 324313 155546 324379 155549
rect 213913 155544 217242 155546
rect 213913 155488 213918 155544
rect 213974 155488 217242 155544
rect 213913 155486 217242 155488
rect 321908 155544 324379 155546
rect 321908 155488 324318 155544
rect 324374 155488 324379 155544
rect 321908 155486 324379 155488
rect 213913 155483 213979 155486
rect 217182 155108 217242 155486
rect 324313 155483 324379 155486
rect 252461 155410 252527 155413
rect 496997 155410 497063 155413
rect 248952 155408 252527 155410
rect 248952 155352 252466 155408
rect 252522 155352 252527 155408
rect 248952 155350 252527 155352
rect 494316 155408 497063 155410
rect 494316 155352 497002 155408
rect 497058 155352 497063 155408
rect 494316 155350 497063 155352
rect 252461 155347 252527 155350
rect 496997 155347 497063 155350
rect 307661 155274 307727 155277
rect 307661 155272 310040 155274
rect 307661 155216 307666 155272
rect 307722 155216 310040 155272
rect 307661 155214 310040 155216
rect 307661 155211 307727 155214
rect 252369 155002 252435 155005
rect 248952 155000 252435 155002
rect 248952 154944 252374 155000
rect 252430 154944 252435 155000
rect 248952 154942 252435 154944
rect 252369 154939 252435 154942
rect 416773 155002 416839 155005
rect 416773 155000 420164 155002
rect 416773 154944 416778 155000
rect 416834 154944 420164 155000
rect 416773 154942 420164 154944
rect 416773 154939 416839 154942
rect 307477 154866 307543 154869
rect 307477 154864 310040 154866
rect 307477 154808 307482 154864
rect 307538 154808 310040 154864
rect 307477 154806 310040 154808
rect 307477 154803 307543 154806
rect 324405 154730 324471 154733
rect 321908 154728 324471 154730
rect 321908 154672 324410 154728
rect 324466 154672 324471 154728
rect 321908 154670 324471 154672
rect 324405 154667 324471 154670
rect 249885 154458 249951 154461
rect 248952 154456 249951 154458
rect 214005 153914 214071 153917
rect 217182 153914 217242 154428
rect 248952 154400 249890 154456
rect 249946 154400 249951 154456
rect 248952 154398 249951 154400
rect 249885 154395 249951 154398
rect 306925 154458 306991 154461
rect 306925 154456 310040 154458
rect 306925 154400 306930 154456
rect 306986 154400 310040 154456
rect 306925 154398 310040 154400
rect 306925 154395 306991 154398
rect 496997 154322 497063 154325
rect 494316 154320 497063 154322
rect 494316 154264 497002 154320
rect 497058 154264 497063 154320
rect 494316 154262 497063 154264
rect 496997 154259 497063 154262
rect 252461 154050 252527 154053
rect 248952 154048 252527 154050
rect 248952 153992 252466 154048
rect 252522 153992 252527 154048
rect 248952 153990 252527 153992
rect 252461 153987 252527 153990
rect 306741 154050 306807 154053
rect 324313 154050 324379 154053
rect 306741 154048 310040 154050
rect 306741 153992 306746 154048
rect 306802 153992 310040 154048
rect 306741 153990 310040 153992
rect 321908 154048 324379 154050
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 306741 153987 306807 153990
rect 324313 153987 324379 153990
rect 214005 153912 217242 153914
rect 214005 153856 214010 153912
rect 214066 153856 217242 153912
rect 214005 153854 217242 153856
rect 214005 153851 214071 153854
rect 250805 153778 250871 153781
rect 258390 153778 258396 153780
rect 250805 153776 258396 153778
rect 213913 153370 213979 153373
rect 217182 153370 217242 153748
rect 250805 153720 250810 153776
rect 250866 153720 258396 153776
rect 250805 153718 258396 153720
rect 250805 153715 250871 153718
rect 258390 153716 258396 153718
rect 258460 153716 258466 153780
rect 307661 153642 307727 153645
rect 307661 153640 310040 153642
rect 307661 153584 307666 153640
rect 307722 153584 310040 153640
rect 307661 153582 310040 153584
rect 307661 153579 307727 153582
rect 252093 153506 252159 153509
rect 248952 153504 252159 153506
rect 248952 153448 252098 153504
rect 252154 153448 252159 153504
rect 248952 153446 252159 153448
rect 252093 153443 252159 153446
rect 213913 153368 217242 153370
rect 213913 153312 213918 153368
rect 213974 153312 217242 153368
rect 213913 153310 217242 153312
rect 213913 153307 213979 153310
rect 307661 153234 307727 153237
rect 324405 153234 324471 153237
rect 307661 153232 310040 153234
rect 307661 153176 307666 153232
rect 307722 153176 310040 153232
rect 307661 153174 310040 153176
rect 321908 153232 324471 153234
rect 321908 153176 324410 153232
rect 324466 153176 324471 153232
rect 321908 153174 324471 153176
rect 307661 153171 307727 153174
rect 324405 153171 324471 153174
rect 416773 153234 416839 153237
rect 497089 153234 497155 153237
rect 416773 153232 420164 153234
rect 416773 153176 416778 153232
rect 416834 153176 420164 153232
rect 416773 153174 420164 153176
rect 494316 153232 497155 153234
rect 494316 153176 497094 153232
rect 497150 153176 497155 153232
rect 494316 153174 497155 153176
rect 416773 153171 416839 153174
rect 497089 153171 497155 153174
rect 252277 153098 252343 153101
rect 248952 153096 252343 153098
rect 214005 152690 214071 152693
rect 217182 152690 217242 153068
rect 248952 153040 252282 153096
rect 252338 153040 252343 153096
rect 248952 153038 252343 153040
rect 252277 153035 252343 153038
rect 252461 152690 252527 152693
rect 214005 152688 217242 152690
rect 214005 152632 214010 152688
rect 214066 152632 217242 152688
rect 214005 152630 217242 152632
rect 248952 152688 252527 152690
rect 248952 152632 252466 152688
rect 252522 152632 252527 152688
rect 248952 152630 252527 152632
rect 214005 152627 214071 152630
rect 252461 152627 252527 152630
rect 307109 152690 307175 152693
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 307109 152688 310040 152690
rect 307109 152632 307114 152688
rect 307170 152632 310040 152688
rect 307109 152630 310040 152632
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 307109 152627 307175 152630
rect 579797 152627 579863 152630
rect 583520 152540 584960 152630
rect 213913 152010 213979 152013
rect 217182 152010 217242 152524
rect 324313 152418 324379 152421
rect 321908 152416 324379 152418
rect 321908 152360 324318 152416
rect 324374 152360 324379 152416
rect 321908 152358 324379 152360
rect 324313 152355 324379 152358
rect 306833 152282 306899 152285
rect 306833 152280 310040 152282
rect 306833 152224 306838 152280
rect 306894 152224 310040 152280
rect 306833 152222 310040 152224
rect 306833 152219 306899 152222
rect 252369 152146 252435 152149
rect 496997 152146 497063 152149
rect 248952 152144 252435 152146
rect 248952 152088 252374 152144
rect 252430 152088 252435 152144
rect 248952 152086 252435 152088
rect 494316 152144 497063 152146
rect 494316 152088 497002 152144
rect 497058 152088 497063 152144
rect 494316 152086 497063 152088
rect 252369 152083 252435 152086
rect 496997 152083 497063 152086
rect 213913 152008 217242 152010
rect 213913 151952 213918 152008
rect 213974 151952 217242 152008
rect 213913 151950 217242 151952
rect 213913 151947 213979 151950
rect 213453 151874 213519 151877
rect 306649 151874 306715 151877
rect 213453 151872 217058 151874
rect 213453 151816 213458 151872
rect 213514 151830 217058 151872
rect 306649 151872 310040 151874
rect 217182 151830 217242 151844
rect 213514 151816 217242 151830
rect 213453 151814 217242 151816
rect 213453 151811 213519 151814
rect 216998 151770 217242 151814
rect 306649 151816 306654 151872
rect 306710 151816 310040 151872
rect 306649 151814 310040 151816
rect 306649 151811 306715 151814
rect 252461 151738 252527 151741
rect 324313 151738 324379 151741
rect 248952 151736 252527 151738
rect 248952 151680 252466 151736
rect 252522 151680 252527 151736
rect 248952 151678 252527 151680
rect 321908 151736 324379 151738
rect 321908 151680 324318 151736
rect 324374 151680 324379 151736
rect 321908 151678 324379 151680
rect 252461 151675 252527 151678
rect 324313 151675 324379 151678
rect 416773 151602 416839 151605
rect 416773 151600 420164 151602
rect 416773 151544 416778 151600
rect 416834 151544 420164 151600
rect 416773 151542 420164 151544
rect 416773 151539 416839 151542
rect 307477 151466 307543 151469
rect 307477 151464 310040 151466
rect 307477 151408 307482 151464
rect 307538 151408 310040 151464
rect 307477 151406 310040 151408
rect 307477 151403 307543 151406
rect 252461 151194 252527 151197
rect 248952 151192 252527 151194
rect 215017 150786 215083 150789
rect 217182 150786 217242 151164
rect 248952 151136 252466 151192
rect 252522 151136 252527 151192
rect 248952 151134 252527 151136
rect 252461 151131 252527 151134
rect 307661 151058 307727 151061
rect 307661 151056 310040 151058
rect 307661 151000 307666 151056
rect 307722 151000 310040 151056
rect 307661 150998 310040 151000
rect 307661 150995 307727 150998
rect 324405 150922 324471 150925
rect 496997 150922 497063 150925
rect 321908 150920 324471 150922
rect 321908 150864 324410 150920
rect 324466 150864 324471 150920
rect 321908 150862 324471 150864
rect 494316 150920 497063 150922
rect 494316 150864 497002 150920
rect 497058 150864 497063 150920
rect 494316 150862 497063 150864
rect 324405 150859 324471 150862
rect 496997 150859 497063 150862
rect 252277 150786 252343 150789
rect 215017 150784 217242 150786
rect 215017 150728 215022 150784
rect 215078 150728 217242 150784
rect 215017 150726 217242 150728
rect 248952 150784 252343 150786
rect 248952 150728 252282 150784
rect 252338 150728 252343 150784
rect 248952 150726 252343 150728
rect 215017 150723 215083 150726
rect 252277 150723 252343 150726
rect 213913 150650 213979 150653
rect 307569 150650 307635 150653
rect 213913 150648 217242 150650
rect 213913 150592 213918 150648
rect 213974 150592 217242 150648
rect 213913 150590 217242 150592
rect 213913 150587 213979 150590
rect 217182 150484 217242 150590
rect 307569 150648 310040 150650
rect 307569 150592 307574 150648
rect 307630 150592 310040 150648
rect 307569 150590 310040 150592
rect 307569 150587 307635 150590
rect 252461 150242 252527 150245
rect 248952 150240 252527 150242
rect 248952 150184 252466 150240
rect 252522 150184 252527 150240
rect 248952 150182 252527 150184
rect 252461 150179 252527 150182
rect 307569 150242 307635 150245
rect 307569 150240 310040 150242
rect 307569 150184 307574 150240
rect 307630 150184 310040 150240
rect 307569 150182 310040 150184
rect 307569 150179 307635 150182
rect 213913 150106 213979 150109
rect 324313 150106 324379 150109
rect 213913 150104 217242 150106
rect 213913 150048 213918 150104
rect 213974 150048 217242 150104
rect 213913 150046 217242 150048
rect 321908 150104 324379 150106
rect 321908 150048 324318 150104
rect 324374 150048 324379 150104
rect 321908 150046 324379 150048
rect 213913 150043 213979 150046
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect 217182 149804 217242 150046
rect 324313 150043 324379 150046
rect 252277 149834 252343 149837
rect 248952 149832 252343 149834
rect -960 149774 3483 149776
rect 248952 149776 252282 149832
rect 252338 149776 252343 149832
rect 248952 149774 252343 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 252277 149771 252343 149774
rect 307150 149772 307156 149836
rect 307220 149834 307226 149836
rect 416773 149834 416839 149837
rect 496997 149834 497063 149837
rect 307220 149774 310040 149834
rect 416773 149832 420164 149834
rect 416773 149776 416778 149832
rect 416834 149776 420164 149832
rect 416773 149774 420164 149776
rect 494316 149832 497063 149834
rect 494316 149776 497002 149832
rect 497058 149776 497063 149832
rect 494316 149774 497063 149776
rect 307220 149772 307226 149774
rect 416773 149771 416839 149774
rect 496997 149771 497063 149774
rect 251766 149636 251772 149700
rect 251836 149698 251842 149700
rect 276749 149698 276815 149701
rect 251836 149696 276815 149698
rect 251836 149640 276754 149696
rect 276810 149640 276815 149696
rect 251836 149638 276815 149640
rect 251836 149636 251842 149638
rect 276749 149635 276815 149638
rect 214005 149562 214071 149565
rect 214005 149560 217242 149562
rect 214005 149504 214010 149560
rect 214066 149504 217242 149560
rect 214005 149502 217242 149504
rect 214005 149499 214071 149502
rect 217182 149124 217242 149502
rect 324313 149426 324379 149429
rect 321908 149424 324379 149426
rect 321908 149368 324318 149424
rect 324374 149368 324379 149424
rect 321908 149366 324379 149368
rect 324313 149363 324379 149366
rect 252369 149290 252435 149293
rect 248952 149288 252435 149290
rect 248952 149232 252374 149288
rect 252430 149232 252435 149288
rect 248952 149230 252435 149232
rect 252369 149227 252435 149230
rect 307661 149290 307727 149293
rect 307661 149288 310040 149290
rect 307661 149232 307666 149288
rect 307722 149232 310040 149288
rect 307661 149230 310040 149232
rect 307661 149227 307727 149230
rect 213913 148882 213979 148885
rect 252461 148882 252527 148885
rect 213913 148880 217242 148882
rect 213913 148824 213918 148880
rect 213974 148824 217242 148880
rect 213913 148822 217242 148824
rect 248952 148880 252527 148882
rect 248952 148824 252466 148880
rect 252522 148824 252527 148880
rect 248952 148822 252527 148824
rect 213913 148819 213979 148822
rect 217182 148444 217242 148822
rect 252461 148819 252527 148822
rect 307385 148882 307451 148885
rect 307385 148880 310040 148882
rect 307385 148824 307390 148880
rect 307446 148824 310040 148880
rect 307385 148822 310040 148824
rect 307385 148819 307451 148822
rect 496997 148746 497063 148749
rect 494316 148744 497063 148746
rect 494316 148688 497002 148744
rect 497058 148688 497063 148744
rect 494316 148686 497063 148688
rect 496997 148683 497063 148686
rect 324313 148610 324379 148613
rect 321908 148608 324379 148610
rect 321908 148552 324318 148608
rect 324374 148552 324379 148608
rect 321908 148550 324379 148552
rect 324313 148547 324379 148550
rect 307109 148474 307175 148477
rect 307109 148472 310040 148474
rect 307109 148416 307114 148472
rect 307170 148416 310040 148472
rect 307109 148414 310040 148416
rect 307109 148411 307175 148414
rect 252369 148338 252435 148341
rect 248952 148336 252435 148338
rect 248952 148280 252374 148336
rect 252430 148280 252435 148336
rect 248952 148278 252435 148280
rect 252369 148275 252435 148278
rect 416773 148202 416839 148205
rect 416773 148200 420164 148202
rect 416773 148144 416778 148200
rect 416834 148144 420164 148200
rect 416773 148142 420164 148144
rect 416773 148139 416839 148142
rect 213913 148066 213979 148069
rect 307017 148066 307083 148069
rect 213913 148064 217242 148066
rect 213913 148008 213918 148064
rect 213974 148008 217242 148064
rect 213913 148006 217242 148008
rect 213913 148003 213979 148006
rect 217182 147900 217242 148006
rect 307017 148064 310040 148066
rect 307017 148008 307022 148064
rect 307078 148008 310040 148064
rect 307017 148006 310040 148008
rect 307017 148003 307083 148006
rect 251173 147930 251239 147933
rect 248952 147928 251239 147930
rect 248952 147872 251178 147928
rect 251234 147872 251239 147928
rect 248952 147870 251239 147872
rect 251173 147867 251239 147870
rect 323209 147794 323275 147797
rect 321908 147792 323275 147794
rect 321908 147736 323214 147792
rect 323270 147736 323275 147792
rect 321908 147734 323275 147736
rect 323209 147731 323275 147734
rect 307477 147658 307543 147661
rect 495709 147658 495775 147661
rect 307477 147656 310040 147658
rect 307477 147600 307482 147656
rect 307538 147600 310040 147656
rect 307477 147598 310040 147600
rect 494316 147656 495775 147658
rect 494316 147600 495714 147656
rect 495770 147600 495775 147656
rect 494316 147598 495775 147600
rect 307477 147595 307543 147598
rect 495709 147595 495775 147598
rect 252461 147522 252527 147525
rect 248952 147520 252527 147522
rect 248952 147464 252466 147520
rect 252522 147464 252527 147520
rect 248952 147462 252527 147464
rect 252461 147459 252527 147462
rect 307569 147250 307635 147253
rect 307569 147248 310040 147250
rect 214005 146706 214071 146709
rect 217182 146706 217242 147220
rect 307569 147192 307574 147248
rect 307630 147192 310040 147248
rect 307569 147190 310040 147192
rect 307569 147187 307635 147190
rect 324313 147114 324379 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 324313 147051 324379 147054
rect 251449 146978 251515 146981
rect 248952 146976 251515 146978
rect 248952 146920 251454 146976
rect 251510 146920 251515 146976
rect 248952 146918 251515 146920
rect 251449 146915 251515 146918
rect 307661 146842 307727 146845
rect 307661 146840 310040 146842
rect 307661 146784 307666 146840
rect 307722 146784 310040 146840
rect 307661 146782 310040 146784
rect 307661 146779 307727 146782
rect 214005 146704 217242 146706
rect 214005 146648 214010 146704
rect 214066 146648 217242 146704
rect 214005 146646 217242 146648
rect 214005 146643 214071 146646
rect 252369 146570 252435 146573
rect 248952 146568 252435 146570
rect 213913 146434 213979 146437
rect 213913 146432 216874 146434
rect 213913 146376 213918 146432
rect 213974 146376 216874 146432
rect 213913 146374 216874 146376
rect 213913 146371 213979 146374
rect 216814 146298 216874 146374
rect 217366 146298 217426 146540
rect 248952 146512 252374 146568
rect 252430 146512 252435 146568
rect 248952 146510 252435 146512
rect 252369 146507 252435 146510
rect 416773 146570 416839 146573
rect 416773 146568 420164 146570
rect 416773 146512 416778 146568
rect 416834 146512 420164 146568
rect 416773 146510 420164 146512
rect 416773 146507 416839 146510
rect 307661 146434 307727 146437
rect 496997 146434 497063 146437
rect 307661 146432 310040 146434
rect 307661 146376 307666 146432
rect 307722 146376 310040 146432
rect 307661 146374 310040 146376
rect 494316 146432 497063 146434
rect 494316 146376 497002 146432
rect 497058 146376 497063 146432
rect 494316 146374 497063 146376
rect 307661 146371 307727 146374
rect 496997 146371 497063 146374
rect 324313 146298 324379 146301
rect 216814 146238 217426 146298
rect 321908 146296 324379 146298
rect 321908 146240 324318 146296
rect 324374 146240 324379 146296
rect 321908 146238 324379 146240
rect 324313 146235 324379 146238
rect 252461 146026 252527 146029
rect 248952 146024 252527 146026
rect 248952 145968 252466 146024
rect 252522 145968 252527 146024
rect 248952 145966 252527 145968
rect 252461 145963 252527 145966
rect 306557 145890 306623 145893
rect 306557 145888 310040 145890
rect 214649 145346 214715 145349
rect 217182 145346 217242 145860
rect 306557 145832 306562 145888
rect 306618 145832 310040 145888
rect 306557 145830 310040 145832
rect 306557 145827 306623 145830
rect 252369 145618 252435 145621
rect 248952 145616 252435 145618
rect 248952 145560 252374 145616
rect 252430 145560 252435 145616
rect 248952 145558 252435 145560
rect 252369 145555 252435 145558
rect 307293 145482 307359 145485
rect 324405 145482 324471 145485
rect 307293 145480 310040 145482
rect 307293 145424 307298 145480
rect 307354 145424 310040 145480
rect 307293 145422 310040 145424
rect 321908 145480 324471 145482
rect 321908 145424 324410 145480
rect 324466 145424 324471 145480
rect 321908 145422 324471 145424
rect 307293 145419 307359 145422
rect 324405 145419 324471 145422
rect 496997 145346 497063 145349
rect 214649 145344 217242 145346
rect 214649 145288 214654 145344
rect 214710 145288 217242 145344
rect 214649 145286 217242 145288
rect 494316 145344 497063 145346
rect 494316 145288 497002 145344
rect 497058 145288 497063 145344
rect 494316 145286 497063 145288
rect 214649 145283 214715 145286
rect 496997 145283 497063 145286
rect 168230 145012 168236 145076
rect 168300 145074 168306 145076
rect 168300 145014 200130 145074
rect 168300 145012 168306 145014
rect 200070 144938 200130 145014
rect 217366 144938 217426 145180
rect 251173 145074 251239 145077
rect 248952 145072 251239 145074
rect 248952 145016 251178 145072
rect 251234 145016 251239 145072
rect 248952 145014 251239 145016
rect 251173 145011 251239 145014
rect 306966 145012 306972 145076
rect 307036 145074 307042 145076
rect 307036 145014 310040 145074
rect 307036 145012 307042 145014
rect 200070 144878 217426 144938
rect 321502 144876 321508 144940
rect 321572 144876 321578 144940
rect 321510 144772 321570 144876
rect 416773 144802 416839 144805
rect 416773 144800 420164 144802
rect 416773 144744 416778 144800
rect 416834 144744 420164 144800
rect 416773 144742 420164 144744
rect 416773 144739 416839 144742
rect 250437 144666 250503 144669
rect 248952 144664 250503 144666
rect 248952 144608 250442 144664
rect 250498 144608 250503 144664
rect 248952 144606 250503 144608
rect 250437 144603 250503 144606
rect 306557 144666 306623 144669
rect 306557 144664 310040 144666
rect 306557 144608 306562 144664
rect 306618 144608 310040 144664
rect 306557 144606 310040 144608
rect 306557 144603 306623 144606
rect 214005 143986 214071 143989
rect 217182 143986 217242 144500
rect 307477 144258 307543 144261
rect 497089 144258 497155 144261
rect 307477 144256 310040 144258
rect 307477 144200 307482 144256
rect 307538 144200 310040 144256
rect 307477 144198 310040 144200
rect 494316 144256 497155 144258
rect 494316 144200 497094 144256
rect 497150 144200 497155 144256
rect 494316 144198 497155 144200
rect 307477 144195 307543 144198
rect 497089 144195 497155 144198
rect 250621 144122 250687 144125
rect 248952 144120 250687 144122
rect 248952 144064 250626 144120
rect 250682 144064 250687 144120
rect 248952 144062 250687 144064
rect 250621 144059 250687 144062
rect 324313 143986 324379 143989
rect 214005 143984 217242 143986
rect 214005 143928 214010 143984
rect 214066 143928 217242 143984
rect 214005 143926 217242 143928
rect 321908 143984 324379 143986
rect 321908 143928 324318 143984
rect 324374 143928 324379 143984
rect 321908 143926 324379 143928
rect 214005 143923 214071 143926
rect 324313 143923 324379 143926
rect 307661 143850 307727 143853
rect 307661 143848 310040 143850
rect 213913 143578 213979 143581
rect 217366 143578 217426 143820
rect 307661 143792 307666 143848
rect 307722 143792 310040 143848
rect 307661 143790 310040 143792
rect 307661 143787 307727 143790
rect 252461 143714 252527 143717
rect 248952 143712 252527 143714
rect 248952 143656 252466 143712
rect 252522 143656 252527 143712
rect 248952 143654 252527 143656
rect 252461 143651 252527 143654
rect 213913 143576 217426 143578
rect 213913 143520 213918 143576
rect 213974 143520 217426 143576
rect 213913 143518 217426 143520
rect 213913 143515 213979 143518
rect 307569 143442 307635 143445
rect 307569 143440 310040 143442
rect 307569 143384 307574 143440
rect 307630 143384 310040 143440
rect 307569 143382 310040 143384
rect 307569 143379 307635 143382
rect 213913 142762 213979 142765
rect 217182 142762 217242 143276
rect 252461 143170 252527 143173
rect 324313 143170 324379 143173
rect 248952 143168 252527 143170
rect 248952 143112 252466 143168
rect 252522 143112 252527 143168
rect 248952 143110 252527 143112
rect 321908 143168 324379 143170
rect 321908 143112 324318 143168
rect 324374 143112 324379 143168
rect 321908 143110 324379 143112
rect 252461 143107 252527 143110
rect 324313 143107 324379 143110
rect 416773 143170 416839 143173
rect 496997 143170 497063 143173
rect 416773 143168 420164 143170
rect 416773 143112 416778 143168
rect 416834 143112 420164 143168
rect 416773 143110 420164 143112
rect 494316 143168 497063 143170
rect 494316 143112 497002 143168
rect 497058 143112 497063 143168
rect 494316 143110 497063 143112
rect 416773 143107 416839 143110
rect 496997 143107 497063 143110
rect 306557 143034 306623 143037
rect 306557 143032 310040 143034
rect 306557 142976 306562 143032
rect 306618 142976 310040 143032
rect 306557 142974 310040 142976
rect 306557 142971 306623 142974
rect 252369 142762 252435 142765
rect 213913 142760 217242 142762
rect 213913 142704 213918 142760
rect 213974 142704 217242 142760
rect 213913 142702 217242 142704
rect 248952 142760 252435 142762
rect 248952 142704 252374 142760
rect 252430 142704 252435 142760
rect 248952 142702 252435 142704
rect 213913 142699 213979 142702
rect 252369 142699 252435 142702
rect 213269 142354 213335 142357
rect 217182 142354 217242 142596
rect 307661 142490 307727 142493
rect 325601 142490 325667 142493
rect 307661 142488 310040 142490
rect 307661 142432 307666 142488
rect 307722 142432 310040 142488
rect 307661 142430 310040 142432
rect 321908 142488 325667 142490
rect 321908 142432 325606 142488
rect 325662 142432 325667 142488
rect 321908 142430 325667 142432
rect 307661 142427 307727 142430
rect 325601 142427 325667 142430
rect 213269 142352 217242 142354
rect 213269 142296 213274 142352
rect 213330 142296 217242 142352
rect 213269 142294 217242 142296
rect 213269 142291 213335 142294
rect 266302 142218 266308 142220
rect 248952 142158 266308 142218
rect 266302 142156 266308 142158
rect 266372 142156 266378 142220
rect 306925 142082 306991 142085
rect 306925 142080 310040 142082
rect 306925 142024 306930 142080
rect 306986 142024 310040 142080
rect 306925 142022 310040 142024
rect 306925 142019 306991 142022
rect 321553 141946 321619 141949
rect 496997 141946 497063 141949
rect 321510 141944 321619 141946
rect 214005 141402 214071 141405
rect 217182 141402 217242 141916
rect 321510 141888 321558 141944
rect 321614 141888 321619 141944
rect 321510 141883 321619 141888
rect 494316 141944 497063 141946
rect 494316 141888 497002 141944
rect 497058 141888 497063 141944
rect 494316 141886 497063 141888
rect 496997 141883 497063 141886
rect 250805 141810 250871 141813
rect 248952 141808 250871 141810
rect 248952 141752 250810 141808
rect 250866 141752 250871 141808
rect 248952 141750 250871 141752
rect 250805 141747 250871 141750
rect 307017 141674 307083 141677
rect 307017 141672 310040 141674
rect 307017 141616 307022 141672
rect 307078 141616 310040 141672
rect 321510 141644 321570 141883
rect 307017 141614 310040 141616
rect 307017 141611 307083 141614
rect 252461 141402 252527 141405
rect 214005 141400 217242 141402
rect 214005 141344 214010 141400
rect 214066 141344 217242 141400
rect 214005 141342 217242 141344
rect 248952 141400 252527 141402
rect 248952 141344 252466 141400
rect 252522 141344 252527 141400
rect 248952 141342 252527 141344
rect 214005 141339 214071 141342
rect 252461 141339 252527 141342
rect 416773 141402 416839 141405
rect 416773 141400 420164 141402
rect 416773 141344 416778 141400
rect 416834 141344 420164 141400
rect 416773 141342 420164 141344
rect 416773 141339 416839 141342
rect 307569 141266 307635 141269
rect 307569 141264 310040 141266
rect 213913 140858 213979 140861
rect 217182 140858 217242 141236
rect 307569 141208 307574 141264
rect 307630 141208 310040 141264
rect 307569 141206 310040 141208
rect 307569 141203 307635 141206
rect 251173 140858 251239 140861
rect 213913 140856 217242 140858
rect 213913 140800 213918 140856
rect 213974 140800 217242 140856
rect 213913 140798 217242 140800
rect 248952 140856 251239 140858
rect 248952 140800 251178 140856
rect 251234 140800 251239 140856
rect 248952 140798 251239 140800
rect 213913 140795 213979 140798
rect 251173 140795 251239 140798
rect 307661 140858 307727 140861
rect 324313 140858 324379 140861
rect 496813 140858 496879 140861
rect 307661 140856 310040 140858
rect 307661 140800 307666 140856
rect 307722 140800 310040 140856
rect 307661 140798 310040 140800
rect 321908 140856 324379 140858
rect 321908 140800 324318 140856
rect 324374 140800 324379 140856
rect 321908 140798 324379 140800
rect 494316 140856 496879 140858
rect 494316 140800 496818 140856
rect 496874 140800 496879 140856
rect 494316 140798 496879 140800
rect 307661 140795 307727 140798
rect 324313 140795 324379 140798
rect 496813 140795 496879 140798
rect 214557 140042 214623 140045
rect 217182 140042 217242 140556
rect 252461 140450 252527 140453
rect 248952 140448 252527 140450
rect 248952 140392 252466 140448
rect 252522 140392 252527 140448
rect 248952 140390 252527 140392
rect 252461 140387 252527 140390
rect 306557 140450 306623 140453
rect 306557 140448 310040 140450
rect 306557 140392 306562 140448
rect 306618 140392 310040 140448
rect 306557 140390 310040 140392
rect 306557 140387 306623 140390
rect 324313 140178 324379 140181
rect 321908 140176 324379 140178
rect 321908 140120 324318 140176
rect 324374 140120 324379 140176
rect 321908 140118 324379 140120
rect 324313 140115 324379 140118
rect 214557 140040 217242 140042
rect 214557 139984 214562 140040
rect 214618 139984 217242 140040
rect 214557 139982 217242 139984
rect 258901 140042 258967 140045
rect 306966 140042 306972 140044
rect 258901 140040 306972 140042
rect 258901 139984 258906 140040
rect 258962 139984 306972 140040
rect 258901 139982 306972 139984
rect 214557 139979 214623 139982
rect 258901 139979 258967 139982
rect 306966 139980 306972 139982
rect 307036 139980 307042 140044
rect 309504 139938 310132 139998
rect 252369 139906 252435 139909
rect 248952 139904 252435 139906
rect 213913 139498 213979 139501
rect 217182 139498 217242 139876
rect 248952 139848 252374 139904
rect 252430 139848 252435 139904
rect 248952 139846 252435 139848
rect 252369 139843 252435 139846
rect 304206 139708 304212 139772
rect 304276 139770 304282 139772
rect 309504 139770 309564 139938
rect 304276 139710 309564 139770
rect 416773 139770 416839 139773
rect 496813 139770 496879 139773
rect 416773 139768 420164 139770
rect 416773 139712 416778 139768
rect 416834 139712 420164 139768
rect 416773 139710 420164 139712
rect 494316 139768 496879 139770
rect 494316 139712 496818 139768
rect 496874 139712 496879 139768
rect 494316 139710 496879 139712
rect 304276 139708 304282 139710
rect 416773 139707 416839 139710
rect 496813 139707 496879 139710
rect 307661 139634 307727 139637
rect 307661 139632 310040 139634
rect 307661 139576 307666 139632
rect 307722 139576 310040 139632
rect 307661 139574 310040 139576
rect 307661 139571 307727 139574
rect 252553 139498 252619 139501
rect 213913 139496 217242 139498
rect 213913 139440 213918 139496
rect 213974 139440 217242 139496
rect 213913 139438 217242 139440
rect 248952 139496 252619 139498
rect 248952 139440 252558 139496
rect 252614 139440 252619 139496
rect 248952 139438 252619 139440
rect 213913 139435 213979 139438
rect 252553 139435 252619 139438
rect 324313 139362 324379 139365
rect 321908 139360 324379 139362
rect 321908 139304 324318 139360
rect 324374 139304 324379 139360
rect 321908 139302 324379 139304
rect 324313 139299 324379 139302
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 214005 138818 214071 138821
rect 217182 138818 217242 139196
rect 306557 139090 306623 139093
rect 306557 139088 310040 139090
rect 306557 139032 306562 139088
rect 306618 139032 310040 139088
rect 306557 139030 310040 139032
rect 306557 139027 306623 139030
rect 252461 138954 252527 138957
rect 248952 138952 252527 138954
rect 248952 138896 252466 138952
rect 252522 138896 252527 138952
rect 248952 138894 252527 138896
rect 252461 138891 252527 138894
rect 214005 138816 217242 138818
rect 214005 138760 214010 138816
rect 214066 138760 217242 138816
rect 214005 138758 217242 138760
rect 214005 138755 214071 138758
rect 306925 138682 306991 138685
rect 496813 138682 496879 138685
rect 306925 138680 310040 138682
rect 213913 138138 213979 138141
rect 217182 138138 217242 138652
rect 306925 138624 306930 138680
rect 306986 138624 310040 138680
rect 306925 138622 310040 138624
rect 494316 138680 496879 138682
rect 494316 138624 496818 138680
rect 496874 138624 496879 138680
rect 494316 138622 496879 138624
rect 306925 138619 306991 138622
rect 496813 138619 496879 138622
rect 251817 138546 251883 138549
rect 324405 138546 324471 138549
rect 248952 138544 251883 138546
rect 248952 138488 251822 138544
rect 251878 138488 251883 138544
rect 248952 138486 251883 138488
rect 321908 138544 324471 138546
rect 321908 138488 324410 138544
rect 324466 138488 324471 138544
rect 321908 138486 324471 138488
rect 251817 138483 251883 138486
rect 324405 138483 324471 138486
rect 307661 138274 307727 138277
rect 307661 138272 310040 138274
rect 307661 138216 307666 138272
rect 307722 138216 310040 138272
rect 307661 138214 310040 138216
rect 307661 138211 307727 138214
rect 213913 138136 217242 138138
rect 213913 138080 213918 138136
rect 213974 138080 217242 138136
rect 213913 138078 217242 138080
rect 213913 138075 213979 138078
rect 252461 138002 252527 138005
rect 248952 138000 252527 138002
rect 213913 137458 213979 137461
rect 217182 137458 217242 137972
rect 248952 137944 252466 138000
rect 252522 137944 252527 138000
rect 248952 137942 252527 137944
rect 252461 137939 252527 137942
rect 416773 138002 416839 138005
rect 416773 138000 420164 138002
rect 416773 137944 416778 138000
rect 416834 137944 420164 138000
rect 416773 137942 420164 137944
rect 416773 137939 416839 137942
rect 307661 137866 307727 137869
rect 323025 137866 323091 137869
rect 307661 137864 310040 137866
rect 307661 137808 307666 137864
rect 307722 137808 310040 137864
rect 307661 137806 310040 137808
rect 321908 137864 323091 137866
rect 321908 137808 323030 137864
rect 323086 137808 323091 137864
rect 321908 137806 323091 137808
rect 307661 137803 307727 137806
rect 323025 137803 323091 137806
rect 256734 137594 256740 137596
rect 248952 137534 256740 137594
rect 256734 137532 256740 137534
rect 256804 137532 256810 137596
rect 213913 137456 217242 137458
rect 213913 137400 213918 137456
rect 213974 137400 217242 137456
rect 213913 137398 217242 137400
rect 307109 137458 307175 137461
rect 496813 137458 496879 137461
rect 307109 137456 310040 137458
rect 307109 137400 307114 137456
rect 307170 137400 310040 137456
rect 307109 137398 310040 137400
rect 494316 137456 496879 137458
rect 494316 137400 496818 137456
rect 496874 137400 496879 137456
rect 494316 137398 496879 137400
rect 213913 137395 213979 137398
rect 307109 137395 307175 137398
rect 496813 137395 496879 137398
rect 278313 137322 278379 137325
rect 307150 137322 307156 137324
rect 278313 137320 307156 137322
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 214005 136778 214071 136781
rect 217182 136778 217242 137292
rect 278313 137264 278318 137320
rect 278374 137264 307156 137320
rect 278313 137262 307156 137264
rect 278313 137259 278379 137262
rect 307150 137260 307156 137262
rect 307220 137260 307226 137324
rect 249742 137050 249748 137052
rect 248952 136990 249748 137050
rect 249742 136988 249748 136990
rect 249812 136988 249818 137052
rect 306966 136988 306972 137052
rect 307036 137050 307042 137052
rect 324313 137050 324379 137053
rect 307036 136990 310040 137050
rect 321908 137048 324379 137050
rect 321908 136992 324318 137048
rect 324374 136992 324379 137048
rect 321908 136990 324379 136992
rect 307036 136988 307042 136990
rect 324313 136987 324379 136990
rect 214005 136776 217242 136778
rect 214005 136720 214010 136776
rect 214066 136720 217242 136776
rect 214005 136718 217242 136720
rect 214005 136715 214071 136718
rect 250529 136642 250595 136645
rect 248952 136640 250595 136642
rect 214005 136098 214071 136101
rect 217182 136098 217242 136612
rect 248952 136584 250534 136640
rect 250590 136584 250595 136640
rect 248952 136582 250595 136584
rect 250529 136579 250595 136582
rect 307477 136642 307543 136645
rect 307477 136640 310040 136642
rect 307477 136584 307482 136640
rect 307538 136584 310040 136640
rect 307477 136582 310040 136584
rect 307477 136579 307543 136582
rect 324313 136370 324379 136373
rect 321908 136368 324379 136370
rect 321908 136312 324318 136368
rect 324374 136312 324379 136368
rect 321908 136310 324379 136312
rect 324313 136307 324379 136310
rect 416773 136370 416839 136373
rect 496813 136370 496879 136373
rect 416773 136368 420164 136370
rect 416773 136312 416778 136368
rect 416834 136312 420164 136368
rect 416773 136310 420164 136312
rect 494316 136368 496879 136370
rect 494316 136312 496818 136368
rect 496874 136312 496879 136368
rect 494316 136310 496879 136312
rect 416773 136307 416839 136310
rect 496813 136307 496879 136310
rect 252461 136234 252527 136237
rect 248952 136232 252527 136234
rect 248952 136176 252466 136232
rect 252522 136176 252527 136232
rect 248952 136174 252527 136176
rect 252461 136171 252527 136174
rect 306557 136234 306623 136237
rect 306557 136232 310040 136234
rect 306557 136176 306562 136232
rect 306618 136176 310040 136232
rect 306557 136174 310040 136176
rect 306557 136171 306623 136174
rect 325601 136098 325667 136101
rect 214005 136096 217242 136098
rect 214005 136040 214010 136096
rect 214066 136040 217242 136096
rect 214005 136038 217242 136040
rect 321878 136096 325667 136098
rect 321878 136040 325606 136096
rect 325662 136040 325667 136096
rect 321878 136038 325667 136040
rect 214005 136035 214071 136038
rect 214741 135554 214807 135557
rect 217182 135554 217242 135932
rect 252369 135690 252435 135693
rect 248952 135688 252435 135690
rect 248952 135632 252374 135688
rect 252430 135632 252435 135688
rect 248952 135630 252435 135632
rect 252369 135627 252435 135630
rect 307661 135690 307727 135693
rect 307661 135688 310040 135690
rect 307661 135632 307666 135688
rect 307722 135632 310040 135688
rect 307661 135630 310040 135632
rect 307661 135627 307727 135630
rect 214741 135552 217242 135554
rect 214741 135496 214746 135552
rect 214802 135496 217242 135552
rect 321878 135524 321938 136038
rect 325601 136035 325667 136038
rect 214741 135494 217242 135496
rect 214741 135491 214807 135494
rect 213913 135418 213979 135421
rect 213913 135416 217242 135418
rect 213913 135360 213918 135416
rect 213974 135360 217242 135416
rect 213913 135358 217242 135360
rect 213913 135355 213979 135358
rect 217182 135252 217242 135358
rect 252277 135282 252343 135285
rect 248952 135280 252343 135282
rect 248952 135224 252282 135280
rect 252338 135224 252343 135280
rect 248952 135222 252343 135224
rect 252277 135219 252343 135222
rect 307109 135282 307175 135285
rect 496997 135282 497063 135285
rect 307109 135280 310040 135282
rect 307109 135224 307114 135280
rect 307170 135224 310040 135280
rect 307109 135222 310040 135224
rect 494316 135280 497063 135282
rect 494316 135224 497002 135280
rect 497058 135224 497063 135280
rect 494316 135222 497063 135224
rect 307109 135219 307175 135222
rect 496997 135219 497063 135222
rect 307569 134874 307635 134877
rect 307569 134872 310040 134874
rect 307569 134816 307574 134872
rect 307630 134816 310040 134872
rect 307569 134814 310040 134816
rect 307569 134811 307635 134814
rect 252461 134738 252527 134741
rect 248952 134736 252527 134738
rect 248952 134680 252466 134736
rect 252522 134680 252527 134736
rect 248952 134678 252527 134680
rect 252461 134675 252527 134678
rect 170438 134132 170444 134196
rect 170508 134194 170514 134196
rect 217182 134194 217242 134572
rect 307661 134466 307727 134469
rect 307661 134464 310040 134466
rect 307661 134408 307666 134464
rect 307722 134408 310040 134464
rect 307661 134406 310040 134408
rect 307661 134403 307727 134406
rect 252369 134330 252435 134333
rect 248952 134328 252435 134330
rect 248952 134272 252374 134328
rect 252430 134272 252435 134328
rect 248952 134270 252435 134272
rect 252369 134267 252435 134270
rect 170508 134134 217242 134194
rect 321878 134194 321938 134708
rect 417325 134602 417391 134605
rect 419165 134602 419231 134605
rect 417325 134600 420164 134602
rect 417325 134544 417330 134600
rect 417386 134544 419170 134600
rect 419226 134544 420164 134600
rect 417325 134542 420164 134544
rect 417325 134539 417391 134542
rect 419165 134539 419231 134542
rect 330334 134194 330340 134196
rect 321878 134134 330340 134194
rect 170508 134132 170514 134134
rect 330334 134132 330340 134134
rect 330404 134132 330410 134196
rect 496813 134194 496879 134197
rect 494316 134192 496879 134194
rect 494316 134136 496818 134192
rect 496874 134136 496879 134192
rect 494316 134134 496879 134136
rect 496813 134131 496879 134134
rect 213913 134058 213979 134061
rect 307017 134058 307083 134061
rect 322974 134058 322980 134060
rect 213913 134056 217242 134058
rect 213913 134000 213918 134056
rect 213974 134000 217242 134056
rect 213913 133998 217242 134000
rect 213913 133995 213979 133998
rect 217182 133892 217242 133998
rect 307017 134056 310040 134058
rect 307017 134000 307022 134056
rect 307078 134000 310040 134056
rect 307017 133998 310040 134000
rect 321908 133998 322980 134058
rect 307017 133995 307083 133998
rect 322974 133996 322980 133998
rect 323044 133996 323050 134060
rect 252461 133786 252527 133789
rect 248952 133784 252527 133786
rect 248952 133728 252466 133784
rect 252522 133728 252527 133784
rect 248952 133726 252527 133728
rect 252461 133723 252527 133726
rect 306925 133650 306991 133653
rect 306925 133648 310040 133650
rect 306925 133592 306930 133648
rect 306986 133592 310040 133648
rect 306925 133590 310040 133592
rect 306925 133587 306991 133590
rect 252369 133378 252435 133381
rect 248952 133376 252435 133378
rect 166206 132772 166212 132836
rect 166276 132834 166282 132836
rect 217182 132834 217242 133348
rect 248952 133320 252374 133376
rect 252430 133320 252435 133376
rect 248952 133318 252435 133320
rect 252369 133315 252435 133318
rect 306557 133242 306623 133245
rect 324313 133242 324379 133245
rect 306557 133240 310040 133242
rect 306557 133184 306562 133240
rect 306618 133184 310040 133240
rect 306557 133182 310040 133184
rect 321908 133240 324379 133242
rect 321908 133184 324318 133240
rect 324374 133184 324379 133240
rect 321908 133182 324379 133184
rect 306557 133179 306623 133182
rect 324313 133179 324379 133182
rect 419349 132970 419415 132973
rect 495433 132970 495499 132973
rect 419349 132968 420164 132970
rect 419349 132912 419354 132968
rect 419410 132912 420164 132968
rect 419349 132910 420164 132912
rect 494316 132968 495499 132970
rect 494316 132912 495438 132968
rect 495494 132912 495499 132968
rect 494316 132910 495499 132912
rect 419349 132907 419415 132910
rect 495433 132907 495499 132910
rect 252277 132834 252343 132837
rect 166276 132774 217242 132834
rect 248952 132832 252343 132834
rect 248952 132776 252282 132832
rect 252338 132776 252343 132832
rect 248952 132774 252343 132776
rect 166276 132772 166282 132774
rect 252277 132771 252343 132774
rect 213913 132562 213979 132565
rect 213913 132560 216874 132562
rect 213913 132504 213918 132560
rect 213974 132510 216874 132560
rect 217366 132510 217426 132668
rect 302734 132636 302740 132700
rect 302804 132698 302810 132700
rect 302804 132638 310040 132698
rect 302804 132636 302810 132638
rect 213974 132504 217426 132510
rect 213913 132502 217426 132504
rect 213913 132499 213979 132502
rect 216814 132450 217426 132502
rect 252461 132426 252527 132429
rect 324313 132426 324379 132429
rect 248952 132424 252527 132426
rect 248952 132368 252466 132424
rect 252522 132368 252527 132424
rect 248952 132366 252527 132368
rect 321908 132424 324379 132426
rect 321908 132368 324318 132424
rect 324374 132368 324379 132424
rect 321908 132366 324379 132368
rect 252461 132363 252527 132366
rect 324313 132363 324379 132366
rect 307477 132290 307543 132293
rect 307477 132288 310040 132290
rect 307477 132232 307482 132288
rect 307538 132232 310040 132288
rect 307477 132230 310040 132232
rect 307477 132227 307543 132230
rect 494237 132154 494303 132157
rect 494237 132152 494346 132154
rect 494237 132096 494242 132152
rect 494298 132096 494346 132152
rect 494237 132091 494346 132096
rect 168966 131412 168972 131476
rect 169036 131474 169042 131476
rect 217182 131474 217242 131988
rect 252369 131882 252435 131885
rect 248952 131880 252435 131882
rect 248952 131824 252374 131880
rect 252430 131824 252435 131880
rect 248952 131822 252435 131824
rect 252369 131819 252435 131822
rect 307569 131882 307635 131885
rect 307569 131880 310040 131882
rect 307569 131824 307574 131880
rect 307630 131824 310040 131880
rect 494286 131852 494346 132091
rect 307569 131822 310040 131824
rect 307569 131819 307635 131822
rect 324405 131746 324471 131749
rect 321908 131744 324471 131746
rect 321908 131688 324410 131744
rect 324466 131688 324471 131744
rect 321908 131686 324471 131688
rect 324405 131683 324471 131686
rect 252093 131474 252159 131477
rect 169036 131414 217242 131474
rect 248952 131472 252159 131474
rect 248952 131416 252098 131472
rect 252154 131416 252159 131472
rect 248952 131414 252159 131416
rect 169036 131412 169042 131414
rect 252093 131411 252159 131414
rect 307661 131474 307727 131477
rect 307661 131472 310040 131474
rect 307661 131416 307666 131472
rect 307722 131416 310040 131472
rect 307661 131414 310040 131416
rect 307661 131411 307727 131414
rect 417601 131338 417667 131341
rect 419717 131338 419783 131341
rect 417601 131336 420164 131338
rect 213913 131202 213979 131205
rect 213913 131200 216874 131202
rect 213913 131144 213918 131200
rect 213974 131144 216874 131200
rect 213913 131142 216874 131144
rect 213913 131139 213979 131142
rect 216814 131066 216874 131142
rect 217366 131066 217426 131308
rect 417601 131280 417606 131336
rect 417662 131280 419722 131336
rect 419778 131280 420164 131336
rect 417601 131278 420164 131280
rect 417601 131275 417667 131278
rect 419717 131275 419783 131278
rect 216814 131006 217426 131066
rect 307477 131066 307543 131069
rect 494329 131066 494395 131069
rect 307477 131064 310040 131066
rect 307477 131008 307482 131064
rect 307538 131008 310040 131064
rect 307477 131006 310040 131008
rect 494286 131064 494395 131066
rect 494286 131008 494334 131064
rect 494390 131008 494395 131064
rect 307477 131003 307543 131006
rect 494286 131003 494395 131008
rect 252369 130930 252435 130933
rect 324313 130930 324379 130933
rect 248952 130928 252435 130930
rect 248952 130872 252374 130928
rect 252430 130872 252435 130928
rect 248952 130870 252435 130872
rect 321908 130928 324379 130930
rect 321908 130872 324318 130928
rect 324374 130872 324379 130928
rect 321908 130870 324379 130872
rect 252369 130867 252435 130870
rect 324313 130867 324379 130870
rect 494286 130764 494346 131003
rect 214649 130114 214715 130117
rect 217182 130114 217242 130628
rect 309550 130554 310132 130614
rect 252461 130522 252527 130525
rect 248952 130520 252527 130522
rect 248952 130464 252466 130520
rect 252522 130464 252527 130520
rect 248952 130462 252527 130464
rect 252461 130459 252527 130462
rect 252277 130114 252343 130117
rect 214649 130112 217242 130114
rect 214649 130056 214654 130112
rect 214710 130056 217242 130112
rect 214649 130054 217242 130056
rect 248952 130112 252343 130114
rect 248952 130056 252282 130112
rect 252338 130056 252343 130112
rect 248952 130054 252343 130056
rect 214649 130051 214715 130054
rect 252277 130051 252343 130054
rect 299974 130052 299980 130116
rect 300044 130114 300050 130116
rect 309550 130114 309610 130554
rect 300044 130054 309610 130114
rect 309734 130146 310132 130206
rect 300044 130052 300050 130054
rect 307569 129978 307635 129981
rect 309734 129978 309794 130146
rect 324405 130114 324471 130117
rect 321908 130112 324471 130114
rect 321908 130056 324410 130112
rect 324466 130056 324471 130112
rect 321908 130054 324471 130056
rect 324405 130051 324471 130054
rect 307569 129976 309794 129978
rect 213913 129842 213979 129845
rect 213913 129840 216874 129842
rect 213913 129784 213918 129840
rect 213974 129784 216874 129840
rect 213913 129782 216874 129784
rect 213913 129779 213979 129782
rect 216814 129706 216874 129782
rect 217366 129706 217426 129948
rect 307569 129920 307574 129976
rect 307630 129920 309794 129976
rect 307569 129918 309794 129920
rect 307569 129915 307635 129918
rect 307661 129842 307727 129845
rect 307661 129840 310040 129842
rect 307661 129784 307666 129840
rect 307722 129784 310040 129840
rect 307661 129782 310040 129784
rect 307661 129779 307727 129782
rect 496813 129706 496879 129709
rect 216814 129646 217426 129706
rect 494316 129704 496879 129706
rect 494316 129648 496818 129704
rect 496874 129648 496879 129704
rect 494316 129646 496879 129648
rect 496813 129643 496879 129646
rect 252461 129570 252527 129573
rect 248952 129568 252527 129570
rect 248952 129512 252466 129568
rect 252522 129512 252527 129568
rect 248952 129510 252527 129512
rect 252461 129507 252527 129510
rect 416773 129570 416839 129573
rect 416773 129568 420164 129570
rect 416773 129512 416778 129568
rect 416834 129512 420164 129568
rect 416773 129510 420164 129512
rect 416773 129507 416839 129510
rect 324313 129434 324379 129437
rect 321908 129432 324379 129434
rect 321908 129376 324318 129432
rect 324374 129376 324379 129432
rect 321908 129374 324379 129376
rect 324313 129371 324379 129374
rect 66069 129298 66135 129301
rect 68142 129298 68816 129304
rect 66069 129296 68816 129298
rect 66069 129240 66074 129296
rect 66130 129244 68816 129296
rect 307661 129298 307727 129301
rect 307661 129296 310040 129298
rect 66130 129240 68202 129244
rect 66069 129238 68202 129240
rect 66069 129235 66135 129238
rect 213913 128890 213979 128893
rect 217182 128890 217242 129268
rect 307661 129240 307666 129296
rect 307722 129240 310040 129296
rect 307661 129238 310040 129240
rect 307661 129235 307727 129238
rect 252369 129162 252435 129165
rect 248952 129160 252435 129162
rect 248952 129104 252374 129160
rect 252430 129104 252435 129160
rect 248952 129102 252435 129104
rect 252369 129099 252435 129102
rect 213913 128888 217242 128890
rect 213913 128832 213918 128888
rect 213974 128832 217242 128888
rect 213913 128830 217242 128832
rect 306925 128890 306991 128893
rect 306925 128888 310040 128890
rect 306925 128832 306930 128888
rect 306986 128832 310040 128888
rect 306925 128830 310040 128832
rect 213913 128827 213979 128830
rect 306925 128827 306991 128830
rect 170254 128556 170260 128620
rect 170324 128618 170330 128620
rect 170324 128558 200130 128618
rect 170324 128556 170330 128558
rect 200070 128482 200130 128558
rect 217366 128482 217426 128724
rect 288934 128692 288940 128756
rect 289004 128754 289010 128756
rect 289004 128694 296730 128754
rect 289004 128692 289010 128694
rect 252277 128618 252343 128621
rect 248952 128616 252343 128618
rect 248952 128560 252282 128616
rect 252338 128560 252343 128616
rect 248952 128558 252343 128560
rect 252277 128555 252343 128558
rect 200070 128422 217426 128482
rect 296670 128482 296730 128694
rect 324405 128618 324471 128621
rect 321908 128616 324471 128618
rect 321908 128560 324410 128616
rect 324466 128560 324471 128616
rect 321908 128558 324471 128560
rect 324405 128555 324471 128558
rect 496905 128482 496971 128485
rect 296670 128422 310040 128482
rect 494316 128480 496971 128482
rect 494316 128424 496910 128480
rect 496966 128424 496971 128480
rect 494316 128422 496971 128424
rect 496905 128419 496971 128422
rect 252461 128210 252527 128213
rect 248952 128208 252527 128210
rect 248952 128152 252466 128208
rect 252522 128152 252527 128208
rect 248952 128150 252527 128152
rect 252461 128147 252527 128150
rect 65517 128074 65583 128077
rect 68142 128074 68816 128080
rect 65517 128072 68816 128074
rect 65517 128016 65522 128072
rect 65578 128020 68816 128072
rect 307477 128074 307543 128077
rect 307477 128072 310040 128074
rect 65578 128016 68202 128020
rect 65517 128014 68202 128016
rect 65517 128011 65583 128014
rect 217182 127530 217242 128044
rect 307477 128016 307482 128072
rect 307538 128016 310040 128072
rect 307477 128014 310040 128016
rect 307477 128011 307543 128014
rect 419809 127938 419875 127941
rect 419809 127936 420164 127938
rect 419809 127880 419814 127936
rect 419870 127880 420164 127936
rect 419809 127878 420164 127880
rect 419809 127875 419875 127878
rect 494094 127876 494100 127940
rect 494164 127876 494170 127940
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 252277 127666 252343 127669
rect 248952 127664 252343 127666
rect 248952 127608 252282 127664
rect 252338 127608 252343 127664
rect 248952 127606 252343 127608
rect 252277 127603 252343 127606
rect 307569 127666 307635 127669
rect 307569 127664 310040 127666
rect 307569 127608 307574 127664
rect 307630 127608 310040 127664
rect 307569 127606 310040 127608
rect 307569 127603 307635 127606
rect 200070 127470 217242 127530
rect 166390 127060 166396 127124
rect 166460 127122 166466 127124
rect 200070 127122 200130 127470
rect 494102 127364 494162 127876
rect 166460 127062 200130 127122
rect 213913 127122 213979 127125
rect 217182 127122 217242 127364
rect 252369 127258 252435 127261
rect 248952 127256 252435 127258
rect 248952 127200 252374 127256
rect 252430 127200 252435 127256
rect 248952 127198 252435 127200
rect 252369 127195 252435 127198
rect 307661 127258 307727 127261
rect 307661 127256 310040 127258
rect 307661 127200 307666 127256
rect 307722 127200 310040 127256
rect 307661 127198 310040 127200
rect 307661 127195 307727 127198
rect 324405 127122 324471 127125
rect 213913 127120 217242 127122
rect 213913 127064 213918 127120
rect 213974 127064 217242 127120
rect 213913 127062 217242 127064
rect 321908 127120 324471 127122
rect 321908 127064 324410 127120
rect 324466 127064 324471 127120
rect 321908 127062 324471 127064
rect 166460 127060 166466 127062
rect 213913 127059 213979 127062
rect 324405 127059 324471 127062
rect 307569 126850 307635 126853
rect 307569 126848 310040 126850
rect 307569 126792 307574 126848
rect 307630 126792 310040 126848
rect 307569 126790 310040 126792
rect 307569 126787 307635 126790
rect 252461 126714 252527 126717
rect 248952 126712 252527 126714
rect 67357 126306 67423 126309
rect 68142 126306 68816 126312
rect 67357 126304 68816 126306
rect 67357 126248 67362 126304
rect 67418 126252 68816 126304
rect 67418 126248 68202 126252
rect 67357 126246 68202 126248
rect 67357 126243 67423 126246
rect 214005 126170 214071 126173
rect 217182 126170 217242 126684
rect 248952 126656 252466 126712
rect 252522 126656 252527 126712
rect 248952 126654 252527 126656
rect 252461 126651 252527 126654
rect 309550 126338 310132 126398
rect 252369 126306 252435 126309
rect 248952 126304 252435 126306
rect 248952 126248 252374 126304
rect 252430 126248 252435 126304
rect 248952 126246 252435 126248
rect 252369 126243 252435 126246
rect 214005 126168 217242 126170
rect 214005 126112 214010 126168
rect 214066 126112 217242 126168
rect 214005 126110 217242 126112
rect 214005 126107 214071 126110
rect 213913 125762 213979 125765
rect 217182 125762 217242 126004
rect 291694 125836 291700 125900
rect 291764 125898 291770 125900
rect 309550 125898 309610 126338
rect 327022 126306 327028 126308
rect 321908 126246 327028 126306
rect 327022 126244 327028 126246
rect 327092 126244 327098 126308
rect 496813 126306 496879 126309
rect 494316 126304 496879 126306
rect 494316 126248 496818 126304
rect 496874 126248 496879 126304
rect 494316 126246 496879 126248
rect 496813 126243 496879 126246
rect 418521 126170 418587 126173
rect 418521 126168 420164 126170
rect 418521 126112 418526 126168
rect 418582 126112 420164 126168
rect 418521 126110 420164 126112
rect 418521 126107 418587 126110
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 291764 125838 309610 125898
rect 583520 125884 584960 125974
rect 291764 125836 291770 125838
rect 309734 125794 310132 125854
rect 252277 125762 252343 125765
rect 213913 125760 217242 125762
rect 213913 125704 213918 125760
rect 213974 125704 217242 125760
rect 213913 125702 217242 125704
rect 248952 125760 252343 125762
rect 248952 125704 252282 125760
rect 252338 125704 252343 125760
rect 248952 125702 252343 125704
rect 213913 125699 213979 125702
rect 252277 125699 252343 125702
rect 307661 125762 307727 125765
rect 309734 125762 309794 125794
rect 307661 125760 309794 125762
rect 307661 125704 307666 125760
rect 307722 125704 309794 125760
rect 307661 125702 309794 125704
rect 307661 125699 307727 125702
rect 307477 125490 307543 125493
rect 324313 125490 324379 125493
rect 307477 125488 310040 125490
rect 307477 125432 307482 125488
rect 307538 125432 310040 125488
rect 307477 125430 310040 125432
rect 321908 125488 324379 125490
rect 321908 125432 324318 125488
rect 324374 125432 324379 125488
rect 321908 125430 324379 125432
rect 307477 125427 307543 125430
rect 324313 125427 324379 125430
rect 252461 125354 252527 125357
rect 248952 125352 252527 125354
rect 66161 125218 66227 125221
rect 68142 125218 68816 125224
rect 66161 125216 68816 125218
rect 66161 125160 66166 125216
rect 66222 125164 68816 125216
rect 66222 125160 68202 125164
rect 66161 125158 68202 125160
rect 66161 125155 66227 125158
rect 214005 124810 214071 124813
rect 217182 124810 217242 125324
rect 248952 125296 252466 125352
rect 252522 125296 252527 125352
rect 248952 125294 252527 125296
rect 252461 125291 252527 125294
rect 496813 125218 496879 125221
rect 494316 125216 496879 125218
rect 494316 125160 496818 125216
rect 496874 125160 496879 125216
rect 494316 125158 496879 125160
rect 496813 125155 496879 125158
rect 307569 125082 307635 125085
rect 307569 125080 310040 125082
rect 307569 125024 307574 125080
rect 307630 125024 310040 125080
rect 307569 125022 310040 125024
rect 307569 125019 307635 125022
rect 252001 124810 252067 124813
rect 324405 124810 324471 124813
rect 214005 124808 217242 124810
rect 214005 124752 214010 124808
rect 214066 124752 217242 124808
rect 214005 124750 217242 124752
rect 248952 124808 252067 124810
rect 248952 124752 252006 124808
rect 252062 124752 252067 124808
rect 248952 124750 252067 124752
rect 321908 124808 324471 124810
rect 321908 124752 324410 124808
rect 324466 124752 324471 124808
rect 321908 124750 324471 124752
rect 214005 124747 214071 124750
rect 252001 124747 252067 124750
rect 324405 124747 324471 124750
rect 307661 124674 307727 124677
rect 307661 124672 310040 124674
rect 213913 124402 213979 124405
rect 217182 124402 217242 124644
rect 307661 124616 307666 124672
rect 307722 124616 310040 124672
rect 307661 124614 310040 124616
rect 307661 124611 307727 124614
rect 418521 124538 418587 124541
rect 418521 124536 420164 124538
rect 418521 124480 418526 124536
rect 418582 124480 420164 124536
rect 418521 124478 420164 124480
rect 418521 124475 418587 124478
rect 252185 124402 252251 124405
rect 213913 124400 217242 124402
rect 213913 124344 213918 124400
rect 213974 124344 217242 124400
rect 213913 124342 217242 124344
rect 248952 124400 252251 124402
rect 248952 124344 252190 124400
rect 252246 124344 252251 124400
rect 248952 124342 252251 124344
rect 213913 124339 213979 124342
rect 252185 124339 252251 124342
rect 307661 124266 307727 124269
rect 307661 124264 310040 124266
rect 307661 124208 307666 124264
rect 307722 124208 310040 124264
rect 307661 124206 310040 124208
rect 307661 124203 307727 124206
rect 496813 124130 496879 124133
rect 494316 124128 496879 124130
rect -960 123572 480 123812
rect 67541 123586 67607 123589
rect 68142 123586 68816 123592
rect 67541 123584 68816 123586
rect 67541 123528 67546 123584
rect 67602 123532 68816 123584
rect 214005 123586 214071 123589
rect 217182 123586 217242 124100
rect 494316 124072 496818 124128
rect 496874 124072 496879 124128
rect 494316 124070 496879 124072
rect 496813 124067 496879 124070
rect 252461 123994 252527 123997
rect 324313 123994 324379 123997
rect 248952 123992 252527 123994
rect 248952 123936 252466 123992
rect 252522 123936 252527 123992
rect 248952 123934 252527 123936
rect 321908 123992 324379 123994
rect 321908 123936 324318 123992
rect 324374 123936 324379 123992
rect 321908 123934 324379 123936
rect 252461 123931 252527 123934
rect 324313 123931 324379 123934
rect 309550 123754 310132 123814
rect 309550 123722 309610 123754
rect 214005 123584 217242 123586
rect 67602 123528 68202 123532
rect 67541 123526 68202 123528
rect 214005 123528 214010 123584
rect 214066 123528 217242 123584
rect 214005 123526 217242 123528
rect 296670 123662 309610 123722
rect 67541 123523 67607 123526
rect 214005 123523 214071 123526
rect 252369 123450 252435 123453
rect 248952 123448 252435 123450
rect 213913 123178 213979 123181
rect 217182 123178 217242 123420
rect 248952 123392 252374 123448
rect 252430 123392 252435 123448
rect 248952 123390 252435 123392
rect 252369 123387 252435 123390
rect 213913 123176 217242 123178
rect 213913 123120 213918 123176
rect 213974 123120 217242 123176
rect 213913 123118 217242 123120
rect 213913 123115 213979 123118
rect 255814 123116 255820 123180
rect 255884 123178 255890 123180
rect 296670 123178 296730 123662
rect 307569 123450 307635 123453
rect 307569 123448 310040 123450
rect 307569 123392 307574 123448
rect 307630 123392 310040 123448
rect 307569 123390 310040 123392
rect 307569 123387 307635 123390
rect 324957 123178 325023 123181
rect 255884 123118 296730 123178
rect 321908 123176 325023 123178
rect 321908 123120 324962 123176
rect 325018 123120 325023 123176
rect 321908 123118 325023 123120
rect 255884 123116 255890 123118
rect 324957 123115 325023 123118
rect 252277 123042 252343 123045
rect 248952 123040 252343 123042
rect 248952 122984 252282 123040
rect 252338 122984 252343 123040
rect 248952 122982 252343 122984
rect 252277 122979 252343 122982
rect 307661 123042 307727 123045
rect 307661 123040 310040 123042
rect 307661 122984 307666 123040
rect 307722 122984 310040 123040
rect 307661 122982 310040 122984
rect 307661 122979 307727 122982
rect 496905 122906 496971 122909
rect 494316 122904 496971 122906
rect 494316 122848 496910 122904
rect 496966 122848 496971 122904
rect 494316 122846 496971 122848
rect 496905 122843 496971 122846
rect 419533 122770 419599 122773
rect 419533 122768 420164 122770
rect 67449 122634 67515 122637
rect 68142 122634 68816 122640
rect 67449 122632 68816 122634
rect 67449 122576 67454 122632
rect 67510 122580 68816 122632
rect 67510 122576 68202 122580
rect 67449 122574 68202 122576
rect 67449 122571 67515 122574
rect 214005 122226 214071 122229
rect 217182 122226 217242 122740
rect 419533 122712 419538 122768
rect 419594 122712 420164 122768
rect 419533 122710 420164 122712
rect 419533 122707 419599 122710
rect 252461 122498 252527 122501
rect 248952 122496 252527 122498
rect 248952 122440 252466 122496
rect 252522 122440 252527 122496
rect 248952 122438 252527 122440
rect 252461 122435 252527 122438
rect 307569 122498 307635 122501
rect 324313 122498 324379 122501
rect 307569 122496 310040 122498
rect 307569 122440 307574 122496
rect 307630 122440 310040 122496
rect 307569 122438 310040 122440
rect 321908 122496 324379 122498
rect 321908 122440 324318 122496
rect 324374 122440 324379 122496
rect 321908 122438 324379 122440
rect 307569 122435 307635 122438
rect 324313 122435 324379 122438
rect 214005 122224 217242 122226
rect 214005 122168 214010 122224
rect 214066 122168 217242 122224
rect 214005 122166 217242 122168
rect 214005 122163 214071 122166
rect 252369 122090 252435 122093
rect 248952 122088 252435 122090
rect 213913 121546 213979 121549
rect 217182 121546 217242 122060
rect 248952 122032 252374 122088
rect 252430 122032 252435 122088
rect 248952 122030 252435 122032
rect 252369 122027 252435 122030
rect 306741 122090 306807 122093
rect 306741 122088 310040 122090
rect 306741 122032 306746 122088
rect 306802 122032 310040 122088
rect 306741 122030 310040 122032
rect 306741 122027 306807 122030
rect 495617 121818 495683 121821
rect 494316 121816 495683 121818
rect 494316 121760 495622 121816
rect 495678 121760 495683 121816
rect 494316 121758 495683 121760
rect 495617 121755 495683 121758
rect 307661 121682 307727 121685
rect 323117 121682 323183 121685
rect 307661 121680 310040 121682
rect 307661 121624 307666 121680
rect 307722 121624 310040 121680
rect 307661 121622 310040 121624
rect 321908 121680 323183 121682
rect 321908 121624 323122 121680
rect 323178 121624 323183 121680
rect 321908 121622 323183 121624
rect 307661 121619 307727 121622
rect 323117 121619 323183 121622
rect 252277 121546 252343 121549
rect 213913 121544 217242 121546
rect 213913 121488 213918 121544
rect 213974 121488 217242 121544
rect 213913 121486 217242 121488
rect 248952 121544 252343 121546
rect 248952 121488 252282 121544
rect 252338 121488 252343 121544
rect 248952 121486 252343 121488
rect 213913 121483 213979 121486
rect 252277 121483 252343 121486
rect 67633 120866 67699 120869
rect 68142 120866 68816 120872
rect 67633 120864 68816 120866
rect 67633 120808 67638 120864
rect 67694 120812 68816 120864
rect 213913 120866 213979 120869
rect 217182 120866 217242 121380
rect 307293 121274 307359 121277
rect 307293 121272 310040 121274
rect 307293 121216 307298 121272
rect 307354 121216 310040 121272
rect 307293 121214 310040 121216
rect 307293 121211 307359 121214
rect 252093 121138 252159 121141
rect 248952 121136 252159 121138
rect 248952 121080 252098 121136
rect 252154 121080 252159 121136
rect 248952 121078 252159 121080
rect 252093 121075 252159 121078
rect 417509 121138 417575 121141
rect 417509 121136 420164 121138
rect 417509 121080 417514 121136
rect 417570 121080 420164 121136
rect 417509 121078 420164 121080
rect 417509 121075 417575 121078
rect 213913 120864 217242 120866
rect 67694 120808 68202 120812
rect 67633 120806 68202 120808
rect 213913 120808 213918 120864
rect 213974 120808 217242 120864
rect 213913 120806 217242 120808
rect 307569 120866 307635 120869
rect 324313 120866 324379 120869
rect 307569 120864 310040 120866
rect 307569 120808 307574 120864
rect 307630 120808 310040 120864
rect 307569 120806 310040 120808
rect 321908 120864 324379 120866
rect 321908 120808 324318 120864
rect 324374 120808 324379 120864
rect 321908 120806 324379 120808
rect 67633 120803 67699 120806
rect 213913 120803 213979 120806
rect 307569 120803 307635 120806
rect 324313 120803 324379 120806
rect 496813 120730 496879 120733
rect 494316 120728 496879 120730
rect 214005 120322 214071 120325
rect 217182 120322 217242 120700
rect 494316 120672 496818 120728
rect 496874 120672 496879 120728
rect 494316 120670 496879 120672
rect 496813 120667 496879 120670
rect 252461 120594 252527 120597
rect 248952 120592 252527 120594
rect 248952 120536 252466 120592
rect 252522 120536 252527 120592
rect 248952 120534 252527 120536
rect 252461 120531 252527 120534
rect 307661 120458 307727 120461
rect 307661 120456 310040 120458
rect 307661 120400 307666 120456
rect 307722 120400 310040 120456
rect 307661 120398 310040 120400
rect 307661 120395 307727 120398
rect 214005 120320 217242 120322
rect 214005 120264 214010 120320
rect 214066 120264 217242 120320
rect 214005 120262 217242 120264
rect 214005 120259 214071 120262
rect 251909 120186 251975 120189
rect 324405 120186 324471 120189
rect 248952 120184 251975 120186
rect 248952 120128 251914 120184
rect 251970 120128 251975 120184
rect 248952 120126 251975 120128
rect 321908 120184 324471 120186
rect 321908 120128 324410 120184
rect 324466 120128 324471 120184
rect 321908 120126 324471 120128
rect 251909 120123 251975 120126
rect 324405 120123 324471 120126
rect 306557 120050 306623 120053
rect 306557 120048 310040 120050
rect 214005 119642 214071 119645
rect 217182 119642 217242 120020
rect 306557 119992 306562 120048
rect 306618 119992 310040 120048
rect 306557 119990 310040 119992
rect 306557 119987 306623 119990
rect 321645 119914 321711 119917
rect 321645 119912 321754 119914
rect 321645 119856 321650 119912
rect 321706 119856 321754 119912
rect 321645 119851 321754 119856
rect 252461 119642 252527 119645
rect 214005 119640 217242 119642
rect 214005 119584 214010 119640
rect 214066 119584 217242 119640
rect 214005 119582 217242 119584
rect 248952 119640 252527 119642
rect 248952 119584 252466 119640
rect 252522 119584 252527 119640
rect 248952 119582 252527 119584
rect 214005 119579 214071 119582
rect 252461 119579 252527 119582
rect 307661 119642 307727 119645
rect 307661 119640 310040 119642
rect 307661 119584 307666 119640
rect 307722 119584 310040 119640
rect 307661 119582 310040 119584
rect 307661 119579 307727 119582
rect 214097 119098 214163 119101
rect 217182 119098 217242 119476
rect 321694 119340 321754 119851
rect 496813 119642 496879 119645
rect 494316 119640 496879 119642
rect 494316 119584 496818 119640
rect 496874 119584 496879 119640
rect 494316 119582 496879 119584
rect 496813 119579 496879 119582
rect 416773 119370 416839 119373
rect 416773 119368 420164 119370
rect 416773 119312 416778 119368
rect 416834 119312 420164 119368
rect 416773 119310 420164 119312
rect 416773 119307 416839 119310
rect 252277 119234 252343 119237
rect 248952 119232 252343 119234
rect 248952 119176 252282 119232
rect 252338 119176 252343 119232
rect 248952 119174 252343 119176
rect 252277 119171 252343 119174
rect 214097 119096 217242 119098
rect 214097 119040 214102 119096
rect 214158 119040 217242 119096
rect 214097 119038 217242 119040
rect 214097 119035 214163 119038
rect 309550 118994 310132 119054
rect 213913 118962 213979 118965
rect 305729 118962 305795 118965
rect 309550 118962 309610 118994
rect 213913 118960 217242 118962
rect 213913 118904 213918 118960
rect 213974 118904 217242 118960
rect 213913 118902 217242 118904
rect 213913 118899 213979 118902
rect 217182 118796 217242 118902
rect 305729 118960 309610 118962
rect 305729 118904 305734 118960
rect 305790 118904 309610 118960
rect 305729 118902 309610 118904
rect 305729 118899 305795 118902
rect 252369 118826 252435 118829
rect 248952 118824 252435 118826
rect 248952 118768 252374 118824
rect 252430 118768 252435 118824
rect 248952 118766 252435 118768
rect 252369 118763 252435 118766
rect 307569 118690 307635 118693
rect 307569 118688 310040 118690
rect 307569 118632 307574 118688
rect 307630 118632 310040 118688
rect 307569 118630 310040 118632
rect 307569 118627 307635 118630
rect 324313 118554 324379 118557
rect 321908 118552 324379 118554
rect 321908 118496 324318 118552
rect 324374 118496 324379 118552
rect 321908 118494 324379 118496
rect 324313 118491 324379 118494
rect 496813 118418 496879 118421
rect 494316 118416 496879 118418
rect 494316 118360 496818 118416
rect 496874 118360 496879 118416
rect 494316 118358 496879 118360
rect 496813 118355 496879 118358
rect 252461 118282 252527 118285
rect 248952 118280 252527 118282
rect 248952 118224 252466 118280
rect 252522 118224 252527 118280
rect 248952 118222 252527 118224
rect 252461 118219 252527 118222
rect 307293 118282 307359 118285
rect 307293 118280 310040 118282
rect 307293 118224 307298 118280
rect 307354 118224 310040 118280
rect 307293 118222 310040 118224
rect 307293 118219 307359 118222
rect 214005 117602 214071 117605
rect 217182 117602 217242 118116
rect 252369 117874 252435 117877
rect 324405 117874 324471 117877
rect 248952 117872 252435 117874
rect 248952 117816 252374 117872
rect 252430 117816 252435 117872
rect 321908 117872 324471 117874
rect 248952 117814 252435 117816
rect 252369 117811 252435 117814
rect 309550 117770 310132 117830
rect 321908 117816 324410 117872
rect 324466 117816 324471 117872
rect 321908 117814 324471 117816
rect 324405 117811 324471 117814
rect 214005 117600 217242 117602
rect 214005 117544 214010 117600
rect 214066 117544 217242 117600
rect 214005 117542 217242 117544
rect 305821 117602 305887 117605
rect 309550 117602 309610 117770
rect 416957 117738 417023 117741
rect 416957 117736 420164 117738
rect 416957 117680 416962 117736
rect 417018 117680 420164 117736
rect 416957 117678 420164 117680
rect 416957 117675 417023 117678
rect 305821 117600 309610 117602
rect 305821 117544 305826 117600
rect 305882 117544 309610 117600
rect 305821 117542 309610 117544
rect 214005 117539 214071 117542
rect 305821 117539 305887 117542
rect 307661 117466 307727 117469
rect 307661 117464 310040 117466
rect 213913 117330 213979 117333
rect 213913 117328 216874 117330
rect 213913 117272 213918 117328
rect 213974 117272 216874 117328
rect 213913 117270 216874 117272
rect 213913 117267 213979 117270
rect 216814 117194 216874 117270
rect 217366 117194 217426 117436
rect 307661 117408 307666 117464
rect 307722 117408 310040 117464
rect 307661 117406 310040 117408
rect 307661 117403 307727 117406
rect 252277 117330 252343 117333
rect 496905 117330 496971 117333
rect 248952 117328 252343 117330
rect 248952 117272 252282 117328
rect 252338 117272 252343 117328
rect 248952 117270 252343 117272
rect 494316 117328 496971 117330
rect 494316 117272 496910 117328
rect 496966 117272 496971 117328
rect 494316 117270 496971 117272
rect 252277 117267 252343 117270
rect 496905 117267 496971 117270
rect 216814 117134 217426 117194
rect 307477 117058 307543 117061
rect 307477 117056 310040 117058
rect 307477 117000 307482 117056
rect 307538 117000 310040 117056
rect 307477 116998 310040 117000
rect 307477 116995 307543 116998
rect 251766 116922 251772 116924
rect 248952 116862 251772 116922
rect 251766 116860 251772 116862
rect 251836 116860 251842 116924
rect 214005 116242 214071 116245
rect 217182 116242 217242 116756
rect 307569 116650 307635 116653
rect 307569 116648 310040 116650
rect 307569 116592 307574 116648
rect 307630 116592 310040 116648
rect 307569 116590 310040 116592
rect 307569 116587 307635 116590
rect 321878 116514 321938 117028
rect 331438 116514 331444 116516
rect 321878 116454 331444 116514
rect 331438 116452 331444 116454
rect 331508 116452 331514 116516
rect 252461 116378 252527 116381
rect 324313 116378 324379 116381
rect 248952 116376 252527 116378
rect 248952 116320 252466 116376
rect 252522 116320 252527 116376
rect 248952 116318 252527 116320
rect 321908 116376 324379 116378
rect 321908 116320 324318 116376
rect 324374 116320 324379 116376
rect 321908 116318 324379 116320
rect 252461 116315 252527 116318
rect 324313 116315 324379 116318
rect 214005 116240 217242 116242
rect 214005 116184 214010 116240
rect 214066 116184 217242 116240
rect 214005 116182 217242 116184
rect 307661 116242 307727 116245
rect 496997 116242 497063 116245
rect 307661 116240 310040 116242
rect 307661 116184 307666 116240
rect 307722 116184 310040 116240
rect 307661 116182 310040 116184
rect 494316 116240 497063 116242
rect 494316 116184 497002 116240
rect 497058 116184 497063 116240
rect 494316 116182 497063 116184
rect 214005 116179 214071 116182
rect 307661 116179 307727 116182
rect 496997 116179 497063 116182
rect 213913 115970 213979 115973
rect 213913 115968 216874 115970
rect 213913 115912 213918 115968
rect 213974 115912 216874 115968
rect 213913 115910 216874 115912
rect 213913 115907 213979 115910
rect 216814 115834 216874 115910
rect 217366 115834 217426 116076
rect 252369 115970 252435 115973
rect 248952 115968 252435 115970
rect 248952 115912 252374 115968
rect 252430 115912 252435 115968
rect 248952 115910 252435 115912
rect 252369 115907 252435 115910
rect 338614 115908 338620 115972
rect 338684 115970 338690 115972
rect 420134 115970 420194 116076
rect 338684 115910 420194 115970
rect 338684 115908 338690 115910
rect 216814 115774 217426 115834
rect 307293 115698 307359 115701
rect 307293 115696 310040 115698
rect 307293 115640 307298 115696
rect 307354 115640 310040 115696
rect 307293 115638 310040 115640
rect 307293 115635 307359 115638
rect 324313 115562 324379 115565
rect 321908 115560 324379 115562
rect 321908 115504 324318 115560
rect 324374 115504 324379 115560
rect 321908 115502 324379 115504
rect 324313 115499 324379 115502
rect 252461 115426 252527 115429
rect 248952 115424 252527 115426
rect 214005 115018 214071 115021
rect 217182 115018 217242 115396
rect 248952 115368 252466 115424
rect 252522 115368 252527 115424
rect 248952 115366 252527 115368
rect 252461 115363 252527 115366
rect 307569 115290 307635 115293
rect 307569 115288 310040 115290
rect 307569 115232 307574 115288
rect 307630 115232 310040 115288
rect 307569 115230 310040 115232
rect 307569 115227 307635 115230
rect 496813 115154 496879 115157
rect 494316 115152 496879 115154
rect 494316 115096 496818 115152
rect 496874 115096 496879 115152
rect 494316 115094 496879 115096
rect 496813 115091 496879 115094
rect 252369 115018 252435 115021
rect 214005 115016 217242 115018
rect 214005 114960 214010 115016
rect 214066 114960 217242 115016
rect 214005 114958 217242 114960
rect 248952 115016 252435 115018
rect 248952 114960 252374 115016
rect 252430 114960 252435 115016
rect 248952 114958 252435 114960
rect 214005 114955 214071 114958
rect 252369 114955 252435 114958
rect 307661 114882 307727 114885
rect 307661 114880 310040 114882
rect 213913 114610 213979 114613
rect 217182 114610 217242 114852
rect 307661 114824 307666 114880
rect 307722 114824 310040 114880
rect 307661 114822 310040 114824
rect 307661 114819 307727 114822
rect 324405 114746 324471 114749
rect 321908 114744 324471 114746
rect 321908 114688 324410 114744
rect 324466 114688 324471 114744
rect 321908 114686 324471 114688
rect 324405 114683 324471 114686
rect 213913 114608 217242 114610
rect 213913 114552 213918 114608
rect 213974 114552 217242 114608
rect 213913 114550 217242 114552
rect 213913 114547 213979 114550
rect 252461 114474 252527 114477
rect 248952 114472 252527 114474
rect 248952 114416 252466 114472
rect 252522 114416 252527 114472
rect 248952 114414 252527 114416
rect 252461 114411 252527 114414
rect 306557 114474 306623 114477
rect 306557 114472 310040 114474
rect 306557 114416 306562 114472
rect 306618 114416 310040 114472
rect 306557 114414 310040 114416
rect 306557 114411 306623 114414
rect 416773 114338 416839 114341
rect 416773 114336 420164 114338
rect 416773 114280 416778 114336
rect 416834 114280 420164 114336
rect 416773 114278 420164 114280
rect 416773 114275 416839 114278
rect 214005 113658 214071 113661
rect 217182 113658 217242 114172
rect 253197 114066 253263 114069
rect 248952 114064 253263 114066
rect 248952 114008 253202 114064
rect 253258 114008 253263 114064
rect 248952 114006 253263 114008
rect 253197 114003 253263 114006
rect 309317 114066 309383 114069
rect 309317 114064 310040 114066
rect 309317 114008 309322 114064
rect 309378 114008 310040 114064
rect 309317 114006 310040 114008
rect 309317 114003 309383 114006
rect 321878 113661 321938 114036
rect 496813 113930 496879 113933
rect 494316 113928 496879 113930
rect 494316 113872 496818 113928
rect 496874 113872 496879 113928
rect 494316 113870 496879 113872
rect 496813 113867 496879 113870
rect 214005 113656 217242 113658
rect 214005 113600 214010 113656
rect 214066 113600 217242 113656
rect 214005 113598 217242 113600
rect 214005 113595 214071 113598
rect 307150 113596 307156 113660
rect 307220 113658 307226 113660
rect 307220 113598 310040 113658
rect 321829 113656 321938 113661
rect 321829 113600 321834 113656
rect 321890 113600 321938 113656
rect 321829 113598 321938 113600
rect 307220 113596 307226 113598
rect 321829 113595 321895 113598
rect 252277 113522 252343 113525
rect 248952 113520 252343 113522
rect 213913 113250 213979 113253
rect 217182 113250 217242 113492
rect 248952 113464 252282 113520
rect 252338 113464 252343 113520
rect 248952 113462 252343 113464
rect 252277 113459 252343 113462
rect 304390 113460 304396 113524
rect 304460 113522 304466 113524
rect 304460 113462 309380 113522
rect 304460 113460 304466 113462
rect 213913 113248 217242 113250
rect 213913 113192 213918 113248
rect 213974 113192 217242 113248
rect 213913 113190 217242 113192
rect 307661 113250 307727 113253
rect 309320 113250 309380 113462
rect 324313 113250 324379 113253
rect 307661 113248 309150 113250
rect 307661 113192 307666 113248
rect 307722 113192 309150 113248
rect 307661 113190 309150 113192
rect 309320 113190 310040 113250
rect 321908 113248 324379 113250
rect 321908 113192 324318 113248
rect 324374 113192 324379 113248
rect 321908 113190 324379 113192
rect 213913 113187 213979 113190
rect 307661 113187 307727 113190
rect 252277 113114 252343 113117
rect 248952 113112 252343 113114
rect 248952 113056 252282 113112
rect 252338 113056 252343 113112
rect 248952 113054 252343 113056
rect 309090 113114 309150 113190
rect 324313 113187 324379 113190
rect 309317 113114 309383 113117
rect 309090 113112 309383 113114
rect 309090 113056 309322 113112
rect 309378 113056 309383 113112
rect 309090 113054 309383 113056
rect 252277 113051 252343 113054
rect 309317 113051 309383 113054
rect 496813 112842 496879 112845
rect 494316 112840 496879 112842
rect 213453 112298 213519 112301
rect 217182 112298 217242 112812
rect 494316 112784 496818 112840
rect 496874 112784 496879 112840
rect 494316 112782 496879 112784
rect 496813 112779 496879 112782
rect 580257 112842 580323 112845
rect 583520 112842 584960 112932
rect 580257 112840 584960 112842
rect 580257 112784 580262 112840
rect 580318 112784 584960 112840
rect 580257 112782 584960 112784
rect 580257 112779 580323 112782
rect 252369 112706 252435 112709
rect 248952 112704 252435 112706
rect 248952 112648 252374 112704
rect 252430 112648 252435 112704
rect 248952 112646 252435 112648
rect 252369 112643 252435 112646
rect 307477 112706 307543 112709
rect 416773 112706 416839 112709
rect 307477 112704 310040 112706
rect 307477 112648 307482 112704
rect 307538 112648 310040 112704
rect 307477 112646 310040 112648
rect 416773 112704 420164 112706
rect 416773 112648 416778 112704
rect 416834 112648 420164 112704
rect 583520 112692 584960 112782
rect 416773 112646 420164 112648
rect 307477 112643 307543 112646
rect 416773 112643 416839 112646
rect 324313 112434 324379 112437
rect 321908 112432 324379 112434
rect 321908 112376 324318 112432
rect 324374 112376 324379 112432
rect 321908 112374 324379 112376
rect 324313 112371 324379 112374
rect 213453 112296 217242 112298
rect 213453 112240 213458 112296
rect 213514 112240 217242 112296
rect 213453 112238 217242 112240
rect 307569 112298 307635 112301
rect 307569 112296 310040 112298
rect 307569 112240 307574 112296
rect 307630 112240 310040 112296
rect 307569 112238 310040 112240
rect 213453 112235 213519 112238
rect 307569 112235 307635 112238
rect 252461 112162 252527 112165
rect 248952 112160 252527 112162
rect 213913 111890 213979 111893
rect 217182 111890 217242 112132
rect 248952 112104 252466 112160
rect 252522 112104 252527 112160
rect 248952 112102 252527 112104
rect 252461 112099 252527 112102
rect 213913 111888 217242 111890
rect 213913 111832 213918 111888
rect 213974 111832 217242 111888
rect 213913 111830 217242 111832
rect 307661 111890 307727 111893
rect 307661 111888 310040 111890
rect 307661 111832 307666 111888
rect 307722 111832 310040 111888
rect 307661 111830 310040 111832
rect 213913 111827 213979 111830
rect 307661 111827 307727 111830
rect 168005 111754 168071 111757
rect 252369 111754 252435 111757
rect 322933 111754 322999 111757
rect 496813 111754 496879 111757
rect 164694 111752 168071 111754
rect 164694 111696 168010 111752
rect 168066 111696 168071 111752
rect 164694 111694 168071 111696
rect 248952 111752 252435 111754
rect 248952 111696 252374 111752
rect 252430 111696 252435 111752
rect 248952 111694 252435 111696
rect 321908 111752 322999 111754
rect 321908 111696 322938 111752
rect 322994 111696 322999 111752
rect 321908 111694 322999 111696
rect 494316 111752 496879 111754
rect 494316 111696 496818 111752
rect 496874 111696 496879 111752
rect 494316 111694 496879 111696
rect 168005 111691 168071 111694
rect 252369 111691 252435 111694
rect 322933 111691 322999 111694
rect 496813 111691 496879 111694
rect 307293 111482 307359 111485
rect 307293 111480 310040 111482
rect 214005 110938 214071 110941
rect 217182 110938 217242 111452
rect 307293 111424 307298 111480
rect 307354 111424 310040 111480
rect 307293 111422 310040 111424
rect 307293 111419 307359 111422
rect 251173 111210 251239 111213
rect 248952 111208 251239 111210
rect 248952 111152 251178 111208
rect 251234 111152 251239 111208
rect 248952 111150 251239 111152
rect 251173 111147 251239 111150
rect 252502 111012 252508 111076
rect 252572 111074 252578 111076
rect 293401 111074 293467 111077
rect 252572 111072 293467 111074
rect 252572 111016 293406 111072
rect 293462 111016 293467 111072
rect 252572 111014 293467 111016
rect 252572 111012 252578 111014
rect 293401 111011 293467 111014
rect 306741 111074 306807 111077
rect 306741 111072 310040 111074
rect 306741 111016 306746 111072
rect 306802 111016 310040 111072
rect 306741 111014 310040 111016
rect 306741 111011 306807 111014
rect 214005 110936 217242 110938
rect 214005 110880 214010 110936
rect 214066 110880 217242 110936
rect 416773 110938 416839 110941
rect 416773 110936 420164 110938
rect 214005 110878 217242 110880
rect 214005 110875 214071 110878
rect 252461 110802 252527 110805
rect 248952 110800 252527 110802
rect -960 110666 480 110756
rect 3693 110666 3759 110669
rect -960 110664 3759 110666
rect -960 110608 3698 110664
rect 3754 110608 3759 110664
rect -960 110606 3759 110608
rect -960 110516 480 110606
rect 3693 110603 3759 110606
rect 213913 110530 213979 110533
rect 217366 110530 217426 110772
rect 248952 110744 252466 110800
rect 252522 110744 252527 110800
rect 248952 110742 252527 110744
rect 252461 110739 252527 110742
rect 307661 110666 307727 110669
rect 321878 110666 321938 110908
rect 416773 110880 416778 110936
rect 416834 110880 420164 110936
rect 416773 110878 420164 110880
rect 416773 110875 416839 110878
rect 334198 110666 334204 110668
rect 307661 110664 310040 110666
rect 307661 110608 307666 110664
rect 307722 110608 310040 110664
rect 307661 110606 310040 110608
rect 321878 110606 334204 110666
rect 307661 110603 307727 110606
rect 334198 110604 334204 110606
rect 334268 110604 334274 110668
rect 496905 110666 496971 110669
rect 494316 110664 496971 110666
rect 494316 110608 496910 110664
rect 496966 110608 496971 110664
rect 494316 110606 496971 110608
rect 496905 110603 496971 110606
rect 213913 110528 217426 110530
rect 213913 110472 213918 110528
rect 213974 110472 217426 110528
rect 213913 110470 217426 110472
rect 213913 110467 213979 110470
rect 252461 110258 252527 110261
rect 248952 110256 252527 110258
rect 168097 110122 168163 110125
rect 164694 110120 168163 110122
rect 164694 110064 168102 110120
rect 168158 110064 168163 110120
rect 164694 110062 168163 110064
rect 168097 110059 168163 110062
rect 214741 109714 214807 109717
rect 217182 109714 217242 110228
rect 248952 110200 252466 110256
rect 252522 110200 252527 110256
rect 248952 110198 252527 110200
rect 252461 110195 252527 110198
rect 307569 110258 307635 110261
rect 307569 110256 310040 110258
rect 307569 110200 307574 110256
rect 307630 110200 310040 110256
rect 307569 110198 310040 110200
rect 307569 110195 307635 110198
rect 252502 109850 252508 109852
rect 248952 109790 252508 109850
rect 252502 109788 252508 109790
rect 252572 109788 252578 109852
rect 306925 109850 306991 109853
rect 306925 109848 310040 109850
rect 306925 109792 306930 109848
rect 306986 109792 310040 109848
rect 306925 109790 310040 109792
rect 306925 109787 306991 109790
rect 214741 109712 217242 109714
rect 214741 109656 214746 109712
rect 214802 109656 217242 109712
rect 214741 109654 217242 109656
rect 214741 109651 214807 109654
rect 321878 109578 321938 110092
rect 213913 109306 213979 109309
rect 217182 109306 217242 109548
rect 321878 109518 325710 109578
rect 324313 109442 324379 109445
rect 321908 109440 324379 109442
rect 321908 109384 324318 109440
rect 324374 109384 324379 109440
rect 321908 109382 324379 109384
rect 324313 109379 324379 109382
rect 251725 109306 251791 109309
rect 213913 109304 217242 109306
rect 213913 109248 213918 109304
rect 213974 109248 217242 109304
rect 213913 109246 217242 109248
rect 248952 109304 251791 109306
rect 248952 109248 251730 109304
rect 251786 109248 251791 109304
rect 248952 109246 251791 109248
rect 213913 109243 213979 109246
rect 251725 109243 251791 109246
rect 307661 109306 307727 109309
rect 307661 109304 310040 109306
rect 307661 109248 307666 109304
rect 307722 109248 310040 109304
rect 307661 109246 310040 109248
rect 307661 109243 307727 109246
rect 325650 109170 325710 109518
rect 496813 109442 496879 109445
rect 494316 109440 496879 109442
rect 494316 109384 496818 109440
rect 496874 109384 496879 109440
rect 494316 109382 496879 109384
rect 496813 109379 496879 109382
rect 417417 109306 417483 109309
rect 417417 109304 420164 109306
rect 417417 109248 417422 109304
rect 417478 109248 420164 109304
rect 417417 109246 420164 109248
rect 417417 109243 417483 109246
rect 339534 109170 339540 109172
rect 325650 109110 339540 109170
rect 339534 109108 339540 109110
rect 339604 109108 339610 109172
rect 252461 108898 252527 108901
rect 248952 108896 252527 108898
rect 167637 108762 167703 108765
rect 164694 108760 167703 108762
rect 164694 108704 167642 108760
rect 167698 108704 167703 108760
rect 164694 108702 167703 108704
rect 167637 108699 167703 108702
rect 214005 108354 214071 108357
rect 217182 108354 217242 108868
rect 248952 108840 252466 108896
rect 252522 108840 252527 108896
rect 248952 108838 252527 108840
rect 252461 108835 252527 108838
rect 307477 108898 307543 108901
rect 307477 108896 310040 108898
rect 307477 108840 307482 108896
rect 307538 108840 310040 108896
rect 307477 108838 310040 108840
rect 307477 108835 307543 108838
rect 324313 108626 324379 108629
rect 321908 108624 324379 108626
rect 321908 108568 324318 108624
rect 324374 108568 324379 108624
rect 321908 108566 324379 108568
rect 324313 108563 324379 108566
rect 309550 108386 310132 108446
rect 252369 108354 252435 108357
rect 214005 108352 217242 108354
rect 214005 108296 214010 108352
rect 214066 108296 217242 108352
rect 214005 108294 217242 108296
rect 248952 108352 252435 108354
rect 248952 108296 252374 108352
rect 252430 108296 252435 108352
rect 248952 108294 252435 108296
rect 214005 108291 214071 108294
rect 252369 108291 252435 108294
rect 213913 107946 213979 107949
rect 217182 107946 217242 108188
rect 251909 107946 251975 107949
rect 213913 107944 217242 107946
rect 213913 107888 213918 107944
rect 213974 107888 217242 107944
rect 213913 107886 217242 107888
rect 248952 107944 251975 107946
rect 248952 107888 251914 107944
rect 251970 107888 251975 107944
rect 248952 107886 251975 107888
rect 213913 107883 213979 107886
rect 251909 107883 251975 107886
rect 305913 107946 305979 107949
rect 309550 107946 309610 108386
rect 496997 108354 497063 108357
rect 494316 108352 497063 108354
rect 494316 108296 497002 108352
rect 497058 108296 497063 108352
rect 494316 108294 497063 108296
rect 496997 108291 497063 108294
rect 305913 107944 309610 107946
rect 305913 107888 305918 107944
rect 305974 107888 309610 107944
rect 305913 107886 309610 107888
rect 309734 107978 310132 108038
rect 305913 107883 305979 107886
rect 307569 107810 307635 107813
rect 309734 107810 309794 107978
rect 325601 107810 325667 107813
rect 307569 107808 309794 107810
rect 307569 107752 307574 107808
rect 307630 107752 309794 107808
rect 307569 107750 309794 107752
rect 321908 107808 325667 107810
rect 321908 107752 325606 107808
rect 325662 107752 325667 107808
rect 321908 107750 325667 107752
rect 307569 107747 307635 107750
rect 325601 107747 325667 107750
rect 307661 107674 307727 107677
rect 307661 107672 310040 107674
rect 307661 107616 307666 107672
rect 307722 107616 310040 107672
rect 307661 107614 310040 107616
rect 307661 107611 307727 107614
rect 252461 107538 252527 107541
rect 248952 107536 252527 107538
rect 214005 106994 214071 106997
rect 217182 106994 217242 107508
rect 248952 107480 252466 107536
rect 252522 107480 252527 107536
rect 248952 107478 252527 107480
rect 252461 107475 252527 107478
rect 416773 107538 416839 107541
rect 416773 107536 420164 107538
rect 416773 107480 416778 107536
rect 416834 107480 420164 107536
rect 416773 107478 420164 107480
rect 416773 107475 416839 107478
rect 307661 107266 307727 107269
rect 497089 107266 497155 107269
rect 307661 107264 310040 107266
rect 307661 107208 307666 107264
rect 307722 107208 310040 107264
rect 307661 107206 310040 107208
rect 494316 107264 497155 107266
rect 494316 107208 497094 107264
rect 497150 107208 497155 107264
rect 494316 107206 497155 107208
rect 307661 107203 307727 107206
rect 497089 107203 497155 107206
rect 326654 107130 326660 107132
rect 321908 107070 326660 107130
rect 326654 107068 326660 107070
rect 326724 107068 326730 107132
rect 252369 106994 252435 106997
rect 214005 106992 217242 106994
rect 214005 106936 214010 106992
rect 214066 106936 217242 106992
rect 214005 106934 217242 106936
rect 248952 106992 252435 106994
rect 248952 106936 252374 106992
rect 252430 106936 252435 106992
rect 248952 106934 252435 106936
rect 214005 106931 214071 106934
rect 252369 106931 252435 106934
rect 306741 106858 306807 106861
rect 306741 106856 310040 106858
rect 213913 106450 213979 106453
rect 217182 106450 217242 106828
rect 306741 106800 306746 106856
rect 306802 106800 310040 106856
rect 306741 106798 310040 106800
rect 306741 106795 306807 106798
rect 252461 106586 252527 106589
rect 248952 106584 252527 106586
rect 248952 106528 252466 106584
rect 252522 106528 252527 106584
rect 248952 106526 252527 106528
rect 252461 106523 252527 106526
rect 213913 106448 217242 106450
rect 213913 106392 213918 106448
rect 213974 106392 217242 106448
rect 213913 106390 217242 106392
rect 307477 106450 307543 106453
rect 307477 106448 310040 106450
rect 307477 106392 307482 106448
rect 307538 106392 310040 106448
rect 307477 106390 310040 106392
rect 213913 106387 213979 106390
rect 307477 106387 307543 106390
rect 328494 106314 328500 106316
rect 321908 106254 328500 106314
rect 328494 106252 328500 106254
rect 328564 106252 328570 106316
rect 496813 106178 496879 106181
rect 494316 106176 496879 106178
rect 214005 105770 214071 105773
rect 217182 105770 217242 106148
rect 494316 106120 496818 106176
rect 496874 106120 496879 106176
rect 494316 106118 496879 106120
rect 496813 106115 496879 106118
rect 250713 106042 250779 106045
rect 248952 106040 250779 106042
rect 248952 105984 250718 106040
rect 250774 105984 250779 106040
rect 248952 105982 250779 105984
rect 250713 105979 250779 105982
rect 307569 105906 307635 105909
rect 416773 105906 416839 105909
rect 307569 105904 310040 105906
rect 307569 105848 307574 105904
rect 307630 105848 310040 105904
rect 307569 105846 310040 105848
rect 416773 105904 420164 105906
rect 416773 105848 416778 105904
rect 416834 105848 420164 105904
rect 416773 105846 420164 105848
rect 307569 105843 307635 105846
rect 416773 105843 416839 105846
rect 214005 105768 217242 105770
rect 214005 105712 214010 105768
rect 214066 105712 217242 105768
rect 214005 105710 217242 105712
rect 214005 105707 214071 105710
rect 252277 105634 252343 105637
rect 248952 105632 252343 105634
rect 214097 105226 214163 105229
rect 217182 105226 217242 105604
rect 248952 105576 252282 105632
rect 252338 105576 252343 105632
rect 248952 105574 252343 105576
rect 252277 105571 252343 105574
rect 306741 105498 306807 105501
rect 324313 105498 324379 105501
rect 306741 105496 310040 105498
rect 306741 105440 306746 105496
rect 306802 105440 310040 105496
rect 306741 105438 310040 105440
rect 321908 105496 324379 105498
rect 321908 105440 324318 105496
rect 324374 105440 324379 105496
rect 321908 105438 324379 105440
rect 306741 105435 306807 105438
rect 324313 105435 324379 105438
rect 214097 105224 217242 105226
rect 214097 105168 214102 105224
rect 214158 105168 217242 105224
rect 214097 105166 217242 105168
rect 214097 105163 214163 105166
rect 213913 105090 213979 105093
rect 252001 105090 252067 105093
rect 213913 105088 217242 105090
rect 213913 105032 213918 105088
rect 213974 105032 217242 105088
rect 213913 105030 217242 105032
rect 248952 105088 252067 105090
rect 248952 105032 252006 105088
rect 252062 105032 252067 105088
rect 248952 105030 252067 105032
rect 213913 105027 213979 105030
rect 217182 104924 217242 105030
rect 252001 105027 252067 105030
rect 307661 105090 307727 105093
rect 307661 105088 310040 105090
rect 307661 105032 307666 105088
rect 307722 105032 310040 105088
rect 307661 105030 310040 105032
rect 307661 105027 307727 105030
rect 495433 104954 495499 104957
rect 494316 104952 495499 104954
rect 494316 104896 495438 104952
rect 495494 104896 495499 104952
rect 494316 104894 495499 104896
rect 495433 104891 495499 104894
rect 323025 104818 323091 104821
rect 321908 104816 323091 104818
rect 321908 104760 323030 104816
rect 323086 104760 323091 104816
rect 321908 104758 323091 104760
rect 323025 104755 323091 104758
rect 252277 104682 252343 104685
rect 248952 104680 252343 104682
rect 248952 104624 252282 104680
rect 252338 104624 252343 104680
rect 248952 104622 252343 104624
rect 252277 104619 252343 104622
rect 307477 104682 307543 104685
rect 307477 104680 310040 104682
rect 307477 104624 307482 104680
rect 307538 104624 310040 104680
rect 307477 104622 310040 104624
rect 307477 104619 307543 104622
rect 321737 104546 321803 104549
rect 321694 104544 321803 104546
rect 321694 104488 321742 104544
rect 321798 104488 321803 104544
rect 321694 104483 321803 104488
rect 306925 104274 306991 104277
rect 306925 104272 310040 104274
rect 213913 103866 213979 103869
rect 217182 103866 217242 104244
rect 306925 104216 306930 104272
rect 306986 104216 310040 104272
rect 306925 104214 310040 104216
rect 306925 104211 306991 104214
rect 252369 104138 252435 104141
rect 248952 104136 252435 104138
rect 248952 104080 252374 104136
rect 252430 104080 252435 104136
rect 248952 104078 252435 104080
rect 252369 104075 252435 104078
rect 321694 103972 321754 104483
rect 416773 104138 416839 104141
rect 416773 104136 420164 104138
rect 416773 104080 416778 104136
rect 416834 104080 420164 104136
rect 416773 104078 420164 104080
rect 416773 104075 416839 104078
rect 213913 103864 217242 103866
rect 213913 103808 213918 103864
rect 213974 103808 217242 103864
rect 213913 103806 217242 103808
rect 306741 103866 306807 103869
rect 496905 103866 496971 103869
rect 306741 103864 310040 103866
rect 306741 103808 306746 103864
rect 306802 103808 310040 103864
rect 306741 103806 310040 103808
rect 494316 103864 496971 103866
rect 494316 103808 496910 103864
rect 496966 103808 496971 103864
rect 494316 103806 496971 103808
rect 213913 103803 213979 103806
rect 306741 103803 306807 103806
rect 496905 103803 496971 103806
rect 252461 103730 252527 103733
rect 200070 103670 217242 103730
rect 248952 103728 252527 103730
rect 248952 103672 252466 103728
rect 252522 103672 252527 103728
rect 248952 103670 252527 103672
rect 172094 103532 172100 103596
rect 172164 103594 172170 103596
rect 200070 103594 200130 103670
rect 172164 103534 200130 103594
rect 217182 103564 217242 103670
rect 252461 103667 252527 103670
rect 172164 103532 172170 103534
rect 307569 103458 307635 103461
rect 307569 103456 310040 103458
rect 307569 103400 307574 103456
rect 307630 103400 310040 103456
rect 307569 103398 310040 103400
rect 307569 103395 307635 103398
rect 252461 103186 252527 103189
rect 248952 103184 252527 103186
rect 248952 103128 252466 103184
rect 252522 103128 252527 103184
rect 248952 103126 252527 103128
rect 252461 103123 252527 103126
rect 307661 103050 307727 103053
rect 307661 103048 310040 103050
rect 307661 102992 307666 103048
rect 307722 102992 310040 103048
rect 307661 102990 310040 102992
rect 307661 102987 307727 102990
rect 213913 102642 213979 102645
rect 217182 102642 217242 102884
rect 321878 102781 321938 103156
rect 251817 102778 251883 102781
rect 248952 102776 251883 102778
rect 248952 102720 251822 102776
rect 251878 102720 251883 102776
rect 248952 102718 251883 102720
rect 321878 102776 321987 102781
rect 495433 102778 495499 102781
rect 321878 102720 321926 102776
rect 321982 102720 321987 102776
rect 321878 102718 321987 102720
rect 494316 102776 495499 102778
rect 494316 102720 495438 102776
rect 495494 102720 495499 102776
rect 494316 102718 495499 102720
rect 251817 102715 251883 102718
rect 321921 102715 321987 102718
rect 495433 102715 495499 102718
rect 213913 102640 217242 102642
rect 213913 102584 213918 102640
rect 213974 102584 217242 102640
rect 213913 102582 217242 102584
rect 213913 102579 213979 102582
rect 214414 102444 214420 102508
rect 214484 102506 214490 102508
rect 306557 102506 306623 102509
rect 416773 102506 416839 102509
rect 214484 102446 217426 102506
rect 214484 102444 214490 102446
rect 65977 102370 66043 102373
rect 68142 102370 68816 102376
rect 65977 102368 68816 102370
rect 65977 102312 65982 102368
rect 66038 102316 68816 102368
rect 66038 102312 68202 102316
rect 65977 102310 68202 102312
rect 65977 102307 66043 102310
rect 217366 102204 217426 102446
rect 306557 102504 310040 102506
rect 306557 102448 306562 102504
rect 306618 102448 310040 102504
rect 416773 102504 420164 102506
rect 306557 102446 310040 102448
rect 306557 102443 306623 102446
rect 321694 102237 321754 102476
rect 416773 102448 416778 102504
rect 416834 102448 420164 102504
rect 416773 102446 420164 102448
rect 416773 102443 416839 102446
rect 252369 102234 252435 102237
rect 248952 102232 252435 102234
rect 248952 102176 252374 102232
rect 252430 102176 252435 102232
rect 248952 102174 252435 102176
rect 321694 102232 321803 102237
rect 321694 102176 321742 102232
rect 321798 102176 321803 102232
rect 321694 102174 321803 102176
rect 252369 102171 252435 102174
rect 321737 102171 321803 102174
rect 306557 102098 306623 102101
rect 306557 102096 310040 102098
rect 306557 102040 306562 102096
rect 306618 102040 310040 102096
rect 306557 102038 310040 102040
rect 306557 102035 306623 102038
rect 252461 101826 252527 101829
rect 248952 101824 252527 101826
rect 248952 101768 252466 101824
rect 252522 101768 252527 101824
rect 248952 101766 252527 101768
rect 252461 101763 252527 101766
rect 309133 101826 309199 101829
rect 309726 101826 309732 101828
rect 309133 101824 309732 101826
rect 309133 101768 309138 101824
rect 309194 101768 309732 101824
rect 309133 101766 309732 101768
rect 309133 101763 309199 101766
rect 309726 101764 309732 101766
rect 309796 101764 309802 101828
rect 307477 101690 307543 101693
rect 498377 101690 498443 101693
rect 307477 101688 310040 101690
rect 307477 101632 307482 101688
rect 307538 101632 310040 101688
rect 494316 101688 498443 101690
rect 307477 101630 310040 101632
rect 307477 101627 307543 101630
rect 169150 101356 169156 101420
rect 169220 101418 169226 101420
rect 214557 101418 214623 101421
rect 169220 101416 214623 101418
rect 169220 101360 214562 101416
rect 214618 101360 214623 101416
rect 169220 101358 214623 101360
rect 169220 101356 169226 101358
rect 214557 101355 214623 101358
rect 214833 101146 214899 101149
rect 217182 101146 217242 101524
rect 251725 101418 251791 101421
rect 248952 101416 251791 101418
rect 248952 101360 251730 101416
rect 251786 101360 251791 101416
rect 248952 101358 251791 101360
rect 251725 101355 251791 101358
rect 307569 101282 307635 101285
rect 307569 101280 310040 101282
rect 307569 101224 307574 101280
rect 307630 101224 310040 101280
rect 307569 101222 310040 101224
rect 307569 101219 307635 101222
rect 321694 101149 321754 101660
rect 494316 101632 498382 101688
rect 498438 101632 498443 101688
rect 494316 101630 498443 101632
rect 498377 101627 498443 101630
rect 214833 101144 217242 101146
rect 214833 101088 214838 101144
rect 214894 101088 217242 101144
rect 214833 101086 217242 101088
rect 321645 101144 321754 101149
rect 321645 101088 321650 101144
rect 321706 101088 321754 101144
rect 321645 101086 321754 101088
rect 214833 101083 214899 101086
rect 321645 101083 321711 101086
rect 213913 100874 213979 100877
rect 213913 100872 216874 100874
rect 213913 100816 213918 100872
rect 213974 100816 216874 100872
rect 213913 100814 216874 100816
rect 213913 100811 213979 100814
rect 67725 100738 67791 100741
rect 68142 100738 68816 100744
rect 67725 100736 68816 100738
rect 67725 100680 67730 100736
rect 67786 100684 68816 100736
rect 216814 100738 216874 100814
rect 217366 100738 217426 100980
rect 252369 100874 252435 100877
rect 248952 100872 252435 100874
rect 248952 100816 252374 100872
rect 252430 100816 252435 100872
rect 248952 100814 252435 100816
rect 252369 100811 252435 100814
rect 307661 100874 307727 100877
rect 324405 100874 324471 100877
rect 307661 100872 310040 100874
rect 307661 100816 307666 100872
rect 307722 100816 310040 100872
rect 307661 100814 310040 100816
rect 321908 100872 324471 100874
rect 321908 100816 324410 100872
rect 324466 100816 324471 100872
rect 321908 100814 324471 100816
rect 307661 100811 307727 100814
rect 324405 100811 324471 100814
rect 416773 100874 416839 100877
rect 416773 100872 420164 100874
rect 416773 100816 416778 100872
rect 416834 100816 420164 100872
rect 416773 100814 420164 100816
rect 416773 100811 416839 100814
rect 67786 100680 68202 100684
rect 67725 100678 68202 100680
rect 216814 100678 217426 100738
rect 67725 100675 67791 100678
rect 252461 100466 252527 100469
rect 248952 100464 252527 100466
rect 248952 100408 252466 100464
rect 252522 100408 252527 100464
rect 248952 100406 252527 100408
rect 252461 100403 252527 100406
rect 307477 100466 307543 100469
rect 307477 100464 310040 100466
rect 307477 100408 307482 100464
rect 307538 100408 310040 100464
rect 307477 100406 310040 100408
rect 307477 100403 307543 100406
rect 214097 99786 214163 99789
rect 217182 99786 217242 100300
rect 307569 100058 307635 100061
rect 307569 100056 310040 100058
rect 307569 100000 307574 100056
rect 307630 100000 310040 100056
rect 307569 99998 310040 100000
rect 307569 99995 307635 99998
rect 252277 99922 252343 99925
rect 248952 99920 252343 99922
rect 248952 99864 252282 99920
rect 252338 99864 252343 99920
rect 248952 99862 252343 99864
rect 252277 99859 252343 99862
rect 214097 99784 217242 99786
rect 214097 99728 214102 99784
rect 214158 99728 217242 99784
rect 214097 99726 217242 99728
rect 214097 99723 214163 99726
rect 307661 99650 307727 99653
rect 321369 99650 321435 99653
rect 321510 99650 321570 100164
rect 494102 100061 494162 100572
rect 494053 100056 494162 100061
rect 494053 100000 494058 100056
rect 494114 100000 494162 100056
rect 494053 99998 494162 100000
rect 494053 99995 494119 99998
rect 307661 99648 310040 99650
rect 214281 99514 214347 99517
rect 214281 99512 216874 99514
rect 214281 99456 214286 99512
rect 214342 99456 216874 99512
rect 214281 99454 216874 99456
rect 214281 99451 214347 99454
rect 216814 99378 216874 99454
rect 217366 99378 217426 99620
rect 307661 99592 307666 99648
rect 307722 99592 310040 99648
rect 307661 99590 310040 99592
rect 321369 99648 321570 99650
rect 321369 99592 321374 99648
rect 321430 99592 321570 99648
rect 321369 99590 321570 99592
rect 307661 99587 307727 99590
rect 321369 99587 321435 99590
rect 252369 99514 252435 99517
rect 248952 99512 252435 99514
rect 248952 99456 252374 99512
rect 252430 99456 252435 99512
rect 248952 99454 252435 99456
rect 252369 99451 252435 99454
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 324262 99378 324268 99380
rect 216814 99318 217426 99378
rect 321908 99318 324268 99378
rect 324262 99316 324268 99318
rect 324332 99316 324338 99380
rect 583520 99364 584960 99454
rect 307569 99106 307635 99109
rect 307569 99104 310040 99106
rect 307569 99048 307574 99104
rect 307630 99048 310040 99104
rect 307569 99046 310040 99048
rect 307569 99043 307635 99046
rect 252461 98970 252527 98973
rect 248952 98968 252527 98970
rect 214005 98426 214071 98429
rect 217182 98426 217242 98940
rect 248952 98912 252466 98968
rect 252522 98912 252527 98968
rect 248952 98910 252527 98912
rect 252461 98907 252527 98910
rect 307661 98698 307727 98701
rect 307661 98696 310040 98698
rect 307661 98640 307666 98696
rect 307722 98640 310040 98696
rect 307661 98638 310040 98640
rect 307661 98635 307727 98638
rect 252369 98562 252435 98565
rect 248952 98560 252435 98562
rect 248952 98504 252374 98560
rect 252430 98504 252435 98560
rect 248952 98502 252435 98504
rect 252369 98499 252435 98502
rect 214005 98424 217242 98426
rect 214005 98368 214010 98424
rect 214066 98368 217242 98424
rect 214005 98366 217242 98368
rect 214005 98363 214071 98366
rect 307293 98290 307359 98293
rect 307293 98288 310040 98290
rect 213913 98018 213979 98021
rect 217366 98018 217426 98260
rect 307293 98232 307298 98288
rect 307354 98232 310040 98288
rect 307293 98230 310040 98232
rect 307293 98227 307359 98230
rect 251357 98018 251423 98021
rect 321510 98020 321570 98532
rect 213913 98016 217426 98018
rect 213913 97960 213918 98016
rect 213974 97960 217426 98016
rect 213913 97958 217426 97960
rect 248952 98016 251423 98018
rect 248952 97960 251362 98016
rect 251418 97960 251423 98016
rect 248952 97958 251423 97960
rect 213913 97955 213979 97958
rect 251357 97955 251423 97958
rect 321502 97956 321508 98020
rect 321572 97956 321578 98020
rect 307201 97882 307267 97885
rect 307201 97880 310040 97882
rect 307201 97824 307206 97880
rect 307262 97824 310040 97880
rect 307201 97822 310040 97824
rect 307201 97819 307267 97822
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect 252185 97610 252251 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect 248952 97608 252251 97610
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 216673 97066 216739 97069
rect 217182 97066 217242 97580
rect 248952 97552 252190 97608
rect 252246 97552 252251 97608
rect 248952 97550 252251 97552
rect 252185 97547 252251 97550
rect 307569 97474 307635 97477
rect 307569 97472 310040 97474
rect 307569 97416 307574 97472
rect 307630 97416 310040 97472
rect 307569 97414 310040 97416
rect 307569 97411 307635 97414
rect 321510 97341 321570 97852
rect 252461 97338 252527 97341
rect 262070 97338 262076 97340
rect 252461 97336 262076 97338
rect 252461 97280 252466 97336
rect 252522 97280 262076 97336
rect 252461 97278 262076 97280
rect 252461 97275 252527 97278
rect 262070 97276 262076 97278
rect 262140 97276 262146 97340
rect 321461 97336 321570 97341
rect 321461 97280 321466 97336
rect 321522 97280 321570 97336
rect 321461 97278 321570 97280
rect 321461 97275 321527 97278
rect 269614 97202 269620 97204
rect 258030 97142 269620 97202
rect 249793 97066 249859 97069
rect 258030 97066 258090 97142
rect 269614 97140 269620 97142
rect 269684 97140 269690 97204
rect 216673 97064 217242 97066
rect 216673 97008 216678 97064
rect 216734 97008 217242 97064
rect 216673 97006 217242 97008
rect 248952 97064 258090 97066
rect 248952 97008 249798 97064
rect 249854 97008 258090 97064
rect 248952 97006 258090 97008
rect 307385 97066 307451 97069
rect 307385 97064 310040 97066
rect 307385 97008 307390 97064
rect 307446 97008 310040 97064
rect 307385 97006 310040 97008
rect 216673 97003 216739 97006
rect 249793 97003 249859 97006
rect 307385 97003 307451 97006
rect 214649 96658 214715 96661
rect 217182 96658 217242 96900
rect 321510 96661 321570 97036
rect 252461 96658 252527 96661
rect 214649 96656 217242 96658
rect 214649 96600 214654 96656
rect 214710 96600 217242 96656
rect 214649 96598 217242 96600
rect 248952 96656 252527 96658
rect 248952 96600 252466 96656
rect 252522 96600 252527 96656
rect 248952 96598 252527 96600
rect 214649 96595 214715 96598
rect 252461 96595 252527 96598
rect 307661 96658 307727 96661
rect 307661 96656 310040 96658
rect 307661 96600 307666 96656
rect 307722 96600 310040 96656
rect 307661 96598 310040 96600
rect 321510 96656 321619 96661
rect 321510 96600 321558 96656
rect 321614 96600 321619 96656
rect 321510 96598 321619 96600
rect 307661 96595 307727 96598
rect 321553 96595 321619 96598
rect 214557 95842 214623 95845
rect 217182 95842 217242 96356
rect 251173 96250 251239 96253
rect 248860 96248 251239 96250
rect 248860 96192 251178 96248
rect 251234 96192 251239 96248
rect 248860 96190 251239 96192
rect 251173 96187 251239 96190
rect 307661 96250 307727 96253
rect 307661 96248 310132 96250
rect 307661 96192 307666 96248
rect 307722 96192 310132 96248
rect 307661 96190 310132 96192
rect 307661 96187 307727 96190
rect 214557 95840 217242 95842
rect 214557 95784 214562 95840
rect 214618 95784 217242 95840
rect 214557 95782 217242 95784
rect 214557 95779 214623 95782
rect 173198 95508 173204 95572
rect 173268 95570 173274 95572
rect 321326 95570 321386 96356
rect 173268 95510 321386 95570
rect 173268 95508 173274 95510
rect 67357 94890 67423 94893
rect 206553 94890 206619 94893
rect 67357 94888 206619 94890
rect 67357 94832 67362 94888
rect 67418 94832 206558 94888
rect 206614 94832 206619 94888
rect 67357 94830 206619 94832
rect 67357 94827 67423 94830
rect 206553 94827 206619 94830
rect 66069 94754 66135 94757
rect 173433 94754 173499 94757
rect 66069 94752 173499 94754
rect 66069 94696 66074 94752
rect 66130 94696 173438 94752
rect 173494 94696 173499 94752
rect 66069 94694 173499 94696
rect 66069 94691 66135 94694
rect 173433 94691 173499 94694
rect 151486 94556 151492 94620
rect 151556 94618 151562 94620
rect 151760 94618 151766 94620
rect 151556 94558 151766 94618
rect 151556 94556 151562 94558
rect 151760 94556 151766 94558
rect 151830 94556 151836 94620
rect 246481 94482 246547 94485
rect 255814 94482 255820 94484
rect 246481 94480 255820 94482
rect 246481 94424 246486 94480
rect 246542 94424 255820 94480
rect 246481 94422 255820 94424
rect 246481 94419 246547 94422
rect 255814 94420 255820 94422
rect 255884 94420 255890 94484
rect 126513 94212 126579 94213
rect 152089 94212 152155 94213
rect 126462 94148 126468 94212
rect 126532 94210 126579 94212
rect 126532 94208 126624 94210
rect 126574 94152 126624 94208
rect 126532 94150 126624 94152
rect 126532 94148 126579 94150
rect 152038 94148 152044 94212
rect 152108 94210 152155 94212
rect 152108 94208 152200 94210
rect 152150 94152 152200 94208
rect 152108 94150 152200 94152
rect 152108 94148 152155 94150
rect 126513 94147 126579 94148
rect 152089 94147 152155 94148
rect 112345 94076 112411 94077
rect 126697 94076 126763 94077
rect 112294 94012 112300 94076
rect 112364 94074 112411 94076
rect 112364 94072 112456 94074
rect 112406 94016 112456 94072
rect 112364 94014 112456 94016
rect 112364 94012 112411 94014
rect 126646 94012 126652 94076
rect 126716 94074 126763 94076
rect 126716 94072 126808 94074
rect 126758 94016 126808 94072
rect 126716 94014 126808 94016
rect 126716 94012 126763 94014
rect 112345 94011 112411 94012
rect 126697 94011 126763 94012
rect 96153 93940 96219 93941
rect 96102 93876 96108 93940
rect 96172 93938 96219 93940
rect 96172 93936 96264 93938
rect 96214 93880 96264 93936
rect 96172 93878 96264 93880
rect 96172 93876 96219 93878
rect 96153 93875 96219 93876
rect 4061 93802 4127 93805
rect 495709 93802 495775 93805
rect 4061 93800 495775 93802
rect 4061 93744 4066 93800
rect 4122 93744 495714 93800
rect 495770 93744 495775 93800
rect 4061 93742 495775 93744
rect 4061 93739 4127 93742
rect 495709 93739 495775 93742
rect 59261 93666 59327 93669
rect 203609 93666 203675 93669
rect 59261 93664 203675 93666
rect 59261 93608 59266 93664
rect 59322 93608 203614 93664
rect 203670 93608 203675 93664
rect 59261 93606 203675 93608
rect 59261 93603 59327 93606
rect 203609 93603 203675 93606
rect 100937 93532 101003 93533
rect 109217 93532 109283 93533
rect 116761 93532 116827 93533
rect 121729 93532 121795 93533
rect 133137 93532 133203 93533
rect 151721 93532 151787 93533
rect 100886 93530 100892 93532
rect 100846 93470 100892 93530
rect 100956 93528 101003 93532
rect 109166 93530 109172 93532
rect 100998 93472 101003 93528
rect 100886 93468 100892 93470
rect 100956 93468 101003 93472
rect 109126 93470 109172 93530
rect 109236 93528 109283 93532
rect 116710 93530 116716 93532
rect 109278 93472 109283 93528
rect 109166 93468 109172 93470
rect 109236 93468 109283 93472
rect 116670 93470 116716 93530
rect 116780 93528 116827 93532
rect 121678 93530 121684 93532
rect 116822 93472 116827 93528
rect 116710 93468 116716 93470
rect 116780 93468 116827 93472
rect 121638 93470 121684 93530
rect 121748 93528 121795 93532
rect 133086 93530 133092 93532
rect 121790 93472 121795 93528
rect 121678 93468 121684 93470
rect 121748 93468 121795 93472
rect 133046 93470 133092 93530
rect 133156 93528 133203 93532
rect 151670 93530 151676 93532
rect 133198 93472 133203 93528
rect 133086 93468 133092 93470
rect 133156 93468 133203 93472
rect 151630 93470 151676 93530
rect 151740 93528 151787 93532
rect 151782 93472 151787 93528
rect 151670 93468 151676 93470
rect 151740 93468 151787 93472
rect 100937 93467 101003 93468
rect 109217 93467 109283 93468
rect 116761 93467 116827 93468
rect 121729 93467 121795 93468
rect 133137 93467 133203 93468
rect 151721 93467 151787 93468
rect 188429 93530 188495 93533
rect 324262 93530 324268 93532
rect 188429 93528 324268 93530
rect 188429 93472 188434 93528
rect 188490 93472 324268 93528
rect 188429 93470 324268 93472
rect 188429 93467 188495 93470
rect 324262 93468 324268 93470
rect 324332 93468 324338 93532
rect 103329 93260 103395 93261
rect 110137 93260 110203 93261
rect 103278 93258 103284 93260
rect 103238 93198 103284 93258
rect 103348 93256 103395 93260
rect 110086 93258 110092 93260
rect 103390 93200 103395 93256
rect 103278 93196 103284 93198
rect 103348 93196 103395 93200
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 103329 93195 103395 93196
rect 110137 93195 110203 93196
rect 74809 92444 74875 92445
rect 85849 92444 85915 92445
rect 88057 92444 88123 92445
rect 88977 92444 89043 92445
rect 74758 92442 74764 92444
rect 74718 92382 74764 92442
rect 74828 92440 74875 92444
rect 85798 92442 85804 92444
rect 74870 92384 74875 92440
rect 74758 92380 74764 92382
rect 74828 92380 74875 92384
rect 85758 92382 85804 92442
rect 85868 92440 85915 92444
rect 88006 92442 88012 92444
rect 85910 92384 85915 92440
rect 85798 92380 85804 92382
rect 85868 92380 85915 92384
rect 87966 92382 88012 92442
rect 88076 92440 88123 92444
rect 88926 92442 88932 92444
rect 88118 92384 88123 92440
rect 88006 92380 88012 92382
rect 88076 92380 88123 92384
rect 88886 92382 88932 92442
rect 88996 92440 89043 92444
rect 89038 92384 89043 92440
rect 88926 92380 88932 92382
rect 88996 92380 89043 92384
rect 97206 92380 97212 92444
rect 97276 92442 97282 92444
rect 97533 92442 97599 92445
rect 97276 92440 97599 92442
rect 97276 92384 97538 92440
rect 97594 92384 97599 92440
rect 97276 92382 97599 92384
rect 97276 92380 97282 92382
rect 74809 92379 74875 92380
rect 85849 92379 85915 92380
rect 88057 92379 88123 92380
rect 88977 92379 89043 92380
rect 97533 92379 97599 92382
rect 98494 92380 98500 92444
rect 98564 92442 98570 92444
rect 98821 92442 98887 92445
rect 98564 92440 98887 92442
rect 98564 92384 98826 92440
rect 98882 92384 98887 92440
rect 98564 92382 98887 92384
rect 98564 92380 98570 92382
rect 98821 92379 98887 92382
rect 113030 92380 113036 92444
rect 113100 92442 113106 92444
rect 114461 92442 114527 92445
rect 114921 92444 114987 92445
rect 115473 92444 115539 92445
rect 118049 92444 118115 92445
rect 132401 92444 132467 92445
rect 151537 92444 151603 92445
rect 114870 92442 114876 92444
rect 113100 92440 114527 92442
rect 113100 92384 114466 92440
rect 114522 92384 114527 92440
rect 113100 92382 114527 92384
rect 114830 92382 114876 92442
rect 114940 92440 114987 92444
rect 115422 92442 115428 92444
rect 114982 92384 114987 92440
rect 113100 92380 113106 92382
rect 114461 92379 114527 92382
rect 114870 92380 114876 92382
rect 114940 92380 114987 92384
rect 115382 92382 115428 92442
rect 115492 92440 115539 92444
rect 117998 92442 118004 92444
rect 115534 92384 115539 92440
rect 115422 92380 115428 92382
rect 115492 92380 115539 92384
rect 117958 92382 118004 92442
rect 118068 92440 118115 92444
rect 132350 92442 132356 92444
rect 118110 92384 118115 92440
rect 117998 92380 118004 92382
rect 118068 92380 118115 92384
rect 132310 92382 132356 92442
rect 132420 92440 132467 92444
rect 151486 92442 151492 92444
rect 132462 92384 132467 92440
rect 132350 92380 132356 92382
rect 132420 92380 132467 92384
rect 151446 92382 151492 92442
rect 151556 92440 151603 92444
rect 151598 92384 151603 92440
rect 151486 92380 151492 92382
rect 151556 92380 151603 92384
rect 114921 92379 114987 92380
rect 115473 92379 115539 92380
rect 118049 92379 118115 92380
rect 132401 92379 132467 92380
rect 151537 92379 151603 92380
rect 102726 92244 102732 92308
rect 102796 92306 102802 92308
rect 103237 92306 103303 92309
rect 102796 92304 103303 92306
rect 102796 92248 103242 92304
rect 103298 92248 103303 92304
rect 102796 92246 103303 92248
rect 102796 92244 102802 92246
rect 103237 92243 103303 92246
rect 122046 92244 122052 92308
rect 122116 92306 122122 92308
rect 169150 92306 169156 92308
rect 122116 92246 169156 92306
rect 122116 92244 122122 92246
rect 169150 92244 169156 92246
rect 169220 92244 169226 92308
rect 122833 92172 122899 92173
rect 122782 92108 122788 92172
rect 122852 92170 122899 92172
rect 122852 92168 122944 92170
rect 122894 92112 122944 92168
rect 122852 92110 122944 92112
rect 122852 92108 122899 92110
rect 151302 92108 151308 92172
rect 151372 92170 151378 92172
rect 151629 92170 151695 92173
rect 151372 92168 151695 92170
rect 151372 92112 151634 92168
rect 151690 92112 151695 92168
rect 151372 92110 151695 92112
rect 151372 92108 151378 92110
rect 122833 92107 122899 92108
rect 151629 92107 151695 92110
rect 90214 91700 90220 91764
rect 90284 91762 90290 91764
rect 90725 91762 90791 91765
rect 90284 91760 90791 91762
rect 90284 91704 90730 91760
rect 90786 91704 90791 91760
rect 90284 91702 90791 91704
rect 90284 91700 90290 91702
rect 90725 91699 90791 91702
rect 119286 91564 119292 91628
rect 119356 91626 119362 91628
rect 119797 91626 119863 91629
rect 119356 91624 119863 91626
rect 119356 91568 119802 91624
rect 119858 91568 119863 91624
rect 119356 91566 119863 91568
rect 119356 91564 119362 91566
rect 119797 91563 119863 91566
rect 136030 91564 136036 91628
rect 136100 91626 136106 91628
rect 136449 91626 136515 91629
rect 136100 91624 136515 91626
rect 136100 91568 136454 91624
rect 136510 91568 136515 91624
rect 136100 91566 136515 91568
rect 136100 91564 136106 91566
rect 136449 91563 136515 91566
rect 93894 91292 93900 91356
rect 93964 91354 93970 91356
rect 95049 91354 95115 91357
rect 93964 91352 95115 91354
rect 93964 91296 95054 91352
rect 95110 91296 95115 91352
rect 93964 91294 95115 91296
rect 93964 91292 93970 91294
rect 95049 91291 95115 91294
rect 98126 91292 98132 91356
rect 98196 91354 98202 91356
rect 99189 91354 99255 91357
rect 100569 91356 100635 91357
rect 101857 91356 101923 91357
rect 100518 91354 100524 91356
rect 98196 91352 99255 91354
rect 98196 91296 99194 91352
rect 99250 91296 99255 91352
rect 98196 91294 99255 91296
rect 100478 91294 100524 91354
rect 100588 91352 100635 91356
rect 101806 91354 101812 91356
rect 100630 91296 100635 91352
rect 98196 91292 98202 91294
rect 99189 91291 99255 91294
rect 100518 91292 100524 91294
rect 100588 91292 100635 91296
rect 101766 91294 101812 91354
rect 101876 91352 101923 91356
rect 101918 91296 101923 91352
rect 101806 91292 101812 91294
rect 101876 91292 101923 91296
rect 105486 91292 105492 91356
rect 105556 91354 105562 91356
rect 106089 91354 106155 91357
rect 105556 91352 106155 91354
rect 105556 91296 106094 91352
rect 106150 91296 106155 91352
rect 105556 91294 106155 91296
rect 105556 91292 105562 91294
rect 100569 91291 100635 91292
rect 101857 91291 101923 91292
rect 106089 91291 106155 91294
rect 106406 91292 106412 91356
rect 106476 91354 106482 91356
rect 107561 91354 107627 91357
rect 106476 91352 107627 91354
rect 106476 91296 107566 91352
rect 107622 91296 107627 91352
rect 106476 91294 107627 91296
rect 106476 91292 106482 91294
rect 107561 91291 107627 91294
rect 120574 91292 120580 91356
rect 120644 91354 120650 91356
rect 120717 91354 120783 91357
rect 120644 91352 120783 91354
rect 120644 91296 120722 91352
rect 120778 91296 120783 91352
rect 120644 91294 120783 91296
rect 120644 91292 120650 91294
rect 120717 91291 120783 91294
rect 124029 91356 124095 91357
rect 124029 91352 124076 91356
rect 124140 91354 124146 91356
rect 124029 91296 124034 91352
rect 124029 91292 124076 91296
rect 124140 91294 124186 91354
rect 124140 91292 124146 91294
rect 124438 91292 124444 91356
rect 124508 91354 124514 91356
rect 125409 91354 125475 91357
rect 124508 91352 125475 91354
rect 124508 91296 125414 91352
rect 125470 91296 125475 91352
rect 124508 91294 125475 91296
rect 124508 91292 124514 91294
rect 124029 91291 124095 91292
rect 125409 91291 125475 91294
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85481 91218 85547 91221
rect 86769 91220 86835 91221
rect 86718 91218 86724 91220
rect 84396 91216 85547 91218
rect 84396 91160 85486 91216
rect 85542 91160 85547 91216
rect 84396 91158 85547 91160
rect 86678 91158 86724 91218
rect 86788 91216 86835 91220
rect 86830 91160 86835 91216
rect 84396 91156 84402 91158
rect 85481 91155 85547 91158
rect 86718 91156 86724 91158
rect 86788 91156 86835 91160
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92381 91218 92447 91221
rect 91388 91216 92447 91218
rect 91388 91160 92386 91216
rect 92442 91160 92447 91216
rect 91388 91158 92447 91160
rect 91388 91156 91394 91158
rect 86769 91155 86835 91156
rect 92381 91155 92447 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96654 91156 96660 91220
rect 96724 91218 96730 91220
rect 97809 91218 97875 91221
rect 96724 91216 97875 91218
rect 96724 91160 97814 91216
rect 97870 91160 97875 91216
rect 96724 91158 97875 91160
rect 96724 91156 96730 91158
rect 97809 91155 97875 91158
rect 99046 91156 99052 91220
rect 99116 91218 99122 91220
rect 99281 91218 99347 91221
rect 99116 91216 99347 91218
rect 99116 91160 99286 91216
rect 99342 91160 99347 91216
rect 99116 91158 99347 91160
rect 99116 91156 99122 91158
rect 99281 91155 99347 91158
rect 99966 91156 99972 91220
rect 100036 91218 100042 91220
rect 100661 91218 100727 91221
rect 102041 91220 102107 91221
rect 104249 91220 104315 91221
rect 101990 91218 101996 91220
rect 100036 91216 100727 91218
rect 100036 91160 100666 91216
rect 100722 91160 100727 91216
rect 100036 91158 100727 91160
rect 101950 91158 101996 91218
rect 102060 91216 102107 91220
rect 104198 91218 104204 91220
rect 102102 91160 102107 91216
rect 100036 91156 100042 91158
rect 100661 91155 100727 91158
rect 101990 91156 101996 91158
rect 102060 91156 102107 91160
rect 104158 91158 104204 91218
rect 104268 91216 104315 91220
rect 104310 91160 104315 91216
rect 104198 91156 104204 91158
rect 104268 91156 104315 91160
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104801 91218 104867 91221
rect 104636 91216 104867 91218
rect 104636 91160 104806 91216
rect 104862 91160 104867 91216
rect 104636 91158 104867 91160
rect 104636 91156 104642 91158
rect 102041 91155 102107 91156
rect 104249 91155 104315 91156
rect 104801 91155 104867 91158
rect 105670 91156 105676 91220
rect 105740 91218 105746 91220
rect 106181 91218 106247 91221
rect 105740 91216 106247 91218
rect 105740 91160 106186 91216
rect 106242 91160 106247 91216
rect 105740 91158 106247 91160
rect 105740 91156 105746 91158
rect 106181 91155 106247 91158
rect 106774 91156 106780 91220
rect 106844 91218 106850 91220
rect 107469 91218 107535 91221
rect 106844 91216 107535 91218
rect 106844 91160 107474 91216
rect 107530 91160 107535 91216
rect 106844 91158 107535 91160
rect 106844 91156 106850 91158
rect 107469 91155 107535 91158
rect 107694 91156 107700 91220
rect 107764 91218 107770 91220
rect 107929 91218 107995 91221
rect 107764 91216 107995 91218
rect 107764 91160 107934 91216
rect 107990 91160 107995 91216
rect 107764 91158 107995 91160
rect 107764 91156 107770 91158
rect 107929 91155 107995 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108941 91218 109007 91221
rect 108132 91216 109007 91218
rect 108132 91160 108946 91216
rect 109002 91160 109007 91216
rect 108132 91158 109007 91160
rect 108132 91156 108138 91158
rect 108941 91155 109007 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110321 91218 110387 91221
rect 110689 91220 110755 91221
rect 110638 91218 110644 91220
rect 109604 91216 110387 91218
rect 109604 91160 110326 91216
rect 110382 91160 110387 91216
rect 109604 91158 110387 91160
rect 110598 91158 110644 91218
rect 110708 91216 110755 91220
rect 110750 91160 110755 91216
rect 109604 91156 109610 91158
rect 110321 91155 110387 91158
rect 110638 91156 110644 91158
rect 110708 91156 110755 91160
rect 111190 91156 111196 91220
rect 111260 91218 111266 91220
rect 111701 91218 111767 91221
rect 111260 91216 111767 91218
rect 111260 91160 111706 91216
rect 111762 91160 111767 91216
rect 111260 91158 111767 91160
rect 111260 91156 111266 91158
rect 110689 91155 110755 91156
rect 111701 91155 111767 91158
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 113081 91218 113147 91221
rect 111996 91216 113147 91218
rect 111996 91160 113086 91216
rect 113142 91160 113147 91216
rect 111996 91158 113147 91160
rect 111996 91156 112002 91158
rect 113081 91155 113147 91158
rect 113214 91156 113220 91220
rect 113284 91218 113290 91220
rect 113357 91218 113423 91221
rect 114369 91220 114435 91221
rect 114318 91218 114324 91220
rect 113284 91216 113423 91218
rect 113284 91160 113362 91216
rect 113418 91160 113423 91216
rect 113284 91158 113423 91160
rect 114278 91158 114324 91218
rect 114388 91216 114435 91220
rect 115749 91220 115815 91221
rect 117129 91220 117195 91221
rect 115749 91218 115796 91220
rect 114430 91160 114435 91216
rect 113284 91156 113290 91158
rect 113357 91155 113423 91158
rect 114318 91156 114324 91158
rect 114388 91156 114435 91160
rect 115704 91216 115796 91218
rect 115704 91160 115754 91216
rect 115704 91158 115796 91160
rect 114369 91155 114435 91156
rect 115749 91156 115796 91158
rect 115860 91156 115866 91220
rect 117078 91218 117084 91220
rect 117038 91158 117084 91218
rect 117148 91216 117195 91220
rect 117190 91160 117195 91216
rect 117078 91156 117084 91158
rect 117148 91156 117195 91160
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118601 91218 118667 91221
rect 118252 91216 118667 91218
rect 118252 91160 118606 91216
rect 118662 91160 118667 91216
rect 118252 91158 118667 91160
rect 118252 91156 118258 91158
rect 115749 91155 115815 91156
rect 117129 91155 117195 91156
rect 118601 91155 118667 91158
rect 119654 91156 119660 91220
rect 119724 91218 119730 91220
rect 119981 91218 120047 91221
rect 119724 91216 120047 91218
rect 119724 91160 119986 91216
rect 120042 91160 120047 91216
rect 119724 91158 120047 91160
rect 119724 91156 119730 91158
rect 119981 91155 120047 91158
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 121361 91218 121427 91221
rect 120276 91216 121427 91218
rect 120276 91160 121366 91216
rect 121422 91160 121427 91216
rect 120276 91158 121427 91160
rect 120276 91156 120282 91158
rect 121361 91155 121427 91158
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 124121 91218 124187 91221
rect 123220 91216 124187 91218
rect 123220 91160 124126 91216
rect 124182 91160 124187 91216
rect 123220 91158 124187 91160
rect 123220 91156 123226 91158
rect 124121 91155 124187 91158
rect 125358 91156 125364 91220
rect 125428 91218 125434 91220
rect 125501 91218 125567 91221
rect 125428 91216 125567 91218
rect 125428 91160 125506 91216
rect 125562 91160 125567 91216
rect 125428 91158 125567 91160
rect 125428 91156 125434 91158
rect 125501 91155 125567 91158
rect 125726 91156 125732 91220
rect 125796 91218 125802 91220
rect 126513 91218 126579 91221
rect 129457 91220 129523 91221
rect 130745 91220 130811 91221
rect 129406 91218 129412 91220
rect 125796 91216 126579 91218
rect 125796 91160 126518 91216
rect 126574 91160 126579 91216
rect 125796 91158 126579 91160
rect 129366 91158 129412 91218
rect 129476 91216 129523 91220
rect 130694 91218 130700 91220
rect 129518 91160 129523 91216
rect 125796 91156 125802 91158
rect 126513 91155 126579 91158
rect 129406 91156 129412 91158
rect 129476 91156 129523 91160
rect 130654 91158 130700 91218
rect 130764 91216 130811 91220
rect 130806 91160 130811 91216
rect 130694 91156 130700 91158
rect 130764 91156 130811 91160
rect 134374 91156 134380 91220
rect 134444 91218 134450 91220
rect 135161 91218 135227 91221
rect 134444 91216 135227 91218
rect 134444 91160 135166 91216
rect 135222 91160 135227 91216
rect 134444 91158 135227 91160
rect 134444 91156 134450 91158
rect 129457 91155 129523 91156
rect 130745 91155 130811 91156
rect 135161 91155 135227 91158
rect 67449 91082 67515 91085
rect 214414 91082 214420 91084
rect 67449 91080 214420 91082
rect 67449 91024 67454 91080
rect 67510 91024 214420 91080
rect 67449 91022 214420 91024
rect 67449 91019 67515 91022
rect 214414 91020 214420 91022
rect 214484 91020 214490 91084
rect 127566 90884 127572 90948
rect 127636 90946 127642 90948
rect 170489 90946 170555 90949
rect 127636 90944 170555 90946
rect 127636 90888 170494 90944
rect 170550 90888 170555 90944
rect 127636 90886 170555 90888
rect 127636 90884 127642 90886
rect 170489 90883 170555 90886
rect 202229 90402 202295 90405
rect 307150 90402 307156 90404
rect 202229 90400 307156 90402
rect 202229 90344 202234 90400
rect 202290 90344 307156 90400
rect 202229 90342 307156 90344
rect 202229 90339 202295 90342
rect 307150 90340 307156 90342
rect 307220 90340 307226 90404
rect 310094 90340 310100 90404
rect 310164 90402 310170 90404
rect 311893 90402 311959 90405
rect 310164 90400 311959 90402
rect 310164 90344 311898 90400
rect 311954 90344 311959 90400
rect 310164 90342 311959 90344
rect 310164 90340 310170 90342
rect 311893 90339 311959 90342
rect 67541 89722 67607 89725
rect 209221 89722 209287 89725
rect 67541 89720 209287 89722
rect 67541 89664 67546 89720
rect 67602 89664 209226 89720
rect 209282 89664 209287 89720
rect 67541 89662 209287 89664
rect 67541 89659 67607 89662
rect 209221 89659 209287 89662
rect 110689 88226 110755 88229
rect 170438 88226 170444 88228
rect 110689 88224 170444 88226
rect 110689 88168 110694 88224
rect 110750 88168 170444 88224
rect 110689 88166 170444 88168
rect 110689 88163 110755 88166
rect 170438 88164 170444 88166
rect 170508 88164 170514 88228
rect 342345 87684 342411 87685
rect 342294 87620 342300 87684
rect 342364 87682 342411 87684
rect 342364 87680 342456 87682
rect 342406 87624 342456 87680
rect 342364 87622 342456 87624
rect 342364 87620 342411 87622
rect 342345 87619 342411 87620
rect 198089 86186 198155 86189
rect 251173 86186 251239 86189
rect 336038 86186 336044 86188
rect 198089 86184 336044 86186
rect 198089 86128 198094 86184
rect 198150 86128 251178 86184
rect 251234 86128 336044 86184
rect 198089 86126 336044 86128
rect 198089 86123 198155 86126
rect 251173 86123 251239 86126
rect 336038 86124 336044 86126
rect 336108 86124 336114 86188
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 130745 85506 130811 85509
rect 168230 85506 168236 85508
rect 130745 85504 168236 85506
rect 130745 85448 130750 85504
rect 130806 85448 168236 85504
rect 130745 85446 168236 85448
rect 130745 85443 130811 85446
rect 168230 85444 168236 85446
rect 168300 85444 168306 85508
rect 170397 84826 170463 84829
rect 306966 84826 306972 84828
rect 170397 84824 306972 84826
rect -960 84690 480 84780
rect 170397 84768 170402 84824
rect 170458 84768 306972 84824
rect 170397 84766 306972 84768
rect 170397 84763 170463 84766
rect 306966 84764 306972 84766
rect 307036 84764 307042 84828
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 66161 84146 66227 84149
rect 172094 84146 172100 84148
rect 66161 84144 172100 84146
rect 66161 84088 66166 84144
rect 66222 84088 172100 84144
rect 66161 84086 172100 84088
rect 66161 84083 66227 84086
rect 172094 84084 172100 84086
rect 172164 84084 172170 84148
rect 99189 82786 99255 82789
rect 166390 82786 166396 82788
rect 99189 82784 166396 82786
rect 99189 82728 99194 82784
rect 99250 82728 166396 82784
rect 99189 82726 166396 82728
rect 99189 82723 99255 82726
rect 166390 82724 166396 82726
rect 166460 82724 166466 82788
rect 262990 82724 262996 82788
rect 263060 82786 263066 82788
rect 335854 82786 335860 82788
rect 263060 82726 335860 82786
rect 263060 82724 263066 82726
rect 335854 82724 335860 82726
rect 335924 82724 335930 82788
rect 262990 81500 262996 81564
rect 263060 81562 263066 81564
rect 263501 81562 263567 81565
rect 263060 81560 263567 81562
rect 263060 81504 263506 81560
rect 263562 81504 263567 81560
rect 263060 81502 263567 81504
rect 263060 81500 263066 81502
rect 263501 81499 263567 81502
rect 106181 81426 106247 81429
rect 168966 81426 168972 81428
rect 106181 81424 168972 81426
rect 106181 81368 106186 81424
rect 106242 81368 168972 81424
rect 106181 81366 168972 81368
rect 106181 81363 106247 81366
rect 168966 81364 168972 81366
rect 169036 81364 169042 81428
rect 266854 81364 266860 81428
rect 266924 81426 266930 81428
rect 267641 81426 267707 81429
rect 338798 81426 338804 81428
rect 266924 81424 338804 81426
rect 266924 81368 267646 81424
rect 267702 81368 338804 81424
rect 266924 81366 338804 81368
rect 266924 81364 266930 81366
rect 267641 81363 267707 81366
rect 338798 81364 338804 81366
rect 338868 81364 338874 81428
rect 99281 80066 99347 80069
rect 170254 80066 170260 80068
rect 99281 80064 170260 80066
rect 99281 80008 99286 80064
rect 99342 80008 170260 80064
rect 99281 80006 170260 80008
rect 99281 80003 99347 80006
rect 170254 80004 170260 80006
rect 170324 80004 170330 80068
rect 108941 79930 109007 79933
rect 166206 79930 166212 79932
rect 108941 79928 166212 79930
rect 108941 79872 108946 79928
rect 109002 79872 166212 79928
rect 108941 79870 166212 79872
rect 108941 79867 109007 79870
rect 166206 79868 166212 79870
rect 166276 79868 166282 79932
rect 309726 77964 309732 78028
rect 309796 78026 309802 78028
rect 310513 78026 310579 78029
rect 309796 78024 310579 78026
rect 309796 77968 310518 78024
rect 310574 77968 310579 78024
rect 309796 77966 310579 77968
rect 309796 77964 309802 77966
rect 310513 77963 310579 77966
rect 173014 77828 173020 77892
rect 173084 77890 173090 77892
rect 246389 77890 246455 77893
rect 173084 77888 246455 77890
rect 173084 77832 246394 77888
rect 246450 77832 246455 77888
rect 173084 77830 246455 77832
rect 173084 77828 173090 77830
rect 246389 77827 246455 77830
rect 39941 77210 40007 77213
rect 321502 77210 321508 77212
rect 39941 77208 321508 77210
rect 39941 77152 39946 77208
rect 40002 77152 321508 77208
rect 39941 77150 321508 77152
rect 39941 77147 40007 77150
rect 321502 77148 321508 77150
rect 321572 77148 321578 77212
rect 12433 76530 12499 76533
rect 304390 76530 304396 76532
rect 12433 76528 304396 76530
rect 12433 76472 12438 76528
rect 12494 76472 304396 76528
rect 12433 76470 304396 76472
rect 12433 76467 12499 76470
rect 304390 76468 304396 76470
rect 304460 76468 304466 76532
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 61694 71028 61700 71092
rect 61764 71090 61770 71092
rect 274173 71090 274239 71093
rect 61764 71088 274239 71090
rect 61764 71032 274178 71088
rect 274234 71032 274239 71088
rect 61764 71030 274239 71032
rect 61764 71028 61770 71030
rect 274173 71027 274239 71030
rect 62982 69532 62988 69596
rect 63052 69594 63058 69596
rect 284334 69594 284340 69596
rect 63052 69534 284340 69594
rect 63052 69532 63058 69534
rect 284334 69532 284340 69534
rect 284404 69532 284410 69596
rect 286317 67554 286383 67557
rect 286961 67554 287027 67557
rect 477493 67554 477559 67557
rect 286317 67552 477559 67554
rect 286317 67496 286322 67552
rect 286378 67496 286966 67552
rect 287022 67496 477498 67552
rect 477554 67496 477559 67552
rect 286317 67494 477559 67496
rect 286317 67491 286383 67494
rect 286961 67491 287027 67494
rect 477493 67491 477559 67494
rect 60590 66812 60596 66876
rect 60660 66874 60666 66876
rect 332593 66874 332659 66877
rect 60660 66872 332659 66874
rect 60660 66816 332598 66872
rect 332654 66816 332659 66872
rect 60660 66814 332659 66816
rect 60660 66812 60666 66814
rect 332593 66811 332659 66814
rect 259545 65652 259611 65653
rect 259494 65588 259500 65652
rect 259564 65650 259611 65652
rect 259564 65648 259656 65650
rect 259606 65592 259656 65648
rect 259564 65590 259656 65592
rect 259564 65588 259611 65590
rect 259545 65587 259611 65588
rect 67633 64154 67699 64157
rect 302734 64154 302740 64156
rect 67633 64152 302740 64154
rect 67633 64096 67638 64152
rect 67694 64096 302740 64152
rect 67633 64094 302740 64096
rect 67633 64091 67699 64094
rect 302734 64092 302740 64094
rect 302804 64092 302810 64156
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 262806 57972 262812 58036
rect 262876 58034 262882 58036
rect 267733 58034 267799 58037
rect 262876 58032 267799 58034
rect 262876 57976 267738 58032
rect 267794 57976 267799 58032
rect 262876 57974 267799 57976
rect 262876 57972 262882 57974
rect 267733 57971 267799 57974
rect 49693 57218 49759 57221
rect 299974 57218 299980 57220
rect 49693 57216 299980 57218
rect 49693 57160 49698 57216
rect 49754 57160 299980 57216
rect 49693 57158 299980 57160
rect 49693 57155 49759 57158
rect 299974 57156 299980 57158
rect 300044 57156 300050 57220
rect 260046 56476 260052 56540
rect 260116 56538 260122 56540
rect 263593 56538 263659 56541
rect 260116 56536 263659 56538
rect 260116 56480 263598 56536
rect 263654 56480 263659 56536
rect 260116 56478 263659 56480
rect 260116 56476 260122 56478
rect 263593 56475 263659 56478
rect 284385 49060 284451 49061
rect 284334 48996 284340 49060
rect 284404 49058 284451 49060
rect 284404 49056 284496 49058
rect 284446 49000 284496 49056
rect 284404 48998 284496 49000
rect 284404 48996 284451 48998
rect 284385 48995 284451 48996
rect 269113 47564 269179 47565
rect 269062 47500 269068 47564
rect 269132 47562 269179 47564
rect 269132 47560 269224 47562
rect 269174 47504 269224 47560
rect 269132 47502 269224 47504
rect 269132 47500 269179 47502
rect 269113 47499 269179 47500
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 31753 46202 31819 46205
rect 334065 46204 334131 46205
rect 288934 46202 288940 46204
rect 31753 46200 288940 46202
rect 31753 46144 31758 46200
rect 31814 46144 288940 46200
rect 31753 46142 288940 46144
rect 31753 46139 31819 46142
rect 288934 46140 288940 46142
rect 289004 46140 289010 46204
rect 334014 46140 334020 46204
rect 334084 46202 334131 46204
rect 334084 46200 334176 46202
rect 334126 46144 334176 46200
rect 583520 46188 584960 46278
rect 334084 46142 334176 46144
rect 334084 46140 334131 46142
rect 334065 46139 334131 46140
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 268326 43420 268332 43484
rect 268396 43482 268402 43484
rect 318885 43482 318951 43485
rect 320081 43482 320147 43485
rect 268396 43480 320147 43482
rect 268396 43424 318890 43480
rect 318946 43424 320086 43480
rect 320142 43424 320147 43480
rect 268396 43422 320147 43424
rect 268396 43420 268402 43422
rect 318885 43419 318951 43422
rect 320081 43419 320147 43422
rect 298185 43348 298251 43349
rect 298134 43284 298140 43348
rect 298204 43346 298251 43348
rect 298204 43344 298296 43346
rect 298246 43288 298296 43344
rect 298204 43286 298296 43288
rect 298204 43284 298251 43286
rect 298185 43283 298251 43284
rect 273253 41306 273319 41309
rect 274173 41306 274239 41309
rect 345606 41306 345612 41308
rect 273253 41304 345612 41306
rect 273253 41248 273258 41304
rect 273314 41248 274178 41304
rect 274234 41248 345612 41304
rect 273253 41246 345612 41248
rect 273253 41243 273319 41246
rect 274173 41243 274239 41246
rect 345606 41244 345612 41246
rect 345676 41244 345682 41308
rect 302233 40764 302299 40765
rect 302182 40700 302188 40764
rect 302252 40762 302299 40764
rect 302252 40760 302344 40762
rect 302294 40704 302344 40760
rect 302252 40702 302344 40704
rect 302252 40700 302299 40702
rect 302233 40699 302299 40700
rect 299657 39404 299723 39405
rect 299606 39340 299612 39404
rect 299676 39402 299723 39404
rect 299676 39400 299768 39402
rect 299718 39344 299768 39400
rect 299676 39342 299768 39344
rect 299676 39340 299723 39342
rect 299657 39339 299723 39340
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 2865 28250 2931 28253
rect 304206 28250 304212 28252
rect 2865 28248 304212 28250
rect 2865 28192 2870 28248
rect 2926 28192 304212 28248
rect 2865 28190 304212 28192
rect 2865 28187 2931 28190
rect 304206 28188 304212 28190
rect 304276 28188 304282 28252
rect 270585 27028 270651 27029
rect 270534 26964 270540 27028
rect 270604 27026 270651 27028
rect 270604 27024 270696 27026
rect 270646 26968 270696 27024
rect 270604 26966 270696 26968
rect 270604 26964 270651 26966
rect 270585 26963 270651 26964
rect 9673 26890 9739 26893
rect 291694 26890 291700 26892
rect 9673 26888 291700 26890
rect 9673 26832 9678 26888
rect 9734 26832 291700 26888
rect 9673 26830 291700 26832
rect 9673 26827 9739 26830
rect 291694 26828 291700 26830
rect 291764 26828 291770 26892
rect 263542 24108 263548 24172
rect 263612 24170 263618 24172
rect 263685 24170 263751 24173
rect 263612 24168 263751 24170
rect 263612 24112 263690 24168
rect 263746 24112 263751 24168
rect 263612 24110 263751 24112
rect 263612 24108 263618 24110
rect 263685 24107 263751 24110
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 270534 12684 270540 12748
rect 270604 12746 270610 12748
rect 271781 12746 271847 12749
rect 270604 12744 271847 12746
rect 270604 12688 271786 12744
rect 271842 12688 271847 12744
rect 270604 12686 271847 12688
rect 270604 12684 270610 12686
rect 271781 12683 271847 12686
rect 262806 12276 262812 12340
rect 262876 12338 262882 12340
rect 268377 12338 268443 12341
rect 262876 12336 268443 12338
rect 262876 12280 268382 12336
rect 268438 12280 268443 12336
rect 262876 12278 268443 12280
rect 262876 12276 262882 12278
rect 268377 12275 268443 12278
rect 259494 11732 259500 11796
rect 259564 11794 259570 11796
rect 260741 11794 260807 11797
rect 259564 11792 260807 11794
rect 259564 11736 260746 11792
rect 260802 11736 260807 11792
rect 259564 11734 260807 11736
rect 259564 11732 259570 11734
rect 260741 11731 260807 11734
rect 263542 11732 263548 11796
rect 263612 11794 263618 11796
rect 264605 11794 264671 11797
rect 263612 11792 264671 11794
rect 263612 11736 264610 11792
rect 264666 11736 264671 11792
rect 263612 11734 264671 11736
rect 263612 11732 263618 11734
rect 264605 11731 264671 11734
rect 269062 11732 269068 11796
rect 269132 11794 269138 11796
rect 270309 11794 270375 11797
rect 269132 11792 270375 11794
rect 269132 11736 270314 11792
rect 270370 11736 270375 11792
rect 269132 11734 270375 11736
rect 269132 11732 269138 11734
rect 270309 11731 270375 11734
rect 284334 11732 284340 11796
rect 284404 11794 284410 11796
rect 285581 11794 285647 11797
rect 284404 11792 285647 11794
rect 284404 11736 285586 11792
rect 285642 11736 285647 11792
rect 284404 11734 285647 11736
rect 284404 11732 284410 11734
rect 285581 11731 285647 11734
rect 298134 11732 298140 11796
rect 298204 11794 298210 11796
rect 299381 11794 299447 11797
rect 298204 11792 299447 11794
rect 298204 11736 299386 11792
rect 299442 11736 299447 11792
rect 298204 11734 299447 11736
rect 298204 11732 298210 11734
rect 299381 11731 299447 11734
rect 299606 11732 299612 11796
rect 299676 11794 299682 11796
rect 300761 11794 300827 11797
rect 299676 11792 300827 11794
rect 299676 11736 300766 11792
rect 300822 11736 300827 11792
rect 299676 11734 300827 11736
rect 299676 11732 299682 11734
rect 300761 11731 300827 11734
rect 302182 11732 302188 11796
rect 302252 11794 302258 11796
rect 303521 11794 303587 11797
rect 302252 11792 303587 11794
rect 302252 11736 303526 11792
rect 303582 11736 303587 11792
rect 302252 11734 303587 11736
rect 302252 11732 302258 11734
rect 303521 11731 303587 11734
rect 310094 11732 310100 11796
rect 310164 11794 310170 11796
rect 312629 11794 312695 11797
rect 310164 11792 312695 11794
rect 310164 11736 312634 11792
rect 312690 11736 312695 11792
rect 310164 11734 312695 11736
rect 310164 11732 310170 11734
rect 312629 11731 312695 11734
rect 334014 11732 334020 11796
rect 334084 11794 334090 11796
rect 335077 11794 335143 11797
rect 334084 11792 335143 11794
rect 334084 11736 335082 11792
rect 335138 11736 335143 11792
rect 334084 11734 335143 11736
rect 334084 11732 334090 11734
rect 335077 11731 335143 11734
rect 342294 11732 342300 11796
rect 342364 11794 342370 11796
rect 343357 11794 343423 11797
rect 342364 11792 343423 11794
rect 342364 11736 343362 11792
rect 343418 11736 343423 11792
rect 342364 11734 343423 11736
rect 342364 11732 342370 11734
rect 343357 11731 343423 11734
rect 309726 11596 309732 11660
rect 309796 11658 309802 11660
rect 311433 11658 311499 11661
rect 309796 11656 311499 11658
rect 309796 11600 311438 11656
rect 311494 11600 311499 11656
rect 309796 11598 311499 11600
rect 309796 11596 309802 11598
rect 311433 11595 311499 11598
rect 61878 10916 61884 10980
rect 61948 10978 61954 10980
rect 242893 10978 242959 10981
rect 243537 10978 243603 10981
rect 258441 10980 258507 10981
rect 61948 10976 243603 10978
rect 61948 10920 242898 10976
rect 242954 10920 243542 10976
rect 243598 10920 243603 10976
rect 61948 10918 243603 10920
rect 61948 10916 61954 10918
rect 242893 10915 242959 10918
rect 243537 10915 243603 10918
rect 258390 10916 258396 10980
rect 258460 10978 258507 10980
rect 258460 10976 258552 10978
rect 258502 10920 258552 10976
rect 258460 10918 258552 10920
rect 258460 10916 258507 10918
rect 258441 10915 258507 10916
rect 287646 9556 287652 9620
rect 287716 9618 287722 9620
rect 300117 9618 300183 9621
rect 300669 9618 300735 9621
rect 287716 9616 300735 9618
rect 287716 9560 300122 9616
rect 300178 9560 300674 9616
rect 300730 9560 300735 9616
rect 287716 9558 300735 9560
rect 287716 9556 287722 9558
rect 300117 9555 300183 9558
rect 300669 9555 300735 9558
rect 373993 8938 374059 8941
rect 496854 8938 496860 8940
rect 373993 8936 496860 8938
rect 373993 8880 373998 8936
rect 374054 8880 496860 8936
rect 373993 8878 496860 8880
rect 373993 8875 374059 8878
rect 496854 8876 496860 8878
rect 496924 8876 496930 8940
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 299657 3634 299723 3637
rect 300761 3634 300827 3637
rect 299657 3632 300827 3634
rect 299657 3576 299662 3632
rect 299718 3576 300766 3632
rect 300822 3576 300827 3632
rect 299657 3574 300827 3576
rect 299657 3571 299723 3574
rect 300761 3571 300827 3574
rect 258257 3498 258323 3501
rect 259361 3498 259427 3501
rect 258257 3496 259427 3498
rect 258257 3440 258262 3496
rect 258318 3440 259366 3496
rect 259422 3440 259427 3496
rect 258257 3438 259427 3440
rect 258257 3435 258323 3438
rect 259361 3435 259427 3438
rect 262949 3498 263015 3501
rect 263501 3498 263567 3501
rect 262949 3496 263567 3498
rect 262949 3440 262954 3496
rect 263010 3440 263506 3496
rect 263562 3440 263567 3496
rect 262949 3438 263567 3440
rect 262949 3435 263015 3438
rect 263501 3435 263567 3438
rect 266537 3498 266603 3501
rect 267641 3498 267707 3501
rect 266537 3496 267707 3498
rect 266537 3440 266542 3496
rect 266598 3440 267646 3496
rect 267702 3440 267707 3496
rect 266537 3438 267707 3440
rect 266537 3435 266603 3438
rect 267641 3435 267707 3438
rect 271229 3498 271295 3501
rect 271781 3498 271847 3501
rect 271229 3496 271847 3498
rect 271229 3440 271234 3496
rect 271290 3440 271786 3496
rect 271842 3440 271847 3496
rect 271229 3438 271847 3440
rect 271229 3435 271295 3438
rect 271781 3435 271847 3438
rect 284293 3498 284359 3501
rect 285581 3498 285647 3501
rect 284293 3496 285647 3498
rect 284293 3440 284298 3496
rect 284354 3440 285586 3496
rect 285642 3440 285647 3496
rect 284293 3438 285647 3440
rect 284293 3435 284359 3438
rect 285581 3435 285647 3438
rect 298461 3498 298527 3501
rect 299381 3498 299447 3501
rect 298461 3496 299447 3498
rect 298461 3440 298466 3496
rect 298522 3440 299386 3496
rect 299442 3440 299447 3496
rect 298461 3438 299447 3440
rect 298461 3435 298527 3438
rect 299381 3435 299447 3438
rect 340822 3436 340828 3500
rect 340892 3498 340898 3500
rect 340965 3498 341031 3501
rect 342069 3498 342135 3501
rect 340892 3496 342135 3498
rect 340892 3440 340970 3496
rect 341026 3440 342074 3496
rect 342130 3440 342135 3496
rect 340892 3438 342135 3440
rect 340892 3436 340898 3438
rect 340965 3435 341031 3438
rect 342069 3435 342135 3438
rect 259453 3362 259519 3365
rect 260741 3362 260807 3365
rect 259453 3360 260807 3362
rect 259453 3304 259458 3360
rect 259514 3304 260746 3360
rect 260802 3304 260807 3360
rect 259453 3302 260807 3304
rect 259453 3299 259519 3302
rect 260741 3299 260807 3302
<< via3 >>
rect 111564 643180 111628 643244
rect 114508 586468 114572 586532
rect 53604 586332 53668 586396
rect 57652 583884 57716 583948
rect 118004 579940 118068 580004
rect 111748 577356 111812 577420
rect 107884 576676 107948 576740
rect 121684 572732 121748 572796
rect 66484 571780 66548 571844
rect 105492 571100 105556 571164
rect 65932 570284 65996 570348
rect 129780 570284 129844 570348
rect 66116 568924 66180 568988
rect 107700 563076 107764 563140
rect 69980 557364 70044 557428
rect 68876 553964 68940 554028
rect 111564 553964 111628 554028
rect 61884 549476 61948 549540
rect 125732 545668 125796 545732
rect 109540 541044 109604 541108
rect 107516 539956 107580 540020
rect 103652 538052 103716 538116
rect 109540 537916 109604 537980
rect 59124 537508 59188 537572
rect 57836 537372 57900 537436
rect 101260 537372 101324 537436
rect 53604 536012 53668 536076
rect 107884 535332 107948 535396
rect 108804 534652 108868 534716
rect 44036 529076 44100 529140
rect 114508 500380 114572 500444
rect 114508 500244 114572 500308
rect 111932 500108 111996 500172
rect 110644 499564 110708 499628
rect 136588 498748 136652 498812
rect 60596 494668 60660 494732
rect 52316 493308 52380 493372
rect 50292 492628 50356 492692
rect 48084 491812 48148 491876
rect 111012 491812 111076 491876
rect 99236 491268 99300 491332
rect 115060 491192 115124 491196
rect 115060 491136 115110 491192
rect 115110 491136 115124 491192
rect 115060 491132 115124 491136
rect 118004 489092 118068 489156
rect 118740 488608 118804 488612
rect 118740 488552 118790 488608
rect 118790 488552 118804 488608
rect 118740 488548 118804 488552
rect 99420 488004 99484 488068
rect 53604 487324 53668 487388
rect 57652 487324 57716 487388
rect 111748 485752 111812 485756
rect 111748 485696 111798 485752
rect 111798 485696 111812 485752
rect 111748 485692 111812 485696
rect 123340 485692 123404 485756
rect 70348 484604 70412 484668
rect 99972 484332 100036 484396
rect 123340 483244 123404 483308
rect 117084 481536 117148 481540
rect 117084 481480 117098 481536
rect 117098 481480 117148 481536
rect 117084 481476 117148 481480
rect 121684 481476 121748 481540
rect 69060 481068 69124 481132
rect 61700 480116 61764 480180
rect 104940 479768 105004 479772
rect 104940 479712 104990 479768
rect 104990 479712 105004 479768
rect 104940 479708 105004 479712
rect 65748 477668 65812 477732
rect 65932 477532 65996 477596
rect 62988 477396 63052 477460
rect 129780 477396 129844 477460
rect 106780 476172 106844 476236
rect 108988 476172 109052 476236
rect 55076 473996 55140 474060
rect 66484 473996 66548 474060
rect 66484 473724 66548 473788
rect 66668 473316 66732 473380
rect 107700 470596 107764 470660
rect 66116 470520 66180 470524
rect 66116 470464 66130 470520
rect 66130 470464 66180 470520
rect 66116 470460 66180 470464
rect 68140 454684 68204 454748
rect 68876 454684 68940 454748
rect 125732 453324 125796 453388
rect 107516 449440 107580 449444
rect 107516 449384 107530 449440
rect 107530 449384 107580 449440
rect 107516 449380 107580 449384
rect 61884 448564 61948 448628
rect 103836 445708 103900 445772
rect 128676 444892 128740 444956
rect 103836 444348 103900 444412
rect 114508 443668 114572 443732
rect 99420 442308 99484 442372
rect 110644 442308 110708 442372
rect 101260 441764 101324 441828
rect 99972 439724 100036 439788
rect 60596 439452 60660 439516
rect 70348 439452 70412 439516
rect 69060 438908 69124 438972
rect 111932 439452 111996 439516
rect 124812 438908 124876 438972
rect 57836 438092 57900 438156
rect 59124 437412 59188 437476
rect 106780 437412 106844 437476
rect 69060 433800 69124 433804
rect 69060 433744 69074 433800
rect 69074 433744 69124 433800
rect 69060 433740 69124 433744
rect 44036 433196 44100 433260
rect 115060 400208 115124 400212
rect 115060 400152 115110 400208
rect 115110 400152 115124 400208
rect 115060 400148 115124 400152
rect 48084 397972 48148 398036
rect 99052 397972 99116 398036
rect 111012 390628 111076 390692
rect 53604 390492 53668 390556
rect 136588 390492 136652 390556
rect 118740 389812 118804 389876
rect 53604 389132 53668 389196
rect 268332 389132 268396 389196
rect 52316 388316 52380 388380
rect 58572 388376 58636 388380
rect 58572 388320 58586 388376
rect 58586 388320 58636 388376
rect 58572 388316 58636 388320
rect 119292 387908 119356 387972
rect 119476 387772 119540 387836
rect 50292 387636 50356 387700
rect 54892 386956 54956 387020
rect 120028 386956 120092 387020
rect 299612 386956 299676 387020
rect 122604 386548 122668 386612
rect 262996 386412 263060 386476
rect 117820 386276 117884 386340
rect 61700 385052 61764 385116
rect 115796 385188 115860 385252
rect 65932 384780 65996 384844
rect 118004 384916 118068 384980
rect 115796 384508 115860 384572
rect 259500 384508 259564 384572
rect 65932 383888 65996 383892
rect 65932 383832 65946 383888
rect 65946 383832 65996 383888
rect 65932 383828 65996 383832
rect 122052 382196 122116 382260
rect 61884 380972 61948 381036
rect 62988 380972 63052 381036
rect 55076 380156 55140 380220
rect 129780 380156 129844 380220
rect 61700 379612 61764 379676
rect 66668 379612 66732 379676
rect 123340 378932 123404 378996
rect 60596 377980 60660 378044
rect 69980 377708 70044 377772
rect 60596 376756 60660 376820
rect 117084 376756 117148 376820
rect 262812 374580 262876 374644
rect 66116 373900 66180 373964
rect 287652 373220 287716 373284
rect 66116 372812 66180 372876
rect 117820 372676 117884 372740
rect 123340 372676 123404 372740
rect 335860 371316 335924 371380
rect 69060 370500 69124 370564
rect 119476 370500 119540 370564
rect 119292 369004 119356 369068
rect 62988 368324 63052 368388
rect 122052 368324 122116 368388
rect 68876 366012 68940 366076
rect 118924 364788 118988 364852
rect 65932 360980 65996 361044
rect 65380 360028 65444 360092
rect 65932 360028 65996 360092
rect 68140 357444 68204 357508
rect 123340 349692 123404 349756
rect 57100 347652 57164 347716
rect 126100 342408 126164 342412
rect 126100 342352 126150 342408
rect 126150 342352 126164 342408
rect 126100 342348 126164 342352
rect 70532 340988 70596 341052
rect 128676 339356 128740 339420
rect 55076 338132 55140 338196
rect 57836 337996 57900 338060
rect 120028 337996 120092 338060
rect 70532 335956 70596 336020
rect 258396 333236 258460 333300
rect 54892 332012 54956 332076
rect 270540 331740 270604 331804
rect 173020 330516 173084 330580
rect 68876 330380 68940 330444
rect 269068 329020 269132 329084
rect 70900 327660 70964 327724
rect 302188 326436 302252 326500
rect 65380 326300 65444 326364
rect 263548 326300 263612 326364
rect 309732 322084 309796 322148
rect 334020 319364 334084 319428
rect 342300 318004 342364 318068
rect 340828 316644 340892 316708
rect 124812 315964 124876 316028
rect 118740 315284 118804 315348
rect 124812 314740 124876 314804
rect 125732 314740 125796 314804
rect 122604 314256 122668 314260
rect 122604 314200 122618 314256
rect 122618 314200 122668 314256
rect 122604 314196 122668 314200
rect 266860 312428 266924 312492
rect 118924 307728 118988 307732
rect 118924 307672 118938 307728
rect 118938 307672 118988 307728
rect 118924 307668 118988 307672
rect 322980 302228 323044 302292
rect 122604 301412 122668 301476
rect 330340 300868 330404 300932
rect 326660 299508 326724 299572
rect 66116 298692 66180 298756
rect 298140 298692 298204 298756
rect 59124 295972 59188 296036
rect 121684 295564 121748 295628
rect 255268 295428 255332 295492
rect 58572 294476 58636 294540
rect 252508 289852 252572 289916
rect 119292 289444 119356 289508
rect 70532 285364 70596 285428
rect 121684 284336 121748 284340
rect 121684 284280 121698 284336
rect 121698 284280 121748 284336
rect 121684 284276 121748 284280
rect 256740 283460 256804 283524
rect 69060 279652 69124 279716
rect 327028 277748 327092 277812
rect 69244 257212 69308 257276
rect 125732 255308 125796 255372
rect 122604 249596 122668 249660
rect 122788 248236 122852 248300
rect 55076 242796 55140 242860
rect 58572 242796 58636 242860
rect 129780 241572 129844 241636
rect 119292 241164 119356 241228
rect 53604 240212 53668 240276
rect 70532 240212 70596 240276
rect 321508 239396 321572 239460
rect 59124 238580 59188 238644
rect 70532 237900 70596 237964
rect 334204 236540 334268 236604
rect 57100 235860 57164 235924
rect 173204 232596 173268 232660
rect 69060 232460 69124 232524
rect 320220 229740 320284 229804
rect 338620 225660 338684 225724
rect 69244 225524 69308 225588
rect 328500 220084 328564 220148
rect 494100 197916 494164 197980
rect 263732 193836 263796 193900
rect 58572 188260 58636 188324
rect 339540 184180 339604 184244
rect 118740 181324 118804 181388
rect 260052 181324 260116 181388
rect 258396 180100 258460 180164
rect 266308 179964 266372 180028
rect 214420 179420 214484 179484
rect 255452 178604 255516 178668
rect 112116 177924 112180 177988
rect 166212 178060 166276 178124
rect 97028 177712 97092 177716
rect 97028 177656 97078 177712
rect 97078 177656 97092 177712
rect 97028 177652 97092 177656
rect 100708 177652 100772 177716
rect 105676 177652 105740 177716
rect 110644 177712 110708 177716
rect 110644 177656 110694 177712
rect 110694 177656 110708 177712
rect 110644 177652 110708 177656
rect 114324 177712 114388 177716
rect 114324 177656 114374 177712
rect 114374 177656 114388 177712
rect 114324 177652 114388 177656
rect 118372 177652 118436 177716
rect 120764 177652 120828 177716
rect 125732 177652 125796 177716
rect 130700 177712 130764 177716
rect 130700 177656 130750 177712
rect 130750 177656 130764 177712
rect 130700 177652 130764 177656
rect 132356 177712 132420 177716
rect 132356 177656 132406 177712
rect 132406 177656 132420 177712
rect 132356 177652 132420 177656
rect 249380 177516 249444 177580
rect 331444 177380 331508 177444
rect 123156 177108 123220 177172
rect 108068 177032 108132 177036
rect 108068 176976 108118 177032
rect 108118 176976 108132 177032
rect 108068 176972 108132 176976
rect 113220 176972 113284 177036
rect 115796 177032 115860 177036
rect 115796 176976 115846 177032
rect 115846 176976 115860 177032
rect 115796 176972 115860 176976
rect 101996 176836 102060 176900
rect 168236 176836 168300 176900
rect 106964 176760 107028 176764
rect 106964 176704 107014 176760
rect 107014 176704 107028 176760
rect 106964 176700 107028 176704
rect 109540 176700 109604 176764
rect 119476 176760 119540 176764
rect 119476 176704 119526 176760
rect 119526 176704 119540 176760
rect 119476 176700 119540 176704
rect 121868 176700 121932 176764
rect 124444 176760 124508 176764
rect 124444 176704 124494 176760
rect 124494 176704 124508 176760
rect 124444 176700 124508 176704
rect 127020 176700 127084 176764
rect 133092 176760 133156 176764
rect 133092 176704 133142 176760
rect 133142 176704 133156 176760
rect 133092 176700 133156 176704
rect 134380 176760 134444 176764
rect 134380 176704 134430 176760
rect 134430 176704 134444 176760
rect 134380 176700 134444 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 269620 176700 269684 176764
rect 249748 176564 249812 176628
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 249196 175884 249260 175948
rect 98316 175476 98380 175540
rect 104572 175536 104636 175540
rect 104572 175480 104622 175536
rect 104622 175480 104636 175536
rect 104572 175476 104636 175480
rect 116900 175536 116964 175540
rect 116900 175480 116950 175536
rect 116950 175480 116964 175536
rect 116900 175476 116964 175480
rect 128124 175536 128188 175540
rect 128124 175480 128174 175536
rect 128174 175480 128188 175536
rect 128124 175476 128188 175480
rect 129412 175536 129476 175540
rect 129412 175480 129462 175536
rect 129462 175480 129476 175536
rect 129412 175476 129476 175480
rect 148180 175536 148244 175540
rect 148180 175480 148230 175536
rect 148230 175480 148244 175536
rect 148180 175476 148244 175480
rect 158852 175536 158916 175540
rect 158852 175480 158902 175536
rect 158902 175480 158916 175536
rect 158852 175476 158916 175480
rect 262076 175340 262140 175404
rect 335860 174524 335924 174588
rect 249196 174252 249260 174316
rect 249380 173708 249444 173772
rect 336044 172484 336108 172548
rect 496860 173300 496924 173364
rect 321324 169492 321388 169556
rect 335860 168404 335924 168468
rect 255452 166228 255516 166292
rect 338804 165684 338868 165748
rect 166212 162828 166276 162892
rect 345612 162828 345676 162892
rect 214420 162012 214484 162076
rect 168236 160652 168300 160716
rect 263732 160788 263796 160852
rect 252508 159156 252572 159220
rect 255268 157252 255332 157316
rect 258396 153716 258460 153780
rect 307156 149772 307220 149836
rect 251772 149636 251836 149700
rect 168236 145012 168300 145076
rect 306972 145012 307036 145076
rect 321508 144876 321572 144940
rect 266308 142156 266372 142220
rect 306972 139980 307036 140044
rect 304212 139708 304276 139772
rect 256740 137532 256804 137596
rect 307156 137260 307220 137324
rect 249748 136988 249812 137052
rect 306972 136988 307036 137052
rect 170444 134132 170508 134196
rect 330340 134132 330404 134196
rect 322980 133996 323044 134060
rect 166212 132772 166276 132836
rect 302740 132636 302804 132700
rect 168972 131412 169036 131476
rect 299980 130052 300044 130116
rect 170260 128556 170324 128620
rect 288940 128692 289004 128756
rect 494100 127876 494164 127940
rect 166396 127060 166460 127124
rect 291700 125836 291764 125900
rect 327028 126244 327092 126308
rect 255820 123116 255884 123180
rect 251772 116860 251836 116924
rect 331444 116452 331508 116516
rect 338620 115908 338684 115972
rect 307156 113596 307220 113660
rect 304396 113460 304460 113524
rect 252508 111012 252572 111076
rect 334204 110604 334268 110668
rect 252508 109788 252572 109852
rect 339540 109108 339604 109172
rect 326660 107068 326724 107132
rect 328500 106252 328564 106316
rect 172100 103532 172164 103596
rect 214420 102444 214484 102508
rect 309732 101764 309796 101828
rect 169156 101356 169220 101420
rect 324268 99316 324332 99380
rect 321508 97956 321572 98020
rect 262076 97276 262140 97340
rect 269620 97140 269684 97204
rect 173204 95508 173268 95572
rect 151492 94556 151556 94620
rect 151766 94556 151830 94620
rect 255820 94420 255884 94484
rect 126468 94208 126532 94212
rect 126468 94152 126518 94208
rect 126518 94152 126532 94208
rect 126468 94148 126532 94152
rect 152044 94208 152108 94212
rect 152044 94152 152094 94208
rect 152094 94152 152108 94208
rect 152044 94148 152108 94152
rect 112300 94072 112364 94076
rect 112300 94016 112350 94072
rect 112350 94016 112364 94072
rect 112300 94012 112364 94016
rect 126652 94072 126716 94076
rect 126652 94016 126702 94072
rect 126702 94016 126716 94072
rect 126652 94012 126716 94016
rect 96108 93936 96172 93940
rect 96108 93880 96158 93936
rect 96158 93880 96172 93936
rect 96108 93876 96172 93880
rect 100892 93528 100956 93532
rect 100892 93472 100942 93528
rect 100942 93472 100956 93528
rect 100892 93468 100956 93472
rect 109172 93528 109236 93532
rect 109172 93472 109222 93528
rect 109222 93472 109236 93528
rect 109172 93468 109236 93472
rect 116716 93528 116780 93532
rect 116716 93472 116766 93528
rect 116766 93472 116780 93528
rect 116716 93468 116780 93472
rect 121684 93528 121748 93532
rect 121684 93472 121734 93528
rect 121734 93472 121748 93528
rect 121684 93468 121748 93472
rect 133092 93528 133156 93532
rect 133092 93472 133142 93528
rect 133142 93472 133156 93528
rect 133092 93468 133156 93472
rect 151676 93528 151740 93532
rect 151676 93472 151726 93528
rect 151726 93472 151740 93528
rect 151676 93468 151740 93472
rect 324268 93468 324332 93532
rect 103284 93256 103348 93260
rect 103284 93200 103334 93256
rect 103334 93200 103348 93256
rect 103284 93196 103348 93200
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 74764 92440 74828 92444
rect 74764 92384 74814 92440
rect 74814 92384 74828 92440
rect 74764 92380 74828 92384
rect 85804 92440 85868 92444
rect 85804 92384 85854 92440
rect 85854 92384 85868 92440
rect 85804 92380 85868 92384
rect 88012 92440 88076 92444
rect 88012 92384 88062 92440
rect 88062 92384 88076 92440
rect 88012 92380 88076 92384
rect 88932 92440 88996 92444
rect 88932 92384 88982 92440
rect 88982 92384 88996 92440
rect 88932 92380 88996 92384
rect 97212 92380 97276 92444
rect 98500 92380 98564 92444
rect 113036 92380 113100 92444
rect 114876 92440 114940 92444
rect 114876 92384 114926 92440
rect 114926 92384 114940 92440
rect 114876 92380 114940 92384
rect 115428 92440 115492 92444
rect 115428 92384 115478 92440
rect 115478 92384 115492 92440
rect 115428 92380 115492 92384
rect 118004 92440 118068 92444
rect 118004 92384 118054 92440
rect 118054 92384 118068 92440
rect 118004 92380 118068 92384
rect 132356 92440 132420 92444
rect 132356 92384 132406 92440
rect 132406 92384 132420 92440
rect 132356 92380 132420 92384
rect 151492 92440 151556 92444
rect 151492 92384 151542 92440
rect 151542 92384 151556 92440
rect 151492 92380 151556 92384
rect 102732 92244 102796 92308
rect 122052 92244 122116 92308
rect 169156 92244 169220 92308
rect 122788 92168 122852 92172
rect 122788 92112 122838 92168
rect 122838 92112 122852 92168
rect 122788 92108 122852 92112
rect 151308 92108 151372 92172
rect 90220 91700 90284 91764
rect 119292 91564 119356 91628
rect 136036 91564 136100 91628
rect 93900 91292 93964 91356
rect 98132 91292 98196 91356
rect 100524 91352 100588 91356
rect 100524 91296 100574 91352
rect 100574 91296 100588 91352
rect 100524 91292 100588 91296
rect 101812 91352 101876 91356
rect 101812 91296 101862 91352
rect 101862 91296 101876 91352
rect 101812 91292 101876 91296
rect 105492 91292 105556 91356
rect 106412 91292 106476 91356
rect 120580 91292 120644 91356
rect 124076 91352 124140 91356
rect 124076 91296 124090 91352
rect 124090 91296 124140 91352
rect 124076 91292 124140 91296
rect 124444 91292 124508 91356
rect 84332 91156 84396 91220
rect 86724 91216 86788 91220
rect 86724 91160 86774 91216
rect 86774 91160 86788 91216
rect 86724 91156 86788 91160
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91156 95068 91220
rect 96660 91156 96724 91220
rect 99052 91156 99116 91220
rect 99972 91156 100036 91220
rect 101996 91216 102060 91220
rect 101996 91160 102046 91216
rect 102046 91160 102060 91216
rect 101996 91156 102060 91160
rect 104204 91216 104268 91220
rect 104204 91160 104254 91216
rect 104254 91160 104268 91216
rect 104204 91156 104268 91160
rect 104572 91156 104636 91220
rect 105676 91156 105740 91220
rect 106780 91156 106844 91220
rect 107700 91156 107764 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 110644 91216 110708 91220
rect 110644 91160 110694 91216
rect 110694 91160 110708 91216
rect 110644 91156 110708 91160
rect 111196 91156 111260 91220
rect 111932 91156 111996 91220
rect 113220 91156 113284 91220
rect 114324 91216 114388 91220
rect 114324 91160 114374 91216
rect 114374 91160 114388 91216
rect 114324 91156 114388 91160
rect 115796 91216 115860 91220
rect 115796 91160 115810 91216
rect 115810 91160 115860 91216
rect 115796 91156 115860 91160
rect 117084 91216 117148 91220
rect 117084 91160 117134 91216
rect 117134 91160 117148 91216
rect 117084 91156 117148 91160
rect 118188 91156 118252 91220
rect 119660 91156 119724 91220
rect 120212 91156 120276 91220
rect 123156 91156 123220 91220
rect 125364 91156 125428 91220
rect 125732 91156 125796 91220
rect 129412 91216 129476 91220
rect 129412 91160 129462 91216
rect 129462 91160 129476 91216
rect 129412 91156 129476 91160
rect 130700 91216 130764 91220
rect 130700 91160 130750 91216
rect 130750 91160 130764 91216
rect 130700 91156 130764 91160
rect 134380 91156 134444 91220
rect 214420 91020 214484 91084
rect 127572 90884 127636 90948
rect 307156 90340 307220 90404
rect 310100 90340 310164 90404
rect 170444 88164 170508 88228
rect 342300 87680 342364 87684
rect 342300 87624 342350 87680
rect 342350 87624 342364 87680
rect 342300 87620 342364 87624
rect 336044 86124 336108 86188
rect 168236 85444 168300 85508
rect 306972 84764 307036 84828
rect 172100 84084 172164 84148
rect 166396 82724 166460 82788
rect 262996 82724 263060 82788
rect 335860 82724 335924 82788
rect 262996 81500 263060 81564
rect 168972 81364 169036 81428
rect 266860 81364 266924 81428
rect 338804 81364 338868 81428
rect 170260 80004 170324 80068
rect 166212 79868 166276 79932
rect 309732 77964 309796 78028
rect 173020 77828 173084 77892
rect 321508 77148 321572 77212
rect 304396 76468 304460 76532
rect 61700 71028 61764 71092
rect 62988 69532 63052 69596
rect 284340 69532 284404 69596
rect 60596 66812 60660 66876
rect 259500 65648 259564 65652
rect 259500 65592 259550 65648
rect 259550 65592 259564 65648
rect 259500 65588 259564 65592
rect 302740 64092 302804 64156
rect 262812 57972 262876 58036
rect 299980 57156 300044 57220
rect 260052 56476 260116 56540
rect 284340 49056 284404 49060
rect 284340 49000 284390 49056
rect 284390 49000 284404 49056
rect 284340 48996 284404 49000
rect 269068 47560 269132 47564
rect 269068 47504 269118 47560
rect 269118 47504 269132 47560
rect 269068 47500 269132 47504
rect 288940 46140 289004 46204
rect 334020 46200 334084 46204
rect 334020 46144 334070 46200
rect 334070 46144 334084 46200
rect 334020 46140 334084 46144
rect 268332 43420 268396 43484
rect 298140 43344 298204 43348
rect 298140 43288 298190 43344
rect 298190 43288 298204 43344
rect 298140 43284 298204 43288
rect 345612 41244 345676 41308
rect 302188 40760 302252 40764
rect 302188 40704 302238 40760
rect 302238 40704 302252 40760
rect 302188 40700 302252 40704
rect 299612 39400 299676 39404
rect 299612 39344 299662 39400
rect 299662 39344 299676 39400
rect 299612 39340 299676 39344
rect 304212 28188 304276 28252
rect 270540 27024 270604 27028
rect 270540 26968 270590 27024
rect 270590 26968 270604 27024
rect 270540 26964 270604 26968
rect 291700 26828 291764 26892
rect 263548 24108 263612 24172
rect 270540 12684 270604 12748
rect 262812 12276 262876 12340
rect 259500 11732 259564 11796
rect 263548 11732 263612 11796
rect 269068 11732 269132 11796
rect 284340 11732 284404 11796
rect 298140 11732 298204 11796
rect 299612 11732 299676 11796
rect 302188 11732 302252 11796
rect 310100 11732 310164 11796
rect 334020 11732 334084 11796
rect 342300 11732 342364 11796
rect 309732 11596 309796 11660
rect 61884 10916 61948 10980
rect 258396 10976 258460 10980
rect 258396 10920 258446 10976
rect 258446 10920 258460 10976
rect 258396 10916 258460 10920
rect 287652 9556 287716 9620
rect 496860 8876 496924 8940
rect 340828 3436 340892 3500
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 44035 529140 44101 529141
rect 44035 529076 44036 529140
rect 44100 529076 44101 529140
rect 44035 529075 44101 529076
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 44038 433261 44098 529075
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 53603 586396 53669 586397
rect 53603 586332 53604 586396
rect 53668 586332 53669 586396
rect 53603 586331 53669 586332
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 53606 536077 53666 586331
rect 55794 561454 56414 596898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 57651 583948 57717 583949
rect 57651 583884 57652 583948
rect 57716 583884 57717 583948
rect 57651 583883 57717 583884
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 53603 536076 53669 536077
rect 53603 536012 53604 536076
rect 53668 536012 53669 536076
rect 53603 536011 53669 536012
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48083 491876 48149 491877
rect 48083 491812 48084 491876
rect 48148 491812 48149 491876
rect 48083 491811 48149 491812
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 44035 433260 44101 433261
rect 44035 433196 44036 433260
rect 44100 433196 44101 433260
rect 44035 433195 44101 433196
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 48086 398037 48146 491811
rect 48954 482614 49574 518058
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 52315 493372 52381 493373
rect 52315 493308 52316 493372
rect 52380 493308 52381 493372
rect 52315 493307 52381 493308
rect 50291 492692 50357 492693
rect 50291 492628 50292 492692
rect 50356 492628 50357 492692
rect 50291 492627 50357 492628
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48083 398036 48149 398037
rect 48083 397972 48084 398036
rect 48148 397972 48149 398036
rect 48083 397971 48149 397972
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 374614 49574 410058
rect 50294 387701 50354 492627
rect 52318 388381 52378 493307
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 53603 487388 53669 487389
rect 53603 487324 53604 487388
rect 53668 487324 53669 487388
rect 53603 487323 53669 487324
rect 53606 390557 53666 487323
rect 55075 474060 55141 474061
rect 55075 473996 55076 474060
rect 55140 473996 55141 474060
rect 55075 473995 55141 473996
rect 53603 390556 53669 390557
rect 53603 390492 53604 390556
rect 53668 390492 53669 390556
rect 53603 390491 53669 390492
rect 53603 389196 53669 389197
rect 53603 389132 53604 389196
rect 53668 389132 53669 389196
rect 53603 389131 53669 389132
rect 52315 388380 52381 388381
rect 52315 388316 52316 388380
rect 52380 388316 52381 388380
rect 52315 388315 52381 388316
rect 50291 387700 50357 387701
rect 50291 387636 50292 387700
rect 50356 387636 50357 387700
rect 50291 387635 50357 387636
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 53606 240277 53666 389131
rect 54891 387020 54957 387021
rect 54891 386956 54892 387020
rect 54956 386956 54957 387020
rect 54891 386955 54957 386956
rect 54894 332077 54954 386955
rect 55078 380221 55138 473995
rect 55794 453454 56414 488898
rect 57654 487389 57714 583883
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59123 537572 59189 537573
rect 59123 537508 59124 537572
rect 59188 537508 59189 537572
rect 59123 537507 59189 537508
rect 57835 537436 57901 537437
rect 57835 537372 57836 537436
rect 57900 537372 57901 537436
rect 57835 537371 57901 537372
rect 57651 487388 57717 487389
rect 57651 487324 57652 487388
rect 57716 487324 57717 487388
rect 57651 487323 57717 487324
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 57838 438157 57898 537371
rect 57835 438156 57901 438157
rect 57835 438092 57836 438156
rect 57900 438092 57901 438156
rect 57835 438091 57901 438092
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55075 380220 55141 380221
rect 55075 380156 55076 380220
rect 55140 380156 55141 380220
rect 55075 380155 55141 380156
rect 55794 345454 56414 380898
rect 57099 347716 57165 347717
rect 57099 347652 57100 347716
rect 57164 347652 57165 347716
rect 57099 347651 57165 347652
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55075 338196 55141 338197
rect 55075 338132 55076 338196
rect 55140 338132 55141 338196
rect 55075 338131 55141 338132
rect 54891 332076 54957 332077
rect 54891 332012 54892 332076
rect 54956 332012 54957 332076
rect 54891 332011 54957 332012
rect 55078 242861 55138 338131
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55075 242860 55141 242861
rect 55075 242796 55076 242860
rect 55140 242796 55141 242860
rect 55075 242795 55141 242796
rect 53603 240276 53669 240277
rect 53603 240212 53604 240276
rect 53668 240212 53669 240276
rect 53603 240211 53669 240212
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 57102 235925 57162 347651
rect 57838 338061 57898 438091
rect 59126 437477 59186 537507
rect 59514 529174 60134 564618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 584000 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 584000 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 584000 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 584000 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 584000 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 584000 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 584000 99854 604338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 584000 103574 608058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 111563 643244 111629 643245
rect 111563 643180 111564 643244
rect 111628 643180 111629 643244
rect 111563 643179 111629 643180
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 76576 579454 76896 579486
rect 76576 579218 76618 579454
rect 76854 579218 76896 579454
rect 76576 579134 76896 579218
rect 76576 578898 76618 579134
rect 76854 578898 76896 579134
rect 76576 578866 76896 578898
rect 87840 579454 88160 579486
rect 87840 579218 87882 579454
rect 88118 579218 88160 579454
rect 87840 579134 88160 579218
rect 87840 578898 87882 579134
rect 88118 578898 88160 579134
rect 87840 578866 88160 578898
rect 99104 579454 99424 579486
rect 99104 579218 99146 579454
rect 99382 579218 99424 579454
rect 99104 579134 99424 579218
rect 99104 578898 99146 579134
rect 99382 578898 99424 579134
rect 99104 578866 99424 578898
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 107883 576740 107949 576741
rect 107883 576676 107884 576740
rect 107948 576676 107949 576740
rect 107883 576675 107949 576676
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66483 571844 66549 571845
rect 66483 571780 66484 571844
rect 66548 571780 66549 571844
rect 66483 571779 66549 571780
rect 65931 570348 65997 570349
rect 65931 570284 65932 570348
rect 65996 570284 65997 570348
rect 65931 570283 65997 570284
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 61883 549540 61949 549541
rect 61883 549476 61884 549540
rect 61948 549476 61949 549540
rect 61883 549475 61949 549476
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 60595 494732 60661 494733
rect 60595 494668 60596 494732
rect 60660 494668 60661 494732
rect 60595 494667 60661 494668
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59123 437476 59189 437477
rect 59123 437412 59124 437476
rect 59188 437412 59189 437476
rect 59123 437411 59189 437412
rect 59514 421174 60134 456618
rect 60598 439517 60658 494667
rect 61699 480180 61765 480181
rect 61699 480116 61700 480180
rect 61764 480116 61765 480180
rect 61699 480115 61765 480116
rect 60595 439516 60661 439517
rect 60595 439452 60596 439516
rect 60660 439452 60661 439516
rect 60595 439451 60661 439452
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 58571 388380 58637 388381
rect 58571 388316 58572 388380
rect 58636 388316 58637 388380
rect 58571 388315 58637 388316
rect 57835 338060 57901 338061
rect 57835 337996 57836 338060
rect 57900 337996 57901 338060
rect 57835 337995 57901 337996
rect 58574 294541 58634 388315
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 61702 385117 61762 480115
rect 61886 448629 61946 549475
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 62987 477460 63053 477461
rect 62987 477396 62988 477460
rect 63052 477396 63053 477460
rect 62987 477395 63053 477396
rect 61883 448628 61949 448629
rect 61883 448564 61884 448628
rect 61948 448564 61949 448628
rect 61883 448563 61949 448564
rect 61699 385116 61765 385117
rect 61699 385052 61700 385116
rect 61764 385052 61765 385116
rect 61699 385051 61765 385052
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 62990 381037 63050 477395
rect 63234 460894 63854 496338
rect 65747 477732 65813 477733
rect 65747 477668 65748 477732
rect 65812 477668 65813 477732
rect 65747 477667 65813 477668
rect 65750 476130 65810 477667
rect 65934 477597 65994 570283
rect 66115 568988 66181 568989
rect 66115 568924 66116 568988
rect 66180 568924 66181 568988
rect 66115 568923 66181 568924
rect 65931 477596 65997 477597
rect 65931 477532 65932 477596
rect 65996 477532 65997 477596
rect 65931 477531 65997 477532
rect 65750 476070 65994 476130
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 61883 381036 61949 381037
rect 61883 380972 61884 381036
rect 61948 380972 61949 381036
rect 61883 380971 61949 380972
rect 62987 381036 63053 381037
rect 62987 380972 62988 381036
rect 63052 380972 63053 381036
rect 62987 380971 63053 380972
rect 61699 379676 61765 379677
rect 61699 379612 61700 379676
rect 61764 379612 61765 379676
rect 61699 379611 61765 379612
rect 60595 378044 60661 378045
rect 60595 377980 60596 378044
rect 60660 377980 60661 378044
rect 60595 377979 60661 377980
rect 60598 376821 60658 377979
rect 60595 376820 60661 376821
rect 60595 376756 60596 376820
rect 60660 376756 60661 376820
rect 60595 376755 60661 376756
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59123 296036 59189 296037
rect 59123 295972 59124 296036
rect 59188 295972 59189 296036
rect 59123 295971 59189 295972
rect 58571 294540 58637 294541
rect 58571 294476 58572 294540
rect 58636 294476 58637 294540
rect 58571 294475 58637 294476
rect 58571 242860 58637 242861
rect 58571 242796 58572 242860
rect 58636 242796 58637 242860
rect 58571 242795 58637 242796
rect 57099 235924 57165 235925
rect 57099 235860 57100 235924
rect 57164 235860 57165 235924
rect 57099 235859 57165 235860
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 58574 188325 58634 242795
rect 59126 238645 59186 295971
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59123 238644 59189 238645
rect 59123 238580 59124 238644
rect 59188 238580 59189 238644
rect 59123 238579 59189 238580
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 58571 188324 58637 188325
rect 58571 188260 58572 188324
rect 58636 188260 58637 188324
rect 58571 188259 58637 188260
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 60598 66877 60658 376755
rect 61702 71093 61762 379611
rect 61699 71092 61765 71093
rect 61699 71028 61700 71092
rect 61764 71028 61765 71092
rect 61699 71027 61765 71028
rect 60595 66876 60661 66877
rect 60595 66812 60596 66876
rect 60660 66812 60661 66876
rect 60595 66811 60661 66812
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 61886 10981 61946 380971
rect 62987 368388 63053 368389
rect 62987 368324 62988 368388
rect 63052 368324 63053 368388
rect 62987 368323 63053 368324
rect 62990 69597 63050 368323
rect 63234 352894 63854 388338
rect 65934 384845 65994 476070
rect 66118 470525 66178 568923
rect 66486 474061 66546 571779
rect 66954 536614 67574 572058
rect 105491 571164 105557 571165
rect 105491 571100 105492 571164
rect 105556 571100 105557 571164
rect 105491 571099 105557 571100
rect 105494 567210 105554 571099
rect 104942 567150 105554 567210
rect 82208 561454 82528 561486
rect 82208 561218 82250 561454
rect 82486 561218 82528 561454
rect 82208 561134 82528 561218
rect 82208 560898 82250 561134
rect 82486 560898 82528 561134
rect 82208 560866 82528 560898
rect 93472 561454 93792 561486
rect 93472 561218 93514 561454
rect 93750 561218 93792 561454
rect 93472 561134 93792 561218
rect 93472 560898 93514 561134
rect 93750 560898 93792 561134
rect 93472 560866 93792 560898
rect 69979 557428 70045 557429
rect 69979 557364 69980 557428
rect 70044 557364 70045 557428
rect 69979 557363 70045 557364
rect 69982 557290 70042 557363
rect 69982 557230 70410 557290
rect 68875 554028 68941 554029
rect 68875 553964 68876 554028
rect 68940 553964 68941 554028
rect 68875 553963 68941 553964
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66483 474060 66549 474061
rect 66483 473996 66484 474060
rect 66548 473996 66549 474060
rect 66483 473995 66549 473996
rect 66486 473789 66546 473995
rect 66483 473788 66549 473789
rect 66483 473724 66484 473788
rect 66548 473724 66549 473788
rect 66483 473723 66549 473724
rect 66667 473380 66733 473381
rect 66667 473316 66668 473380
rect 66732 473316 66733 473380
rect 66667 473315 66733 473316
rect 66115 470524 66181 470525
rect 66115 470460 66116 470524
rect 66180 470460 66181 470524
rect 66115 470459 66181 470460
rect 65931 384844 65997 384845
rect 65931 384780 65932 384844
rect 65996 384780 65997 384844
rect 65931 384779 65997 384780
rect 65934 383893 65994 384779
rect 65931 383892 65997 383893
rect 65931 383828 65932 383892
rect 65996 383828 65997 383892
rect 65931 383827 65997 383828
rect 66670 379677 66730 473315
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 68878 454749 68938 553963
rect 70350 484669 70410 557230
rect 76576 543454 76896 543486
rect 76576 543218 76618 543454
rect 76854 543218 76896 543454
rect 76576 543134 76896 543218
rect 76576 542898 76618 543134
rect 76854 542898 76896 543134
rect 76576 542866 76896 542898
rect 87840 543454 88160 543486
rect 87840 543218 87882 543454
rect 88118 543218 88160 543454
rect 87840 543134 88160 543218
rect 87840 542898 87882 543134
rect 88118 542898 88160 543134
rect 87840 542866 88160 542898
rect 99104 543454 99424 543486
rect 99104 543218 99146 543454
rect 99382 543218 99424 543454
rect 99104 543134 99424 543218
rect 99104 542898 99146 543134
rect 99382 542898 99424 543134
rect 99104 542866 99424 542898
rect 103651 538116 103717 538117
rect 103651 538052 103652 538116
rect 103716 538052 103717 538116
rect 103651 538051 103717 538052
rect 73794 507454 74414 538000
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 492000 74414 506898
rect 77514 511174 78134 538000
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 492000 78134 510618
rect 81234 514894 81854 538000
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 492000 81854 514338
rect 84954 518614 85574 538000
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 492000 85574 518058
rect 91794 525454 92414 538000
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 492000 92414 524898
rect 95514 529174 96134 538000
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 492000 96134 492618
rect 99234 532894 99854 538000
rect 101259 537436 101325 537437
rect 101259 537372 101260 537436
rect 101324 537372 101325 537436
rect 101259 537371 101325 537372
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 492000 99854 496338
rect 99235 491332 99301 491333
rect 99235 491268 99236 491332
rect 99300 491268 99301 491332
rect 99235 491267 99301 491268
rect 99238 487930 99298 491267
rect 99419 488068 99485 488069
rect 99419 488004 99420 488068
rect 99484 488004 99485 488068
rect 99419 488003 99485 488004
rect 99422 487930 99482 488003
rect 99238 487870 99482 487930
rect 70347 484668 70413 484669
rect 70347 484604 70348 484668
rect 70412 484604 70413 484668
rect 70347 484603 70413 484604
rect 99971 484396 100037 484397
rect 99971 484332 99972 484396
rect 100036 484332 100037 484396
rect 99971 484331 100037 484332
rect 69059 481132 69125 481133
rect 69059 481068 69060 481132
rect 69124 481068 69125 481132
rect 69059 481067 69125 481068
rect 68139 454748 68205 454749
rect 68139 454684 68140 454748
rect 68204 454684 68205 454748
rect 68139 454683 68205 454684
rect 68875 454748 68941 454749
rect 68875 454684 68876 454748
rect 68940 454684 68941 454748
rect 68875 454683 68941 454684
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66667 379676 66733 379677
rect 66667 379612 66668 379676
rect 66732 379612 66733 379676
rect 66667 379611 66733 379612
rect 66115 373964 66181 373965
rect 66115 373900 66116 373964
rect 66180 373900 66181 373964
rect 66115 373899 66181 373900
rect 66118 372877 66178 373899
rect 66115 372876 66181 372877
rect 66115 372812 66116 372876
rect 66180 372812 66181 372876
rect 66115 372811 66181 372812
rect 65931 361044 65997 361045
rect 65931 360980 65932 361044
rect 65996 360980 65997 361044
rect 65931 360979 65997 360980
rect 65934 360093 65994 360979
rect 65379 360092 65445 360093
rect 65379 360028 65380 360092
rect 65444 360028 65445 360092
rect 65379 360027 65445 360028
rect 65931 360092 65997 360093
rect 65931 360028 65932 360092
rect 65996 360028 65997 360092
rect 65931 360027 65997 360028
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 65382 326365 65442 360027
rect 65379 326364 65445 326365
rect 65379 326300 65380 326364
rect 65444 326300 65445 326364
rect 65379 326299 65445 326300
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 66118 298757 66178 372811
rect 66954 356614 67574 392058
rect 68142 357509 68202 454683
rect 69062 438973 69122 481067
rect 75576 471454 75896 471486
rect 75576 471218 75618 471454
rect 75854 471218 75896 471454
rect 75576 471134 75896 471218
rect 75576 470898 75618 471134
rect 75854 470898 75896 471134
rect 75576 470866 75896 470898
rect 84840 471454 85160 471486
rect 84840 471218 84882 471454
rect 85118 471218 85160 471454
rect 84840 471134 85160 471218
rect 84840 470898 84882 471134
rect 85118 470898 85160 471134
rect 84840 470866 85160 470898
rect 94104 471454 94424 471486
rect 94104 471218 94146 471454
rect 94382 471218 94424 471454
rect 94104 471134 94424 471218
rect 94104 470898 94146 471134
rect 94382 470898 94424 471134
rect 94104 470866 94424 470898
rect 80208 453454 80528 453486
rect 80208 453218 80250 453454
rect 80486 453218 80528 453454
rect 80208 453134 80528 453218
rect 80208 452898 80250 453134
rect 80486 452898 80528 453134
rect 80208 452866 80528 452898
rect 89472 453454 89792 453486
rect 89472 453218 89514 453454
rect 89750 453218 89792 453454
rect 89472 453134 89792 453218
rect 89472 452898 89514 453134
rect 89750 452898 89792 453134
rect 89472 452866 89792 452898
rect 99419 442372 99485 442373
rect 99419 442370 99420 442372
rect 99054 442310 99420 442370
rect 70347 439516 70413 439517
rect 70347 439452 70348 439516
rect 70412 439452 70413 439516
rect 70347 439451 70413 439452
rect 69059 438972 69125 438973
rect 69059 438908 69060 438972
rect 69124 438908 69125 438972
rect 69059 438907 69125 438908
rect 69059 433804 69125 433805
rect 69059 433740 69060 433804
rect 69124 433740 69125 433804
rect 69059 433739 69125 433740
rect 69062 370565 69122 433739
rect 69979 377772 70045 377773
rect 69979 377708 69980 377772
rect 70044 377770 70045 377772
rect 70350 377770 70410 439451
rect 73794 435454 74414 438000
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 388000 74414 398898
rect 77514 403174 78134 438000
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 388000 78134 402618
rect 81234 406894 81854 438000
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 388000 81854 406338
rect 84954 410614 85574 438000
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 388000 85574 410058
rect 91794 417454 92414 438000
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 388000 92414 416898
rect 95514 421174 96134 438000
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 388000 96134 420618
rect 99054 398037 99114 442310
rect 99419 442308 99420 442310
rect 99484 442308 99485 442372
rect 99419 442307 99485 442308
rect 99974 439789 100034 484331
rect 101262 441829 101322 537371
rect 102954 536614 103574 538000
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 101259 441828 101325 441829
rect 101259 441764 101260 441828
rect 101324 441764 101325 441828
rect 101259 441763 101325 441764
rect 99971 439788 100037 439789
rect 99971 439724 99972 439788
rect 100036 439724 100037 439788
rect 99971 439723 100037 439724
rect 99234 424894 99854 438000
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99051 398036 99117 398037
rect 99051 397972 99052 398036
rect 99116 397972 99117 398036
rect 99051 397971 99117 397972
rect 99234 388894 99854 424338
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 388000 99854 388338
rect 102954 428614 103574 464058
rect 103654 460950 103714 538051
rect 104942 479773 105002 567150
rect 107699 563140 107765 563141
rect 107699 563076 107700 563140
rect 107764 563076 107765 563140
rect 107699 563075 107765 563076
rect 107515 540020 107581 540021
rect 107515 539956 107516 540020
rect 107580 539956 107581 540020
rect 107515 539955 107581 539956
rect 104939 479772 105005 479773
rect 104939 479708 104940 479772
rect 105004 479708 105005 479772
rect 104939 479707 105005 479708
rect 106779 476236 106845 476237
rect 106779 476172 106780 476236
rect 106844 476172 106845 476236
rect 106779 476171 106845 476172
rect 103654 460890 103898 460950
rect 103838 445773 103898 460890
rect 103835 445772 103901 445773
rect 103835 445708 103836 445772
rect 103900 445708 103901 445772
rect 103835 445707 103901 445708
rect 103838 444413 103898 445707
rect 103835 444412 103901 444413
rect 103835 444348 103836 444412
rect 103900 444348 103901 444412
rect 103835 444347 103901 444348
rect 106782 437477 106842 476171
rect 107518 449445 107578 539955
rect 107702 470661 107762 563075
rect 107886 535397 107946 576675
rect 109794 543454 110414 578898
rect 111566 554029 111626 643179
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 114507 586532 114573 586533
rect 114507 586468 114508 586532
rect 114572 586468 114573 586532
rect 114507 586467 114573 586468
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 111747 577420 111813 577421
rect 111747 577356 111748 577420
rect 111812 577356 111813 577420
rect 111747 577355 111813 577356
rect 111563 554028 111629 554029
rect 111563 553964 111564 554028
rect 111628 553964 111629 554028
rect 111563 553963 111629 553964
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109539 541108 109605 541109
rect 109539 541044 109540 541108
rect 109604 541044 109605 541108
rect 109539 541043 109605 541044
rect 109542 537981 109602 541043
rect 109539 537980 109605 537981
rect 109539 537916 109540 537980
rect 109604 537916 109605 537980
rect 109539 537915 109605 537916
rect 107883 535396 107949 535397
rect 107883 535332 107884 535396
rect 107948 535332 107949 535396
rect 107883 535331 107949 535332
rect 108803 534716 108869 534717
rect 108803 534652 108804 534716
rect 108868 534652 108869 534716
rect 108803 534651 108869 534652
rect 108806 534090 108866 534651
rect 108806 534030 109050 534090
rect 108990 495450 109050 534030
rect 108806 495390 109050 495450
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 108806 485790 108866 495390
rect 108806 485730 109050 485790
rect 108990 476237 109050 485730
rect 108987 476236 109053 476237
rect 108987 476172 108988 476236
rect 109052 476172 109053 476236
rect 108987 476171 109053 476172
rect 109794 471454 110414 506898
rect 110643 499628 110709 499629
rect 110643 499564 110644 499628
rect 110708 499564 110709 499628
rect 110643 499563 110709 499564
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 107699 470660 107765 470661
rect 107699 470596 107700 470660
rect 107764 470596 107765 470660
rect 107699 470595 107765 470596
rect 107515 449444 107581 449445
rect 107515 449380 107516 449444
rect 107580 449380 107581 449444
rect 107515 449379 107581 449380
rect 106779 437476 106845 437477
rect 106779 437412 106780 437476
rect 106844 437412 106845 437476
rect 106779 437411 106845 437412
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 392614 103574 428058
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 388000 103574 392058
rect 109794 435454 110414 470898
rect 110646 442373 110706 499563
rect 111011 491876 111077 491877
rect 111011 491812 111012 491876
rect 111076 491812 111077 491876
rect 111011 491811 111077 491812
rect 110643 442372 110709 442373
rect 110643 442308 110644 442372
rect 110708 442308 110709 442372
rect 110643 442307 110709 442308
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 388000 110414 398898
rect 111014 390693 111074 491811
rect 111750 485757 111810 577355
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 111931 500172 111997 500173
rect 111931 500108 111932 500172
rect 111996 500108 111997 500172
rect 111931 500107 111997 500108
rect 111747 485756 111813 485757
rect 111747 485692 111748 485756
rect 111812 485692 111813 485756
rect 111747 485691 111813 485692
rect 111934 439517 111994 500107
rect 113514 475174 114134 510618
rect 114510 500445 114570 586467
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 118003 580004 118069 580005
rect 118003 579940 118004 580004
rect 118068 579940 118069 580004
rect 118003 579939 118069 579940
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 114507 500444 114573 500445
rect 114507 500380 114508 500444
rect 114572 500380 114573 500444
rect 114507 500379 114573 500380
rect 114507 500308 114573 500309
rect 114507 500244 114508 500308
rect 114572 500244 114573 500308
rect 114507 500243 114573 500244
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 111931 439516 111997 439517
rect 111931 439452 111932 439516
rect 111996 439452 111997 439516
rect 111931 439451 111997 439452
rect 113514 439174 114134 474618
rect 114510 443733 114570 500243
rect 115059 491196 115125 491197
rect 115059 491132 115060 491196
rect 115124 491132 115125 491196
rect 115059 491131 115125 491132
rect 114507 443732 114573 443733
rect 114507 443668 114508 443732
rect 114572 443668 114573 443732
rect 114507 443667 114573 443668
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 111011 390692 111077 390693
rect 111011 390628 111012 390692
rect 111076 390628 111077 390692
rect 111011 390627 111077 390628
rect 113514 388000 114134 402618
rect 115062 400213 115122 491131
rect 117083 481540 117149 481541
rect 117083 481476 117084 481540
rect 117148 481476 117149 481540
rect 117083 481475 117149 481476
rect 115059 400212 115125 400213
rect 115059 400148 115060 400212
rect 115124 400148 115125 400212
rect 115059 400147 115125 400148
rect 115795 385252 115861 385253
rect 115795 385188 115796 385252
rect 115860 385188 115861 385252
rect 115795 385187 115861 385188
rect 115798 384573 115858 385187
rect 115795 384572 115861 384573
rect 115795 384508 115796 384572
rect 115860 384508 115861 384572
rect 115795 384507 115861 384508
rect 89568 381454 89888 381486
rect 89568 381218 89610 381454
rect 89846 381218 89888 381454
rect 89568 381134 89888 381218
rect 89568 380898 89610 381134
rect 89846 380898 89888 381134
rect 89568 380866 89888 380898
rect 70044 377710 70410 377770
rect 70044 377708 70045 377710
rect 69979 377707 70045 377708
rect 117086 376821 117146 481475
rect 117234 478894 117854 514338
rect 118006 489157 118066 579939
rect 120954 554614 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 121683 572796 121749 572797
rect 121683 572732 121684 572796
rect 121748 572732 121749 572796
rect 121683 572731 121749 572732
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 118003 489156 118069 489157
rect 118003 489092 118004 489156
rect 118068 489092 118069 489156
rect 118003 489091 118069 489092
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 388000 117854 406338
rect 117819 386340 117885 386341
rect 117819 386276 117820 386340
rect 117884 386276 117885 386340
rect 117819 386275 117885 386276
rect 117083 376820 117149 376821
rect 117083 376756 117084 376820
rect 117148 376756 117149 376820
rect 117083 376755 117149 376756
rect 117822 372741 117882 386275
rect 118006 384981 118066 489091
rect 118739 488612 118805 488613
rect 118739 488548 118740 488612
rect 118804 488548 118805 488612
rect 118739 488547 118805 488548
rect 118742 389877 118802 488547
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 121686 481541 121746 572731
rect 127794 561454 128414 596898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 129779 570348 129845 570349
rect 129779 570284 129780 570348
rect 129844 570284 129845 570348
rect 129779 570283 129845 570284
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 125731 545732 125797 545733
rect 125731 545668 125732 545732
rect 125796 545668 125797 545732
rect 125731 545667 125797 545668
rect 123339 485756 123405 485757
rect 123339 485692 123340 485756
rect 123404 485692 123405 485756
rect 123339 485691 123405 485692
rect 123342 483309 123402 485691
rect 123339 483308 123405 483309
rect 123339 483244 123340 483308
rect 123404 483244 123405 483308
rect 123339 483243 123405 483244
rect 121683 481540 121749 481541
rect 121683 481476 121684 481540
rect 121748 481476 121749 481540
rect 121683 481475 121749 481476
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 118739 389876 118805 389877
rect 118739 389812 118740 389876
rect 118804 389812 118805 389876
rect 118739 389811 118805 389812
rect 119291 387972 119357 387973
rect 119291 387908 119292 387972
rect 119356 387908 119357 387972
rect 119291 387907 119357 387908
rect 118003 384980 118069 384981
rect 118003 384916 118004 384980
rect 118068 384916 118069 384980
rect 118003 384915 118069 384916
rect 117819 372740 117885 372741
rect 117819 372676 117820 372740
rect 117884 372676 117885 372740
rect 117819 372675 117885 372676
rect 69059 370564 69125 370565
rect 69059 370500 69060 370564
rect 69124 370500 69125 370564
rect 69059 370499 69125 370500
rect 119294 369069 119354 387907
rect 119475 387836 119541 387837
rect 119475 387772 119476 387836
rect 119540 387772 119541 387836
rect 119475 387771 119541 387772
rect 119478 370565 119538 387771
rect 120027 387020 120093 387021
rect 120027 386956 120028 387020
rect 120092 386956 120093 387020
rect 120027 386955 120093 386956
rect 119475 370564 119541 370565
rect 119475 370500 119476 370564
rect 119540 370500 119541 370564
rect 119475 370499 119541 370500
rect 119291 369068 119357 369069
rect 119291 369004 119292 369068
rect 119356 369004 119357 369068
rect 119291 369003 119357 369004
rect 68875 366076 68941 366077
rect 68875 366012 68876 366076
rect 68940 366012 68941 366076
rect 68875 366011 68941 366012
rect 68139 357508 68205 357509
rect 68139 357444 68140 357508
rect 68204 357444 68205 357508
rect 68139 357443 68205 357444
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 68878 330445 68938 366011
rect 118923 364852 118989 364853
rect 118923 364788 118924 364852
rect 118988 364788 118989 364852
rect 118923 364787 118989 364788
rect 74208 363454 74528 363486
rect 74208 363218 74250 363454
rect 74486 363218 74528 363454
rect 74208 363134 74528 363218
rect 74208 362898 74250 363134
rect 74486 362898 74528 363134
rect 74208 362866 74528 362898
rect 104928 363454 105248 363486
rect 104928 363218 104970 363454
rect 105206 363218 105248 363454
rect 104928 363134 105248 363218
rect 104928 362898 104970 363134
rect 105206 362898 105248 363134
rect 104928 362866 105248 362898
rect 89568 345454 89888 345486
rect 89568 345218 89610 345454
rect 89846 345218 89888 345454
rect 89568 345134 89888 345218
rect 89568 344898 89610 345134
rect 89846 344898 89888 345134
rect 89568 344866 89888 344898
rect 70531 341052 70597 341053
rect 70531 340988 70532 341052
rect 70596 340988 70597 341052
rect 70531 340987 70597 340988
rect 70534 336021 70594 340987
rect 70531 336020 70597 336021
rect 70531 335956 70532 336020
rect 70596 335956 70597 336020
rect 70531 335955 70597 335956
rect 68875 330444 68941 330445
rect 68875 330380 68876 330444
rect 68940 330380 68941 330444
rect 68875 330379 68941 330380
rect 70899 327724 70965 327725
rect 70899 327660 70900 327724
rect 70964 327660 70965 327724
rect 70899 327659 70965 327660
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66115 298756 66181 298757
rect 66115 298692 66116 298756
rect 66180 298692 66181 298756
rect 66115 298691 66181 298692
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 66954 284614 67574 320058
rect 70902 287070 70962 327659
rect 73794 327454 74414 338000
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 294000 74414 326898
rect 77514 331174 78134 338000
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 294000 78134 294618
rect 81234 334894 81854 338000
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 294000 81854 298338
rect 84954 302614 85574 338000
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 294000 85574 302058
rect 91794 309454 92414 338000
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 95514 313174 96134 338000
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 294000 96134 312618
rect 99234 316894 99854 338000
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 294000 99854 316338
rect 102954 320614 103574 338000
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 294000 103574 320058
rect 109794 327454 110414 338000
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 113514 331174 114134 338000
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 294000 114134 294618
rect 117234 334894 117854 338000
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 118739 315348 118805 315349
rect 118739 315284 118740 315348
rect 118804 315284 118805 315348
rect 118739 315283 118805 315284
rect 118742 306390 118802 315283
rect 118926 307733 118986 364787
rect 120030 338061 120090 386955
rect 120954 374614 121574 410058
rect 122603 386612 122669 386613
rect 122603 386548 122604 386612
rect 122668 386548 122669 386612
rect 122603 386547 122669 386548
rect 122051 382260 122117 382261
rect 122051 382196 122052 382260
rect 122116 382196 122117 382260
rect 122051 382195 122117 382196
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 122054 368389 122114 382195
rect 122051 368388 122117 368389
rect 122051 368324 122052 368388
rect 122116 368324 122117 368388
rect 122051 368323 122117 368324
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120027 338060 120093 338061
rect 120027 337996 120028 338060
rect 120092 337996 120093 338060
rect 120027 337995 120093 337996
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 118923 307732 118989 307733
rect 118923 307668 118924 307732
rect 118988 307668 118989 307732
rect 118923 307667 118989 307668
rect 118742 306330 119354 306390
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 294000 117854 298338
rect 119294 289509 119354 306330
rect 120954 302614 121574 338058
rect 122606 314261 122666 386547
rect 123342 378997 123402 483243
rect 125734 453389 125794 545667
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 129782 477461 129842 570283
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 129779 477460 129845 477461
rect 129779 477396 129780 477460
rect 129844 477396 129845 477460
rect 129779 477395 129845 477396
rect 125731 453388 125797 453389
rect 125731 453324 125732 453388
rect 125796 453324 125797 453388
rect 125731 453323 125797 453324
rect 125734 451290 125794 453323
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 125734 451230 126162 451290
rect 124811 438972 124877 438973
rect 124811 438908 124812 438972
rect 124876 438908 124877 438972
rect 124811 438907 124877 438908
rect 123339 378996 123405 378997
rect 123339 378932 123340 378996
rect 123404 378932 123405 378996
rect 123339 378931 123405 378932
rect 123339 372740 123405 372741
rect 123339 372676 123340 372740
rect 123404 372676 123405 372740
rect 123339 372675 123405 372676
rect 123342 349757 123402 372675
rect 123339 349756 123405 349757
rect 123339 349692 123340 349756
rect 123404 349692 123405 349756
rect 123339 349691 123405 349692
rect 124814 316029 124874 438907
rect 126102 342413 126162 451230
rect 127794 417454 128414 452898
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 128675 444956 128741 444957
rect 128675 444892 128676 444956
rect 128740 444892 128741 444956
rect 128675 444891 128741 444892
rect 128678 431970 128738 444891
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 128494 431910 128738 431970
rect 128494 364350 128554 431910
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 129779 380220 129845 380221
rect 129779 380156 129780 380220
rect 129844 380156 129845 380220
rect 129779 380155 129845 380156
rect 128494 364290 128738 364350
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 126099 342412 126165 342413
rect 126099 342348 126100 342412
rect 126164 342348 126165 342412
rect 126099 342347 126165 342348
rect 124811 316028 124877 316029
rect 124811 315964 124812 316028
rect 124876 315964 124877 316028
rect 124811 315963 124877 315964
rect 124814 314805 124874 315963
rect 124811 314804 124877 314805
rect 124811 314740 124812 314804
rect 124876 314740 124877 314804
rect 124811 314739 124877 314740
rect 125731 314804 125797 314805
rect 125731 314740 125732 314804
rect 125796 314740 125797 314804
rect 125731 314739 125797 314740
rect 122603 314260 122669 314261
rect 122603 314196 122604 314260
rect 122668 314196 122669 314260
rect 122603 314195 122669 314196
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 294000 121574 302058
rect 122603 301476 122669 301477
rect 122603 301412 122604 301476
rect 122668 301412 122669 301476
rect 122603 301411 122669 301412
rect 121683 295628 121749 295629
rect 121683 295564 121684 295628
rect 121748 295564 121749 295628
rect 121683 295563 121749 295564
rect 119291 289508 119357 289509
rect 119291 289444 119292 289508
rect 119356 289444 119357 289508
rect 119291 289443 119357 289444
rect 70534 287010 70962 287070
rect 70534 285429 70594 287010
rect 70531 285428 70597 285429
rect 70531 285364 70532 285428
rect 70596 285364 70597 285428
rect 70531 285363 70597 285364
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 121686 284341 121746 295563
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 121683 284340 121749 284341
rect 121683 284276 121684 284340
rect 121748 284276 121749 284340
rect 121683 284275 121749 284276
rect 66954 248614 67574 284058
rect 69059 279716 69125 279717
rect 69059 279652 69060 279716
rect 69124 279652 69125 279716
rect 69059 279651 69125 279652
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 69062 232525 69122 279651
rect 89568 273454 89888 273486
rect 89568 273218 89610 273454
rect 89846 273218 89888 273454
rect 89568 273134 89888 273218
rect 89568 272898 89610 273134
rect 89846 272898 89888 273134
rect 89568 272866 89888 272898
rect 69243 257276 69309 257277
rect 69243 257212 69244 257276
rect 69308 257212 69309 257276
rect 69243 257211 69309 257212
rect 69059 232524 69125 232525
rect 69059 232460 69060 232524
rect 69124 232460 69125 232524
rect 69059 232459 69125 232460
rect 69246 225589 69306 257211
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 122606 249661 122666 301411
rect 125734 255373 125794 314739
rect 127794 309454 128414 344898
rect 128678 339421 128738 364290
rect 128675 339420 128741 339421
rect 128675 339356 128676 339420
rect 128740 339356 128741 339420
rect 128675 339355 128741 339356
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 125731 255372 125797 255373
rect 125731 255308 125732 255372
rect 125796 255308 125797 255372
rect 125731 255307 125797 255308
rect 122603 249660 122669 249661
rect 122603 249596 122604 249660
rect 122668 249596 122669 249660
rect 122603 249595 122669 249596
rect 122606 248430 122666 249595
rect 122606 248370 122850 248430
rect 122790 248301 122850 248370
rect 122787 248300 122853 248301
rect 122787 248236 122788 248300
rect 122852 248236 122853 248300
rect 122787 248235 122853 248236
rect 119291 241228 119357 241229
rect 119291 241164 119292 241228
rect 119356 241164 119357 241228
rect 119291 241163 119357 241164
rect 70531 240276 70597 240277
rect 70531 240212 70532 240276
rect 70596 240212 70597 240276
rect 70531 240211 70597 240212
rect 70534 237965 70594 240211
rect 70531 237964 70597 237965
rect 70531 237900 70532 237964
rect 70596 237900 70597 237964
rect 70531 237899 70597 237900
rect 69243 225588 69309 225589
rect 69243 225524 69244 225588
rect 69308 225524 69309 225588
rect 69243 225523 69309 225524
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 223174 78134 238000
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 238000
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 230614 85574 238000
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 238000
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 238000
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177716 97093 177717
rect 97027 177652 97028 177716
rect 97092 177652 97093 177716
rect 97027 177651 97093 177652
rect 97030 175130 97090 177651
rect 99234 176600 99854 208338
rect 102954 212614 103574 238000
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177716 100773 177717
rect 100707 177652 100708 177716
rect 100772 177652 100773 177716
rect 100707 177651 100773 177652
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 98315 175540 98381 175541
rect 98315 175476 98316 175540
rect 98380 175476 98381 175540
rect 98315 175475 98381 175476
rect 96960 175070 97090 175130
rect 98318 175130 98378 175475
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177651
rect 101995 176900 102061 176901
rect 101995 176836 101996 176900
rect 102060 176836 102061 176900
rect 101995 176835 102061 176836
rect 101998 175130 102058 176835
rect 102954 176600 103574 212058
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 105675 177716 105741 177717
rect 105675 177652 105676 177716
rect 105740 177652 105741 177716
rect 105675 177651 105741 177652
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104571 175540 104637 175541
rect 104571 175476 104572 175540
rect 104636 175476 104637 175540
rect 104571 175475 104637 175476
rect 104574 175130 104634 175475
rect 105678 175130 105738 177651
rect 108067 177036 108133 177037
rect 108067 176972 108068 177036
rect 108132 176972 108133 177036
rect 108067 176971 108133 176972
rect 106963 176764 107029 176765
rect 106963 176700 106964 176764
rect 107028 176700 107029 176764
rect 106963 176699 107029 176700
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176699
rect 108070 175130 108130 176971
rect 109539 176764 109605 176765
rect 109539 176700 109540 176764
rect 109604 176700 109605 176764
rect 109539 176699 109605 176700
rect 109542 175130 109602 176699
rect 109794 176600 110414 182898
rect 113514 223174 114134 238000
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 112115 177988 112181 177989
rect 112115 177924 112116 177988
rect 112180 177924 112181 177988
rect 112115 177923 112181 177924
rect 110643 177716 110709 177717
rect 110643 177652 110644 177716
rect 110708 177652 110709 177716
rect 110643 177651 110709 177652
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177651
rect 112118 175130 112178 177923
rect 113219 177036 113285 177037
rect 113219 176972 113220 177036
rect 113284 176972 113285 177036
rect 113219 176971 113285 176972
rect 113222 175130 113282 176971
rect 113514 176600 114134 186618
rect 117234 226894 117854 238000
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 119294 219450 119354 241163
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 114323 177716 114389 177717
rect 114323 177652 114324 177716
rect 114388 177652 114389 177716
rect 114323 177651 114389 177652
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 177651
rect 115795 177036 115861 177037
rect 115795 176972 115796 177036
rect 115860 176972 115861 177036
rect 115795 176971 115861 176972
rect 115798 175130 115858 176971
rect 117234 176600 117854 190338
rect 118742 219390 119354 219450
rect 120954 230614 121574 238000
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 118742 181389 118802 219390
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 118739 181388 118805 181389
rect 118739 181324 118740 181388
rect 118804 181324 118805 181388
rect 118739 181323 118805 181324
rect 118371 177716 118437 177717
rect 118371 177652 118372 177716
rect 118436 177652 118437 177716
rect 118371 177651 118437 177652
rect 120763 177716 120829 177717
rect 120763 177652 120764 177716
rect 120828 177652 120829 177716
rect 120763 177651 120829 177652
rect 116899 175540 116965 175541
rect 116899 175476 116900 175540
rect 116964 175476 116965 175540
rect 116899 175475 116965 175476
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 175475
rect 118374 175130 118434 177651
rect 119475 176764 119541 176765
rect 119475 176700 119476 176764
rect 119540 176700 119541 176764
rect 119475 176699 119541 176700
rect 119478 175130 119538 176699
rect 120766 175130 120826 177651
rect 120954 176600 121574 194058
rect 127794 237454 128414 272898
rect 129782 241637 129842 380155
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 129779 241636 129845 241637
rect 129779 241572 129780 241636
rect 129844 241572 129845 241636
rect 129779 241571 129845 241572
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 125731 177716 125797 177717
rect 125731 177652 125732 177716
rect 125796 177652 125797 177716
rect 125731 177651 125797 177652
rect 123155 177172 123221 177173
rect 123155 177108 123156 177172
rect 123220 177108 123221 177172
rect 123155 177107 123221 177108
rect 121867 176764 121933 176765
rect 121867 176700 121868 176764
rect 121932 176700 121933 176764
rect 121867 176699 121933 176700
rect 121870 175130 121930 176699
rect 123158 175130 123218 177107
rect 124443 176764 124509 176765
rect 124443 176700 124444 176764
rect 124508 176700 124509 176764
rect 124443 176699 124509 176700
rect 124446 175130 124506 176699
rect 125734 175130 125794 177651
rect 127019 176764 127085 176765
rect 127019 176700 127020 176764
rect 127084 176700 127085 176764
rect 127019 176699 127085 176700
rect 127022 175130 127082 176699
rect 127794 176600 128414 200898
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 130699 177716 130765 177717
rect 130699 177652 130700 177716
rect 130764 177652 130765 177716
rect 130699 177651 130765 177652
rect 128123 175540 128189 175541
rect 128123 175476 128124 175540
rect 128188 175476 128189 175540
rect 128123 175475 128189 175476
rect 129411 175540 129477 175541
rect 129411 175476 129412 175540
rect 129476 175476 129477 175540
rect 129411 175475 129477 175476
rect 128126 175130 128186 175475
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 175475
rect 130702 175130 130762 177651
rect 131514 176600 132134 204618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 136587 498812 136653 498813
rect 136587 498748 136588 498812
rect 136652 498748 136653 498812
rect 136587 498747 136653 498748
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 136590 390557 136650 498747
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 136587 390556 136653 390557
rect 136587 390492 136588 390556
rect 136652 390492 136653 390556
rect 136587 390491 136653 390492
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177716 132421 177717
rect 132355 177652 132356 177716
rect 132420 177652 132421 177716
rect 132355 177651 132421 177652
rect 132358 175130 132418 177651
rect 133091 176764 133157 176765
rect 133091 176700 133092 176764
rect 133156 176700 133157 176764
rect 133091 176699 133157 176700
rect 134379 176764 134445 176765
rect 134379 176700 134380 176764
rect 134444 176700 134445 176764
rect 134379 176699 134445 176700
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 176699
rect 134382 175130 134442 176699
rect 135234 176600 135854 208338
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 176600 150134 186618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 176600 164414 200898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 166211 178124 166277 178125
rect 166211 178060 166212 178124
rect 166276 178060 166277 178124
rect 166211 178059 166277 178060
rect 148179 175540 148245 175541
rect 148179 175476 148180 175540
rect 148244 175476 148245 175540
rect 148179 175475 148245 175476
rect 158851 175540 158917 175541
rect 158851 175476 158852 175540
rect 158916 175476 158917 175540
rect 158851 175475 158917 175476
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 175475
rect 158854 175130 158914 175475
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 166214 162893 166274 178059
rect 167514 169174 168134 204618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 173019 330580 173085 330581
rect 173019 330516 173020 330580
rect 173084 330516 173085 330580
rect 173019 330515 173085 330516
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 168235 176900 168301 176901
rect 168235 176836 168236 176900
rect 168300 176836 168301 176900
rect 168235 176835 168301 176836
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 166211 162892 166277 162893
rect 166211 162828 166212 162892
rect 166276 162828 166277 162892
rect 166211 162827 166277 162828
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 167514 133174 168134 168618
rect 168238 160717 168298 176835
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 168235 160716 168301 160717
rect 168235 160652 168236 160716
rect 168300 160652 168301 160716
rect 168235 160651 168301 160652
rect 168235 145076 168301 145077
rect 168235 145012 168236 145076
rect 168300 145012 168301 145076
rect 168235 145011 168301 145012
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 166211 132836 166277 132837
rect 166211 132772 166212 132836
rect 166276 132772 166277 132836
rect 166211 132771 166277 132772
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 62987 69596 63053 69597
rect 62987 69532 62988 69596
rect 63052 69532 63053 69596
rect 62987 69531 63053 69532
rect 63234 64894 63854 100338
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 61883 10980 61949 10981
rect 61883 10916 61884 10980
rect 61948 10916 61949 10980
rect 61883 10915 61949 10916
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 92445 74826 94830
rect 74763 92444 74829 92445
rect 74763 92380 74764 92444
rect 74828 92380 74829 92444
rect 74763 92379 74829 92380
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 91221 84394 94830
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 92445 85866 94830
rect 85803 92444 85869 92445
rect 85803 92380 85804 92444
rect 85868 92380 85869 92444
rect 85803 92379 85869 92380
rect 86726 91221 86786 94830
rect 88014 92445 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 92445 88994 94830
rect 88011 92444 88077 92445
rect 88011 92380 88012 92444
rect 88076 92380 88077 92444
rect 88011 92379 88077 92380
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 90222 91765 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96170 94890
rect 90219 91764 90285 91765
rect 90219 91700 90220 91764
rect 90284 91700 90285 91764
rect 90219 91699 90285 91700
rect 91326 91221 91386 94830
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91357 93962 94830
rect 93899 91356 93965 91357
rect 93899 91292 93900 91356
rect 93964 91292 93965 91356
rect 93899 91291 93965 91292
rect 95006 91221 95066 94830
rect 96110 93941 96170 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96107 93940 96173 93941
rect 96107 93876 96108 93940
rect 96172 93876 96173 93940
rect 96107 93875 96173 93876
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96662 91221 96722 94830
rect 97214 92445 97274 94830
rect 97211 92444 97277 92445
rect 97211 92380 97212 92444
rect 97276 92380 97277 92444
rect 97211 92379 97277 92380
rect 98134 91357 98194 94830
rect 98502 92445 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 98499 92444 98565 92445
rect 98499 92380 98500 92444
rect 98564 92380 98565 92444
rect 98499 92379 98565 92380
rect 98131 91356 98197 91357
rect 98131 91292 98132 91356
rect 98196 91292 98197 91356
rect 98131 91291 98197 91292
rect 99054 91221 99114 94830
rect 96659 91220 96725 91221
rect 96659 91156 96660 91220
rect 96724 91156 96725 91220
rect 96659 91155 96725 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 91221 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 100526 91357 100586 94830
rect 100894 93533 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 100891 93532 100957 93533
rect 100891 93468 100892 93532
rect 100956 93468 100957 93532
rect 100891 93467 100957 93468
rect 101814 91357 101874 94830
rect 100523 91356 100589 91357
rect 100523 91292 100524 91356
rect 100588 91292 100589 91356
rect 100523 91291 100589 91292
rect 101811 91356 101877 91357
rect 101811 91292 101812 91356
rect 101876 91292 101877 91356
rect 101811 91291 101877 91292
rect 101998 91221 102058 94830
rect 102918 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 102918 93870 102978 94830
rect 102734 93810 102978 93870
rect 102734 92309 102794 93810
rect 103286 93261 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 103283 93260 103349 93261
rect 103283 93196 103284 93260
rect 103348 93196 103349 93260
rect 103283 93195 103349 93196
rect 102731 92308 102797 92309
rect 102731 92244 102732 92308
rect 102796 92244 102797 92308
rect 102731 92243 102797 92244
rect 99971 91220 100037 91221
rect 99971 91156 99972 91220
rect 100036 91156 100037 91220
rect 99971 91155 100037 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91221 104266 94830
rect 104574 91221 104634 94830
rect 105494 91357 105554 94830
rect 105491 91356 105557 91357
rect 105491 91292 105492 91356
rect 105556 91292 105557 91356
rect 105491 91291 105557 91292
rect 105678 91221 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 106414 91357 106474 94830
rect 106411 91356 106477 91357
rect 106411 91292 106412 91356
rect 106476 91292 106477 91356
rect 106411 91291 106477 91292
rect 106782 91221 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 107702 91221 107762 94830
rect 108070 91221 108130 94830
rect 109174 93533 109234 94830
rect 109171 93532 109237 93533
rect 109171 93468 109172 93532
rect 109236 93468 109237 93532
rect 109171 93467 109237 93468
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105675 91220 105741 91221
rect 105675 91156 105676 91220
rect 105740 91156 105741 91220
rect 105675 91155 105741 91156
rect 106779 91220 106845 91221
rect 106779 91156 106780 91220
rect 106844 91156 106845 91220
rect 106779 91155 106845 91156
rect 107699 91220 107765 91221
rect 107699 91156 107700 91220
rect 107764 91156 107765 91220
rect 107699 91155 107765 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 91221 111258 94830
rect 111934 91221 111994 94830
rect 112302 94830 112388 94890
rect 113038 94830 113204 94890
rect 113406 94830 113748 94890
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 112302 94077 112362 94830
rect 112299 94076 112365 94077
rect 112299 94012 112300 94076
rect 112364 94012 112365 94076
rect 112299 94011 112365 94012
rect 113038 92445 113098 94830
rect 113406 93870 113466 94830
rect 113222 93810 113466 93870
rect 113035 92444 113101 92445
rect 113035 92380 113036 92444
rect 113100 92380 113101 92444
rect 113035 92379 113101 92380
rect 113222 91221 113282 93810
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 113219 91220 113285 91221
rect 113219 91156 113220 91220
rect 113284 91156 113285 91220
rect 113219 91155 113285 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 94830
rect 114878 92445 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 92445 115490 94830
rect 114875 92444 114941 92445
rect 114875 92380 114876 92444
rect 114940 92380 114941 92444
rect 114875 92379 114941 92380
rect 115427 92444 115493 92445
rect 115427 92380 115428 92444
rect 115492 92380 115493 92444
rect 115427 92379 115493 92380
rect 115798 91221 115858 94830
rect 116718 93533 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 93532 116781 93533
rect 116715 93468 116716 93532
rect 116780 93468 116781 93532
rect 116715 93467 116781 93468
rect 117086 91221 117146 94830
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 92445 118066 94830
rect 118003 92444 118069 92445
rect 118003 92380 118004 92444
rect 118068 92380 118069 92444
rect 118003 92379 118069 92380
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119294 91629 119354 94830
rect 119291 91628 119357 91629
rect 119291 91564 119292 91628
rect 119356 91564 119357 91628
rect 119291 91563 119357 91564
rect 119662 91221 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 120214 91221 120274 94830
rect 120582 91357 120642 94830
rect 121686 93533 121746 94830
rect 121683 93532 121749 93533
rect 121683 93468 121684 93532
rect 121748 93468 121749 93532
rect 121683 93467 121749 93468
rect 120579 91356 120645 91357
rect 120579 91292 120580 91356
rect 120644 91292 120645 91356
rect 120579 91291 120645 91292
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 119659 91220 119725 91221
rect 119659 91156 119660 91220
rect 119724 91156 119725 91220
rect 119659 91155 119725 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 122054 92309 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122051 92308 122117 92309
rect 122051 92244 122052 92308
rect 122116 92244 122117 92308
rect 122051 92243 122117 92244
rect 122606 92170 122666 93810
rect 122787 92172 122853 92173
rect 122787 92170 122788 92172
rect 122606 92110 122788 92170
rect 122787 92108 122788 92110
rect 122852 92108 122853 92172
rect 122787 92107 122853 92108
rect 123158 91221 123218 94830
rect 124078 91357 124138 94830
rect 124446 91357 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 124075 91356 124141 91357
rect 124075 91292 124076 91356
rect 124140 91292 124141 91356
rect 124075 91291 124141 91292
rect 124443 91356 124509 91357
rect 124443 91292 124444 91356
rect 124508 91292 124509 91356
rect 124443 91291 124509 91292
rect 125366 91221 125426 94830
rect 125734 91221 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 126470 94213 126530 94830
rect 126467 94212 126533 94213
rect 126467 94148 126468 94212
rect 126532 94148 126533 94212
rect 126467 94147 126533 94148
rect 126654 94077 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 126651 94076 126717 94077
rect 126651 94012 126652 94076
rect 126716 94012 126717 94076
rect 126651 94011 126717 94012
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 125731 91220 125797 91221
rect 125731 91156 125732 91220
rect 125796 91156 125797 91220
rect 125731 91155 125797 91156
rect 127574 90949 127634 94830
rect 127571 90948 127637 90949
rect 127571 90884 127572 90948
rect 127636 90884 127637 90948
rect 127571 90883 127637 90884
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 91221 130762 94830
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 92445 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133094 93533 133154 94830
rect 133091 93532 133157 93533
rect 133091 93468 133092 93532
rect 133156 93468 133157 93532
rect 133091 93467 133157 93468
rect 132355 92444 132421 92445
rect 132355 92380 132356 92444
rect 132420 92380 132421 92444
rect 132355 92379 132421 92380
rect 134382 91221 134442 94830
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 91629 136098 94830
rect 151310 94830 151556 94890
rect 136035 91628 136101 91629
rect 136035 91564 136036 91628
rect 136100 91564 136101 91628
rect 136035 91563 136101 91564
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 92173 151370 94830
rect 151491 94620 151557 94621
rect 151491 94556 151492 94620
rect 151556 94556 151557 94620
rect 151491 94555 151557 94556
rect 151494 92445 151554 94555
rect 151632 94210 151692 95200
rect 151768 94621 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151765 94620 151831 94621
rect 151765 94556 151766 94620
rect 151830 94556 151831 94620
rect 151765 94555 151831 94556
rect 152046 94213 152106 94830
rect 152043 94212 152109 94213
rect 151632 94150 151738 94210
rect 151678 93533 151738 94150
rect 152043 94148 152044 94212
rect 152108 94148 152109 94212
rect 152043 94147 152109 94148
rect 151675 93532 151741 93533
rect 151675 93468 151676 93532
rect 151740 93468 151741 93532
rect 151675 93467 151741 93468
rect 151491 92444 151557 92445
rect 151491 92380 151492 92444
rect 151556 92380 151557 92444
rect 151491 92379 151557 92380
rect 151307 92172 151373 92173
rect 151307 92108 151308 92172
rect 151372 92108 151373 92172
rect 151307 92107 151373 92108
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 79933 166274 132771
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 166395 127124 166461 127125
rect 166395 127060 166396 127124
rect 166460 127060 166461 127124
rect 166395 127059 166461 127060
rect 166398 82789 166458 127059
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166395 82788 166461 82789
rect 166395 82724 166396 82788
rect 166460 82724 166461 82788
rect 166395 82723 166461 82724
rect 166211 79932 166277 79933
rect 166211 79868 166212 79932
rect 166276 79868 166277 79932
rect 166211 79867 166277 79868
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 168238 85509 168298 145011
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 170443 134196 170509 134197
rect 170443 134132 170444 134196
rect 170508 134132 170509 134196
rect 170443 134131 170509 134132
rect 168971 131476 169037 131477
rect 168971 131412 168972 131476
rect 169036 131412 169037 131476
rect 168971 131411 169037 131412
rect 168235 85508 168301 85509
rect 168235 85444 168236 85508
rect 168300 85444 168301 85508
rect 168235 85443 168301 85444
rect 168974 81429 169034 131411
rect 170259 128620 170325 128621
rect 170259 128556 170260 128620
rect 170324 128556 170325 128620
rect 170259 128555 170325 128556
rect 169155 101420 169221 101421
rect 169155 101356 169156 101420
rect 169220 101356 169221 101420
rect 169155 101355 169221 101356
rect 169158 92309 169218 101355
rect 169155 92308 169221 92309
rect 169155 92244 169156 92308
rect 169220 92244 169221 92308
rect 169155 92243 169221 92244
rect 168971 81428 169037 81429
rect 168971 81364 168972 81428
rect 169036 81364 169037 81428
rect 168971 81363 169037 81364
rect 170262 80069 170322 128555
rect 170446 88229 170506 134131
rect 171234 100894 171854 136338
rect 172099 103596 172165 103597
rect 172099 103532 172100 103596
rect 172164 103532 172165 103596
rect 172099 103531 172165 103532
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 170443 88228 170509 88229
rect 170443 88164 170444 88228
rect 170508 88164 170509 88228
rect 170443 88163 170509 88164
rect 170259 80068 170325 80069
rect 170259 80004 170260 80068
rect 170324 80004 170325 80068
rect 170259 80003 170325 80004
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100338
rect 172102 84149 172162 103531
rect 172099 84148 172165 84149
rect 172099 84084 172100 84148
rect 172164 84084 172165 84148
rect 172099 84083 172165 84084
rect 173022 77893 173082 330515
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 173203 232660 173269 232661
rect 173203 232596 173204 232660
rect 173268 232596 173269 232660
rect 173203 232595 173269 232596
rect 173206 95573 173266 232595
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 173203 95572 173269 95573
rect 173203 95508 173204 95572
rect 173268 95508 173269 95572
rect 173203 95507 173269 95508
rect 173019 77892 173085 77893
rect 173019 77828 173020 77892
rect 173084 77828 173085 77892
rect 173019 77827 173085 77828
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 214419 179484 214485 179485
rect 214419 179420 214420 179484
rect 214484 179420 214485 179484
rect 214419 179419 214485 179420
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 214422 162077 214482 179419
rect 217794 178000 218414 182898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 178000 240134 204618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 178000 243854 208338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 259499 384572 259565 384573
rect 259499 384508 259500 384572
rect 259564 384508 259565 384572
rect 259499 384507 259565 384508
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 258395 333300 258461 333301
rect 258395 333236 258396 333300
rect 258460 333236 258461 333300
rect 258395 333235 258461 333236
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 255267 295492 255333 295493
rect 255267 295428 255268 295492
rect 255332 295428 255333 295492
rect 255267 295427 255333 295428
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 252507 289916 252573 289917
rect 252507 289852 252508 289916
rect 252572 289852 252573 289916
rect 252507 289851 252573 289852
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 178000 247574 212058
rect 249379 177580 249445 177581
rect 249379 177516 249380 177580
rect 249444 177516 249445 177580
rect 249379 177515 249445 177516
rect 249195 175948 249261 175949
rect 249195 175884 249196 175948
rect 249260 175884 249261 175948
rect 249195 175883 249261 175884
rect 249198 174317 249258 175883
rect 249195 174316 249261 174317
rect 249195 174252 249196 174316
rect 249260 174252 249261 174316
rect 249195 174251 249261 174252
rect 249382 173773 249442 177515
rect 249747 176628 249813 176629
rect 249747 176564 249748 176628
rect 249812 176564 249813 176628
rect 249747 176563 249813 176564
rect 249379 173772 249445 173773
rect 249379 173708 249380 173772
rect 249444 173708 249445 173772
rect 249379 173707 249445 173708
rect 227874 165454 228194 165486
rect 227874 165218 227916 165454
rect 228152 165218 228194 165454
rect 227874 165134 228194 165218
rect 227874 164898 227916 165134
rect 228152 164898 228194 165134
rect 227874 164866 228194 164898
rect 237805 165454 238125 165486
rect 237805 165218 237847 165454
rect 238083 165218 238125 165454
rect 237805 165134 238125 165218
rect 237805 164898 237847 165134
rect 238083 164898 238125 165134
rect 237805 164866 238125 164898
rect 214419 162076 214485 162077
rect 214419 162012 214420 162076
rect 214484 162012 214485 162076
rect 214419 162011 214485 162012
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 249750 137053 249810 176563
rect 252510 159221 252570 289851
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 252507 159220 252573 159221
rect 252507 159156 252508 159220
rect 252572 159156 252573 159220
rect 252507 159155 252573 159156
rect 251771 149700 251837 149701
rect 251771 149636 251772 149700
rect 251836 149636 251837 149700
rect 251771 149635 251837 149636
rect 249747 137052 249813 137053
rect 249747 136988 249748 137052
rect 249812 136988 249813 137052
rect 249747 136987 249813 136988
rect 227874 129454 228194 129486
rect 227874 129218 227916 129454
rect 228152 129218 228194 129454
rect 227874 129134 228194 129218
rect 227874 128898 227916 129134
rect 228152 128898 228194 129134
rect 227874 128866 228194 128898
rect 237805 129454 238125 129486
rect 237805 129218 237847 129454
rect 238083 129218 238125 129454
rect 237805 129134 238125 129218
rect 237805 128898 237847 129134
rect 238083 128898 238125 129134
rect 237805 128866 238125 128898
rect 251774 116925 251834 149635
rect 253794 147454 254414 182898
rect 255270 157317 255330 295427
rect 257514 295174 258134 330618
rect 258398 316050 258458 333235
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 256739 283524 256805 283525
rect 256739 283460 256740 283524
rect 256804 283460 256805 283524
rect 256739 283459 256805 283460
rect 255451 178668 255517 178669
rect 255451 178604 255452 178668
rect 255516 178604 255517 178668
rect 255451 178603 255517 178604
rect 255454 166293 255514 178603
rect 255451 166292 255517 166293
rect 255451 166228 255452 166292
rect 255516 166228 255517 166292
rect 255451 166227 255517 166228
rect 255267 157316 255333 157317
rect 255267 157252 255268 157316
rect 255332 157252 255333 157316
rect 255267 157251 255333 157252
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 251771 116924 251837 116925
rect 251771 116860 251772 116924
rect 251836 116860 251837 116924
rect 251771 116859 251837 116860
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 253794 111454 254414 146898
rect 256742 137597 256802 283459
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 256739 137596 256805 137597
rect 256739 137532 256740 137596
rect 256804 137532 256805 137596
rect 256739 137531 256805 137532
rect 255819 123180 255885 123181
rect 255819 123116 255820 123180
rect 255884 123116 255885 123180
rect 255819 123115 255885 123116
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 252507 111076 252573 111077
rect 252507 111012 252508 111076
rect 252572 111012 252573 111076
rect 252507 111011 252573 111012
rect 242771 110866 243091 110898
rect 252510 109853 252570 111011
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 252507 109852 252573 109853
rect 252507 109788 252508 109852
rect 252572 109788 252573 109852
rect 252507 109787 252573 109788
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214419 102508 214485 102509
rect 214419 102444 214420 102508
rect 214484 102444 214485 102508
rect 214419 102443 214485 102444
rect 214422 91085 214482 102443
rect 214419 91084 214485 91085
rect 214419 91020 214420 91084
rect 214484 91020 214485 91084
rect 214419 91019 214485 91020
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 94000
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 94000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 94000
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 75454 254414 110898
rect 255822 94485 255882 123115
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 255819 94484 255885 94485
rect 255819 94420 255820 94484
rect 255884 94420 255885 94484
rect 255819 94419 255885 94420
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 258214 315990 258458 316050
rect 258214 16590 258274 315990
rect 258395 180164 258461 180165
rect 258395 180100 258396 180164
rect 258460 180100 258461 180164
rect 258395 180099 258461 180100
rect 258398 153781 258458 180099
rect 258395 153780 258461 153781
rect 258395 153716 258396 153780
rect 258460 153716 258461 153780
rect 258395 153715 258461 153716
rect 259502 65653 259562 384507
rect 261234 370894 261854 406338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 262995 386476 263061 386477
rect 262995 386412 262996 386476
rect 263060 386412 263061 386476
rect 262995 386411 263061 386412
rect 262811 374644 262877 374645
rect 262811 374580 262812 374644
rect 262876 374580 262877 374644
rect 262811 374579 262877 374580
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 260051 181388 260117 181389
rect 260051 181324 260052 181388
rect 260116 181324 260117 181388
rect 260051 181323 260117 181324
rect 259499 65652 259565 65653
rect 259499 65588 259500 65652
rect 259564 65588 259565 65652
rect 259499 65587 259565 65588
rect 258214 16530 258458 16590
rect 258398 10981 258458 16530
rect 259502 11797 259562 65587
rect 260054 56541 260114 181323
rect 261234 154894 261854 190338
rect 262075 175404 262141 175405
rect 262075 175340 262076 175404
rect 262140 175340 262141 175404
rect 262075 175339 262141 175340
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 262078 97341 262138 175339
rect 262075 97340 262141 97341
rect 262075 97276 262076 97340
rect 262140 97276 262141 97340
rect 262075 97275 262141 97276
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 260051 56540 260117 56541
rect 260051 56476 260052 56540
rect 260116 56476 260117 56540
rect 260051 56475 260117 56476
rect 261234 46894 261854 82338
rect 262814 58037 262874 374579
rect 262998 82789 263058 386411
rect 264954 374614 265574 410058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 268331 389196 268397 389197
rect 268331 389132 268332 389196
rect 268396 389132 268397 389196
rect 268331 389131 268397 389132
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 263547 326364 263613 326365
rect 263547 326300 263548 326364
rect 263612 326300 263613 326364
rect 263547 326299 263613 326300
rect 262995 82788 263061 82789
rect 262995 82724 262996 82788
rect 263060 82724 263061 82788
rect 262995 82723 263061 82724
rect 262998 81565 263058 82723
rect 262995 81564 263061 81565
rect 262995 81500 262996 81564
rect 263060 81500 263061 81564
rect 262995 81499 263061 81500
rect 262811 58036 262877 58037
rect 262811 57972 262812 58036
rect 262876 57972 262877 58036
rect 262811 57971 262877 57972
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 259499 11796 259565 11797
rect 259499 11732 259500 11796
rect 259564 11732 259565 11796
rect 259499 11731 259565 11732
rect 258395 10980 258461 10981
rect 258395 10916 258396 10980
rect 258460 10916 258461 10980
rect 258395 10915 258461 10916
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 46338
rect 262814 12341 262874 57971
rect 263550 24173 263610 326299
rect 264954 302614 265574 338058
rect 266859 312492 266925 312493
rect 266859 312428 266860 312492
rect 266924 312428 266925 312492
rect 266859 312427 266925 312428
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 263731 193900 263797 193901
rect 263731 193836 263732 193900
rect 263796 193836 263797 193900
rect 263731 193835 263797 193836
rect 263734 160853 263794 193835
rect 263731 160852 263797 160853
rect 263731 160788 263732 160852
rect 263796 160788 263797 160852
rect 263731 160787 263797 160788
rect 264954 158614 265574 194058
rect 266307 180028 266373 180029
rect 266307 179964 266308 180028
rect 266372 179964 266373 180028
rect 266307 179963 266373 179964
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 266310 142221 266370 179963
rect 266307 142220 266373 142221
rect 266307 142156 266308 142220
rect 266372 142156 266373 142220
rect 266307 142155 266373 142156
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 266862 81429 266922 312427
rect 266859 81428 266925 81429
rect 266859 81364 266860 81428
rect 266924 81364 266925 81428
rect 266859 81363 266925 81364
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 263547 24172 263613 24173
rect 263547 24108 263548 24172
rect 263612 24108 263613 24172
rect 263547 24107 263613 24108
rect 262811 12340 262877 12341
rect 262811 12276 262812 12340
rect 262876 12276 262877 12340
rect 262811 12275 262877 12276
rect 263550 11797 263610 24107
rect 264954 14614 265574 50058
rect 268334 43485 268394 389131
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 270539 331804 270605 331805
rect 270539 331740 270540 331804
rect 270604 331740 270605 331804
rect 270539 331739 270605 331740
rect 269067 329084 269133 329085
rect 269067 329020 269068 329084
rect 269132 329020 269133 329084
rect 269067 329019 269133 329020
rect 269070 47565 269130 329019
rect 269619 176764 269685 176765
rect 269619 176700 269620 176764
rect 269684 176700 269685 176764
rect 269619 176699 269685 176700
rect 269622 97205 269682 176699
rect 269619 97204 269685 97205
rect 269619 97140 269620 97204
rect 269684 97140 269685 97204
rect 269619 97139 269685 97140
rect 269067 47564 269133 47565
rect 269067 47500 269068 47564
rect 269132 47500 269133 47564
rect 269067 47499 269133 47500
rect 268331 43484 268397 43485
rect 268331 43420 268332 43484
rect 268396 43420 268397 43484
rect 268331 43419 268397 43420
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 263547 11796 263613 11797
rect 263547 11732 263548 11796
rect 263612 11732 263613 11796
rect 263547 11731 263613 11732
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 269070 11797 269130 47499
rect 270542 27029 270602 331739
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 270539 27028 270605 27029
rect 270539 26964 270540 27028
rect 270604 26964 270605 27028
rect 270539 26963 270605 26964
rect 270542 12749 270602 26963
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 270539 12748 270605 12749
rect 270539 12684 270540 12748
rect 270604 12684 270605 12748
rect 270539 12683 270605 12684
rect 269067 11796 269133 11797
rect 269067 11732 269068 11796
rect 269132 11732 269133 11796
rect 269067 11731 269133 11732
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 287651 373284 287717 373285
rect 287651 373220 287652 373284
rect 287716 373220 287717 373284
rect 287651 373219 287717 373220
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 284339 69596 284405 69597
rect 284339 69532 284340 69596
rect 284404 69532 284405 69596
rect 284339 69531 284405 69532
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 284342 49061 284402 69531
rect 284339 49060 284405 49061
rect 284339 48996 284340 49060
rect 284404 48996 284405 49060
rect 284339 48995 284405 48996
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 284342 11797 284402 48995
rect 284339 11796 284405 11797
rect 284339 11732 284340 11796
rect 284404 11732 284405 11796
rect 284339 11731 284405 11732
rect 287654 9621 287714 373219
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 288939 128756 289005 128757
rect 288939 128692 288940 128756
rect 289004 128692 289005 128756
rect 288939 128691 289005 128692
rect 288942 46205 289002 128691
rect 289794 111454 290414 146898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 291699 125900 291765 125901
rect 291699 125836 291700 125900
rect 291764 125836 291765 125900
rect 291699 125835 291765 125836
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 288939 46204 289005 46205
rect 288939 46140 288940 46204
rect 289004 46140 289005 46204
rect 288939 46139 289005 46140
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 287651 9620 287717 9621
rect 287651 9556 287652 9620
rect 287716 9556 287717 9620
rect 287651 9555 287717 9556
rect 289794 3454 290414 38898
rect 291702 26893 291762 125835
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 291699 26892 291765 26893
rect 291699 26828 291700 26892
rect 291764 26828 291765 26892
rect 291699 26827 291765 26828
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 299611 387020 299677 387021
rect 299611 386956 299612 387020
rect 299676 386956 299677 387020
rect 299611 386955 299677 386956
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 298139 298756 298205 298757
rect 298139 298692 298140 298756
rect 298204 298692 298205 298756
rect 298139 298691 298205 298692
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 298142 43349 298202 298691
rect 298139 43348 298205 43349
rect 298139 43284 298140 43348
rect 298204 43284 298205 43348
rect 298139 43283 298205 43284
rect 298142 11797 298202 43283
rect 299614 39405 299674 386955
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 302187 326500 302253 326501
rect 302187 326436 302188 326500
rect 302252 326436 302253 326500
rect 302187 326435 302253 326436
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 299979 130116 300045 130117
rect 299979 130052 299980 130116
rect 300044 130052 300045 130116
rect 299979 130051 300045 130052
rect 299982 57221 300042 130051
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 299979 57220 300045 57221
rect 299979 57156 299980 57220
rect 300044 57156 300045 57220
rect 299979 57155 300045 57156
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 299611 39404 299677 39405
rect 299611 39340 299612 39404
rect 299676 39340 299677 39404
rect 299611 39339 299677 39340
rect 299614 11797 299674 39339
rect 300954 14614 301574 50058
rect 302190 40765 302250 326435
rect 307794 309454 308414 344898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 309731 322148 309797 322149
rect 309731 322084 309732 322148
rect 309796 322084 309797 322148
rect 309731 322083 309797 322084
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 178000 308414 200898
rect 307155 149836 307221 149837
rect 307155 149772 307156 149836
rect 307220 149772 307221 149836
rect 307155 149771 307221 149772
rect 306971 145076 307037 145077
rect 306971 145012 306972 145076
rect 307036 145012 307037 145076
rect 306971 145011 307037 145012
rect 306974 140045 307034 145011
rect 306971 140044 307037 140045
rect 306971 139980 306972 140044
rect 307036 139980 307037 140044
rect 306971 139979 307037 139980
rect 304211 139772 304277 139773
rect 304211 139708 304212 139772
rect 304276 139708 304277 139772
rect 304211 139707 304277 139708
rect 302739 132700 302805 132701
rect 302739 132636 302740 132700
rect 302804 132636 302805 132700
rect 302739 132635 302805 132636
rect 302742 64157 302802 132635
rect 302739 64156 302805 64157
rect 302739 64092 302740 64156
rect 302804 64092 302805 64156
rect 302739 64091 302805 64092
rect 302187 40764 302253 40765
rect 302187 40700 302188 40764
rect 302252 40700 302253 40764
rect 302187 40699 302253 40700
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 298139 11796 298205 11797
rect 298139 11732 298140 11796
rect 298204 11732 298205 11796
rect 298139 11731 298205 11732
rect 299611 11796 299677 11797
rect 299611 11732 299612 11796
rect 299676 11732 299677 11796
rect 299611 11731 299677 11732
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 302190 11797 302250 40699
rect 304214 28253 304274 139707
rect 307158 137325 307218 149771
rect 307155 137324 307221 137325
rect 307155 137260 307156 137324
rect 307220 137260 307221 137324
rect 307155 137259 307221 137260
rect 306971 137052 307037 137053
rect 306971 136988 306972 137052
rect 307036 136988 307037 137052
rect 306971 136987 307037 136988
rect 304395 113524 304461 113525
rect 304395 113460 304396 113524
rect 304460 113460 304461 113524
rect 304395 113459 304461 113460
rect 304398 76533 304458 113459
rect 306974 84829 307034 136987
rect 307155 113660 307221 113661
rect 307155 113596 307156 113660
rect 307220 113596 307221 113660
rect 307155 113595 307221 113596
rect 307158 90405 307218 113595
rect 309734 103530 309794 322083
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 178000 312134 204618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 178000 315854 208338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 322979 302292 323045 302293
rect 322979 302228 322980 302292
rect 323044 302228 323045 302292
rect 322979 302227 323045 302228
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 321507 239460 321573 239461
rect 321507 239396 321508 239460
rect 321572 239396 321573 239460
rect 321507 239395 321573 239396
rect 320219 229804 320285 229805
rect 320219 229740 320220 229804
rect 320284 229740 320285 229804
rect 320219 229739 320285 229740
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 178000 319574 212058
rect 320222 190470 320282 229739
rect 320222 190410 321386 190470
rect 321326 169557 321386 190410
rect 321323 169556 321389 169557
rect 321323 169492 321324 169556
rect 321388 169492 321389 169556
rect 321323 169491 321389 169492
rect 314208 165454 314528 165486
rect 314208 165218 314250 165454
rect 314486 165218 314528 165454
rect 314208 165134 314528 165218
rect 314208 164898 314250 165134
rect 314486 164898 314528 165134
rect 314208 164866 314528 164898
rect 317472 165454 317792 165486
rect 317472 165218 317514 165454
rect 317750 165218 317792 165454
rect 317472 165134 317792 165218
rect 317472 164898 317514 165134
rect 317750 164898 317792 165134
rect 317472 164866 317792 164898
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 321510 144941 321570 239395
rect 321507 144940 321573 144941
rect 321507 144876 321508 144940
rect 321572 144876 321573 144940
rect 321507 144875 321573 144876
rect 322982 134061 323042 302227
rect 325794 291454 326414 326898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 326659 299572 326725 299573
rect 326659 299508 326660 299572
rect 326724 299508 326725 299572
rect 326659 299507 326725 299508
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 322979 134060 323045 134061
rect 322979 133996 322980 134060
rect 323044 133996 323045 134060
rect 322979 133995 323045 133996
rect 314208 129454 314528 129486
rect 314208 129218 314250 129454
rect 314486 129218 314528 129454
rect 314208 129134 314528 129218
rect 314208 128898 314250 129134
rect 314486 128898 314528 129134
rect 314208 128866 314528 128898
rect 317472 129454 317792 129486
rect 317472 129218 317514 129454
rect 317750 129218 317792 129454
rect 317472 129134 317792 129218
rect 317472 128898 317514 129134
rect 317750 128898 317792 129134
rect 317472 128866 317792 128898
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 309366 103470 309794 103530
rect 309366 98970 309426 103470
rect 309731 101828 309797 101829
rect 309731 101764 309732 101828
rect 309796 101764 309797 101828
rect 309731 101763 309797 101764
rect 309734 101690 309794 101763
rect 309734 101630 309978 101690
rect 309366 98910 309794 98970
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307155 90404 307221 90405
rect 307155 90340 307156 90404
rect 307220 90340 307221 90404
rect 307155 90339 307221 90340
rect 306971 84828 307037 84829
rect 306971 84764 306972 84828
rect 307036 84764 307037 84828
rect 306971 84763 307037 84764
rect 304395 76532 304461 76533
rect 304395 76468 304396 76532
rect 304460 76468 304461 76532
rect 304395 76467 304461 76468
rect 307794 57454 308414 92898
rect 309734 78029 309794 98910
rect 309918 93870 309978 101630
rect 324267 99380 324333 99381
rect 324267 99316 324268 99380
rect 324332 99316 324333 99380
rect 324267 99315 324333 99316
rect 321507 98020 321573 98021
rect 321507 97956 321508 98020
rect 321572 97956 321573 98020
rect 321507 97955 321573 97956
rect 309918 93810 310162 93870
rect 310102 90405 310162 93810
rect 310099 90404 310165 90405
rect 310099 90340 310100 90404
rect 310164 90340 310165 90404
rect 310099 90339 310165 90340
rect 309731 78028 309797 78029
rect 309731 77964 309732 78028
rect 309796 77964 309797 78028
rect 309731 77963 309797 77964
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 304211 28252 304277 28253
rect 304211 28188 304212 28252
rect 304276 28188 304277 28252
rect 304211 28187 304277 28188
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 302187 11796 302253 11797
rect 302187 11732 302188 11796
rect 302252 11732 302253 11796
rect 302187 11731 302253 11732
rect 307794 -1306 308414 20898
rect 309734 11661 309794 77963
rect 310102 11797 310162 90339
rect 311514 61174 312134 94000
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 310099 11796 310165 11797
rect 310099 11732 310100 11796
rect 310164 11732 310165 11796
rect 310099 11731 310165 11732
rect 309731 11660 309797 11661
rect 309731 11596 309732 11660
rect 309796 11596 309797 11660
rect 309731 11595 309797 11596
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 64894 315854 94000
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 68614 319574 94000
rect 321510 77213 321570 97955
rect 324270 93533 324330 99315
rect 324267 93532 324333 93533
rect 324267 93468 324268 93532
rect 324332 93468 324333 93532
rect 324267 93467 324333 93468
rect 321507 77212 321573 77213
rect 321507 77148 321508 77212
rect 321572 77148 321573 77212
rect 321507 77147 321573 77148
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 75454 326414 110898
rect 326662 107133 326722 299507
rect 329514 295174 330134 330618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 335859 371380 335925 371381
rect 335859 371316 335860 371380
rect 335924 371316 335925 371380
rect 335859 371315 335925 371316
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 330339 300932 330405 300933
rect 330339 300868 330340 300932
rect 330404 300868 330405 300932
rect 330339 300867 330405 300868
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 327027 277812 327093 277813
rect 327027 277748 327028 277812
rect 327092 277748 327093 277812
rect 327027 277747 327093 277748
rect 327030 126309 327090 277747
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 328499 220148 328565 220149
rect 328499 220084 328500 220148
rect 328564 220084 328565 220148
rect 328499 220083 328565 220084
rect 327027 126308 327093 126309
rect 327027 126244 327028 126308
rect 327092 126244 327093 126308
rect 327027 126243 327093 126244
rect 326659 107132 326725 107133
rect 326659 107068 326660 107132
rect 326724 107068 326725 107132
rect 326659 107067 326725 107068
rect 328502 106317 328562 220083
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 330342 134197 330402 300867
rect 333234 298894 333854 334338
rect 334019 319428 334085 319429
rect 334019 319364 334020 319428
rect 334084 319364 334085 319428
rect 334019 319363 334085 319364
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 331443 177444 331509 177445
rect 331443 177380 331444 177444
rect 331508 177380 331509 177444
rect 331443 177379 331509 177380
rect 330339 134196 330405 134197
rect 330339 134132 330340 134196
rect 330404 134132 330405 134196
rect 330339 134131 330405 134132
rect 331446 116517 331506 177379
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 331443 116516 331509 116517
rect 331443 116452 331444 116516
rect 331508 116452 331509 116516
rect 331443 116451 331509 116452
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 328499 106316 328565 106317
rect 328499 106252 328500 106316
rect 328564 106252 328565 106316
rect 328499 106251 328565 106252
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 334022 46205 334082 319363
rect 334203 236604 334269 236605
rect 334203 236540 334204 236604
rect 334268 236540 334269 236604
rect 334203 236539 334269 236540
rect 334206 110669 334266 236539
rect 335862 174589 335922 371315
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 342299 318068 342365 318069
rect 342299 318004 342300 318068
rect 342364 318004 342365 318068
rect 342299 318003 342365 318004
rect 340827 316708 340893 316709
rect 340827 316644 340828 316708
rect 340892 316644 340893 316708
rect 340827 316643 340893 316644
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 338619 225724 338685 225725
rect 338619 225660 338620 225724
rect 338684 225660 338685 225724
rect 338619 225659 338685 225660
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 335859 174588 335925 174589
rect 335859 174524 335860 174588
rect 335924 174524 335925 174588
rect 335859 174523 335925 174524
rect 336043 172548 336109 172549
rect 336043 172484 336044 172548
rect 336108 172484 336109 172548
rect 336043 172483 336109 172484
rect 335859 168468 335925 168469
rect 335859 168404 335860 168468
rect 335924 168404 335925 168468
rect 335859 168403 335925 168404
rect 334203 110668 334269 110669
rect 334203 110604 334204 110668
rect 334268 110604 334269 110668
rect 334203 110603 334269 110604
rect 335862 82789 335922 168403
rect 336046 86189 336106 172483
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 338622 115973 338682 225659
rect 339539 184244 339605 184245
rect 339539 184180 339540 184244
rect 339604 184180 339605 184244
rect 339539 184179 339605 184180
rect 338803 165748 338869 165749
rect 338803 165684 338804 165748
rect 338868 165684 338869 165748
rect 338803 165683 338869 165684
rect 338619 115972 338685 115973
rect 338619 115908 338620 115972
rect 338684 115908 338685 115972
rect 338619 115907 338685 115908
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336043 86188 336109 86189
rect 336043 86124 336044 86188
rect 336108 86124 336109 86188
rect 336043 86123 336109 86124
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 335859 82788 335925 82789
rect 335859 82724 335860 82788
rect 335924 82724 335925 82788
rect 335859 82723 335925 82724
rect 336954 50614 337574 86058
rect 338806 81429 338866 165683
rect 339542 109173 339602 184179
rect 339539 109172 339605 109173
rect 339539 109108 339540 109172
rect 339604 109108 339605 109172
rect 339539 109107 339605 109108
rect 338803 81428 338869 81429
rect 338803 81364 338804 81428
rect 338868 81364 338869 81428
rect 338803 81363 338869 81364
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 334019 46204 334085 46205
rect 334019 46140 334020 46204
rect 334084 46140 334085 46204
rect 334019 46139 334085 46140
rect 334022 11797 334082 46139
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 334019 11796 334085 11797
rect 334019 11732 334020 11796
rect 334084 11732 334085 11796
rect 334019 11731 334085 11732
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 340830 3501 340890 316643
rect 342302 87685 342362 318003
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 345611 162892 345677 162893
rect 345611 162828 345612 162892
rect 345676 162828 345677 162892
rect 345611 162827 345677 162828
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 342299 87684 342365 87685
rect 342299 87620 342300 87684
rect 342364 87620 342365 87684
rect 342299 87619 342365 87620
rect 342302 11797 342362 87619
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 345614 41309 345674 162827
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 345611 41308 345677 41309
rect 345611 41244 345612 41308
rect 345676 41244 345677 41308
rect 345611 41243 345677 41244
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 342299 11796 342365 11797
rect 342299 11732 342300 11796
rect 342364 11732 342365 11796
rect 342299 11731 342365 11732
rect 340827 3500 340893 3501
rect 340827 3436 340828 3500
rect 340892 3436 340893 3500
rect 340827 3435 340893 3436
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 181600 420134 204618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 181600 423854 208338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 181600 427574 212058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 181600 434414 182898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 181600 438134 186618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 181600 441854 190338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 181600 445574 194058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 181600 452414 200898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 181600 456134 204618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 181600 459854 208338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 181600 463574 212058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 181600 470414 182898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 181600 474134 186618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 181600 477854 190338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 181600 481574 194058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 181600 488414 200898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 181600 492134 204618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 494099 197980 494165 197981
rect 494099 197916 494100 197980
rect 494164 197916 494165 197980
rect 494099 197915 494165 197916
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 439568 165454 439888 165486
rect 439568 165218 439610 165454
rect 439846 165218 439888 165454
rect 439568 165134 439888 165218
rect 439568 164898 439610 165134
rect 439846 164898 439888 165134
rect 439568 164866 439888 164898
rect 470288 165454 470608 165486
rect 470288 165218 470330 165454
rect 470566 165218 470608 165454
rect 470288 165134 470608 165218
rect 470288 164898 470330 165134
rect 470566 164898 470608 165134
rect 470288 164866 470608 164898
rect 424208 147454 424528 147486
rect 424208 147218 424250 147454
rect 424486 147218 424528 147454
rect 424208 147134 424528 147218
rect 424208 146898 424250 147134
rect 424486 146898 424528 147134
rect 424208 146866 424528 146898
rect 454928 147454 455248 147486
rect 454928 147218 454970 147454
rect 455206 147218 455248 147454
rect 454928 147134 455248 147218
rect 454928 146898 454970 147134
rect 455206 146898 455248 147134
rect 454928 146866 455248 146898
rect 485648 147454 485968 147486
rect 485648 147218 485690 147454
rect 485926 147218 485968 147454
rect 485648 147134 485968 147218
rect 485648 146898 485690 147134
rect 485926 146898 485968 147134
rect 485648 146866 485968 146898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 439568 129454 439888 129486
rect 439568 129218 439610 129454
rect 439846 129218 439888 129454
rect 439568 129134 439888 129218
rect 439568 128898 439610 129134
rect 439846 128898 439888 129134
rect 439568 128866 439888 128898
rect 470288 129454 470608 129486
rect 470288 129218 470330 129454
rect 470566 129218 470608 129454
rect 470288 129134 470608 129218
rect 470288 128898 470330 129134
rect 470566 128898 470608 129134
rect 470288 128866 470608 128898
rect 494102 127941 494162 197915
rect 495234 181600 495854 208338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 496859 173364 496925 173365
rect 496859 173300 496860 173364
rect 496924 173300 496925 173364
rect 496859 173299 496925 173300
rect 494099 127940 494165 127941
rect 494099 127876 494100 127940
rect 494164 127876 494165 127940
rect 494099 127875 494165 127876
rect 424208 111454 424528 111486
rect 424208 111218 424250 111454
rect 424486 111218 424528 111454
rect 424208 111134 424528 111218
rect 424208 110898 424250 111134
rect 424486 110898 424528 111134
rect 424208 110866 424528 110898
rect 454928 111454 455248 111486
rect 454928 111218 454970 111454
rect 455206 111218 455248 111454
rect 454928 111134 455248 111218
rect 454928 110898 454970 111134
rect 455206 110898 455248 111134
rect 454928 110866 455248 110898
rect 485648 111454 485968 111486
rect 485648 111218 485690 111454
rect 485926 111218 485968 111454
rect 485648 111134 485968 111218
rect 485648 110898 485690 111134
rect 485926 110898 485968 111134
rect 485648 110866 485968 110898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 97174 420134 98000
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 64894 423854 98000
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 68614 427574 98000
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 75454 434414 98000
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 79174 438134 98000
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 82894 441854 98000
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 86614 445574 98000
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 93454 452414 98000
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 97174 456134 98000
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 64894 459854 98000
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 68614 463574 98000
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 75454 470414 98000
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 79174 474134 98000
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 82894 477854 98000
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 86614 481574 98000
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 93454 488414 98000
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 97174 492134 98000
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 64894 495854 98000
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 496862 8941 496922 173299
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 496859 8940 496925 8941
rect 496859 8876 496860 8940
rect 496924 8876 496925 8940
rect 496859 8875 496925 8876
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 76618 579218 76854 579454
rect 76618 578898 76854 579134
rect 87882 579218 88118 579454
rect 87882 578898 88118 579134
rect 99146 579218 99382 579454
rect 99146 578898 99382 579134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 82250 561218 82486 561454
rect 82250 560898 82486 561134
rect 93514 561218 93750 561454
rect 93514 560898 93750 561134
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 76618 543218 76854 543454
rect 76618 542898 76854 543134
rect 87882 543218 88118 543454
rect 87882 542898 88118 543134
rect 99146 543218 99382 543454
rect 99146 542898 99382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 75618 471218 75854 471454
rect 75618 470898 75854 471134
rect 84882 471218 85118 471454
rect 84882 470898 85118 471134
rect 94146 471218 94382 471454
rect 94146 470898 94382 471134
rect 80250 453218 80486 453454
rect 80250 452898 80486 453134
rect 89514 453218 89750 453454
rect 89514 452898 89750 453134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 89610 381218 89846 381454
rect 89610 380898 89846 381134
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 74250 363218 74486 363454
rect 74250 362898 74486 363134
rect 104970 363218 105206 363454
rect 104970 362898 105206 363134
rect 89610 345218 89846 345454
rect 89610 344898 89846 345134
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 89610 273218 89846 273454
rect 89610 272898 89846 273134
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 227916 165218 228152 165454
rect 227916 164898 228152 165134
rect 237847 165218 238083 165454
rect 237847 164898 238083 165134
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 227916 129218 228152 129454
rect 227916 128898 228152 129134
rect 237847 129218 238083 129454
rect 237847 128898 238083 129134
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 242813 110898 243049 111134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 314250 165218 314486 165454
rect 314250 164898 314486 165134
rect 317514 165218 317750 165454
rect 317514 164898 317750 165134
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 314250 129218 314486 129454
rect 314250 128898 314486 129134
rect 317514 129218 317750 129454
rect 317514 128898 317750 129134
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 439610 165218 439846 165454
rect 439610 164898 439846 165134
rect 470330 165218 470566 165454
rect 470330 164898 470566 165134
rect 424250 147218 424486 147454
rect 424250 146898 424486 147134
rect 454970 147218 455206 147454
rect 454970 146898 455206 147134
rect 485690 147218 485926 147454
rect 485690 146898 485926 147134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 439610 129218 439846 129454
rect 439610 128898 439846 129134
rect 470330 129218 470566 129454
rect 470330 128898 470566 129134
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 424250 111218 424486 111454
rect 424250 110898 424486 111134
rect 454970 111218 455206 111454
rect 454970 110898 455206 111134
rect 485690 111218 485926 111454
rect 485690 110898 485926 111134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 76618 579454
rect 76854 579218 87882 579454
rect 88118 579218 99146 579454
rect 99382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 76618 579134
rect 76854 578898 87882 579134
rect 88118 578898 99146 579134
rect 99382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 82250 561454
rect 82486 561218 93514 561454
rect 93750 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 82250 561134
rect 82486 560898 93514 561134
rect 93750 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 76618 543454
rect 76854 543218 87882 543454
rect 88118 543218 99146 543454
rect 99382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 76618 543134
rect 76854 542898 87882 543134
rect 88118 542898 99146 543134
rect 99382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 75618 471454
rect 75854 471218 84882 471454
rect 85118 471218 94146 471454
rect 94382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 75618 471134
rect 75854 470898 84882 471134
rect 85118 470898 94146 471134
rect 94382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 80250 453454
rect 80486 453218 89514 453454
rect 89750 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 80250 453134
rect 80486 452898 89514 453134
rect 89750 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 89610 381454
rect 89846 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 89610 381134
rect 89846 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 74250 363454
rect 74486 363218 104970 363454
rect 105206 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 74250 363134
rect 74486 362898 104970 363134
rect 105206 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 89610 345454
rect 89846 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 89610 345134
rect 89846 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 89610 273454
rect 89846 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 89610 273134
rect 89846 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 227916 165454
rect 228152 165218 237847 165454
rect 238083 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 314250 165454
rect 314486 165218 317514 165454
rect 317750 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 439610 165454
rect 439846 165218 470330 165454
rect 470566 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 227916 165134
rect 228152 164898 237847 165134
rect 238083 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 314250 165134
rect 314486 164898 317514 165134
rect 317750 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 439610 165134
rect 439846 164898 470330 165134
rect 470566 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 424250 147454
rect 424486 147218 454970 147454
rect 455206 147218 485690 147454
rect 485926 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 424250 147134
rect 424486 146898 454970 147134
rect 455206 146898 485690 147134
rect 485926 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 227916 129454
rect 228152 129218 237847 129454
rect 238083 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 314250 129454
rect 314486 129218 317514 129454
rect 317750 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 439610 129454
rect 439846 129218 470330 129454
rect 470566 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 227916 129134
rect 228152 128898 237847 129134
rect 238083 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 314250 129134
rect 314486 128898 317514 129134
rect 317750 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 439610 129134
rect 439846 128898 470330 129134
rect 470566 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 424250 111454
rect 424486 111218 454970 111454
rect 455206 111218 485690 111454
rect 485926 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 424250 111134
rect 424486 110898 454970 111134
rect 455206 110898 485690 111134
rect 485926 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_frequency_counter  wrapped_frequency_counter_2
timestamp 0
transform 1 0 70000 0 1 440000
box -10 -52 30000 50000
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
use wrapped_hack_soc_dffram  wrapped_hack_soc_dffram_11
timestamp 0
transform 1 0 420000 0 1 100000
box 0 0 74470 79600
use wrapped_rgb_mixer  wrapped_rgb_mixer_3
timestamp 0
transform 1 0 70000 0 1 540000
box -10 -52 36000 42000
use wrapped_vga_clock  wrapped_vga_clock_1
timestamp 0
transform 1 0 70000 0 1 340000
box -10 -52 46000 46000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 294000 74414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 294000 110414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 388000 74414 438000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 492000 74414 538000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 584000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 388000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 181600 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 181600 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 294000 78134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 294000 114134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 388000 78134 438000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 492000 78134 538000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 584000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 388000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 181600 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 181600 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 294000 81854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 294000 117854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 388000 81854 438000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 492000 81854 538000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 584000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 388000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 181600 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 181600 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 294000 85574 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 388000 85574 438000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 492000 85574 538000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 584000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 294000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 181600 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 181600 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 294000 99854 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 388000 99854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 492000 99854 538000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 584000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 178000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 178000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 181600 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 181600 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 181600 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 294000 103574 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 388000 103574 538000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 584000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 178000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 178000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 181600 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 181600 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 294000 92414 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 388000 92414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 492000 92414 538000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 584000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 178000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 178000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 181600 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 181600 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 294000 96134 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 388000 96134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 492000 96134 538000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 584000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 178000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 178000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 181600 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 181600 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 181600 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
