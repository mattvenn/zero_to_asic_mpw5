VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_vgademo_on_fpga
  CLASS BLOCK ;
  FOREIGN wrapped_vgademo_on_fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 296.000 3.270 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 296.000 14.770 300.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.710 296.000 72.270 300.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.690 296.000 78.250 300.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.210 296.000 83.770 300.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.190 296.000 89.750 300.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 296.000 95.270 300.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.690 296.000 101.250 300.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 296.000 106.770 300.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.190 296.000 112.750 300.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.710 296.000 118.270 300.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.690 296.000 124.250 300.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.730 296.000 20.290 300.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.210 296.000 129.770 300.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.190 296.000 135.750 300.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.710 296.000 141.270 300.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.690 296.000 147.250 300.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.670 296.000 153.230 300.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 296.000 158.750 300.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.170 296.000 164.730 300.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.690 296.000 170.250 300.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.670 296.000 176.230 300.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.190 296.000 181.750 300.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 296.000 26.270 300.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.170 296.000 187.730 300.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 296.000 193.250 300.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 296.000 199.230 300.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.190 296.000 204.750 300.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.170 296.000 210.730 300.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.690 296.000 216.250 300.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.670 296.000 222.230 300.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.650 296.000 228.210 300.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.230 296.000 31.790 300.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.210 296.000 37.770 300.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.730 296.000 43.290 300.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 296.000 49.270 300.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.230 296.000 54.790 300.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.210 296.000 60.770 300.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.730 296.000 66.290 300.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 115.340 300.000 116.540 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 150.700 300.000 151.900 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.100 300.000 155.300 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 158.180 300.000 159.380 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 161.580 300.000 162.780 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.980 300.000 166.180 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 168.380 300.000 169.580 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 172.460 300.000 173.660 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 175.860 300.000 177.060 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.260 300.000 180.460 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.660 300.000 183.860 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 118.740 300.000 119.940 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 186.740 300.000 187.940 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.140 300.000 191.340 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.540 300.000 194.740 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 196.940 300.000 198.140 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.020 300.000 202.220 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 204.420 300.000 205.620 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 207.820 300.000 209.020 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.220 300.000 212.420 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 215.300 300.000 216.500 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 218.700 300.000 219.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.140 300.000 123.340 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 222.100 300.000 223.300 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 225.500 300.000 226.700 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.580 300.000 230.780 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.980 300.000 234.180 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 236.380 300.000 237.580 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.780 300.000 240.980 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 243.860 300.000 245.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.260 300.000 248.460 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.540 300.000 126.740 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.620 300.000 130.820 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.020 300.000 134.220 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.420 300.000 137.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 139.820 300.000 141.020 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 143.900 300.000 145.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 147.300 300.000 148.500 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.660 300.000 251.860 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.340 300.000 269.540 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.900 4.000 281.100 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 272.420 300.000 273.620 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.170 296.000 256.730 300.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.980 4.000 285.180 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.150 296.000 262.710 300.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.890 0.000 64.450 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 275.820 300.000 277.020 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 279.220 300.000 280.420 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.670 0.000 107.230 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 254.060 300.000 255.260 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 282.620 300.000 283.820 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.670 296.000 268.230 300.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 286.700 300.000 287.900 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 0.000 150.010 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.650 296.000 274.210 300.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.060 4.000 289.260 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.170 296.000 279.730 300.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.820 4.000 294.020 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.150 296.000 285.710 300.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 290.100 300.000 291.300 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 296.000 233.730 300.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.670 296.000 291.230 300.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 293.500 300.000 294.700 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.230 0.000 192.790 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.010 0.000 235.570 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.650 296.000 297.210 300.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 296.900 300.000 298.100 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.900 4.000 298.100 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.790 0.000 278.350 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.140 300.000 259.340 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 296.000 239.710 300.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 296.000 245.230 300.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.540 300.000 262.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.110 0.000 21.670 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 296.000 251.210 300.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 264.940 300.000 266.140 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.780 4.000 2.980 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.620 4.000 45.820 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.380 4.000 50.580 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.460 4.000 54.660 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.220 4.000 59.420 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.300 4.000 63.500 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.380 4.000 67.580 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.140 4.000 72.340 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.220 4.000 76.420 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.980 4.000 81.180 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.060 4.000 85.260 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.860 4.000 7.060 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.140 4.000 89.340 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.900 4.000 94.100 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.980 4.000 98.180 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.740 4.000 102.940 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.820 4.000 107.020 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.900 4.000 111.100 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.660 4.000 115.860 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.740 4.000 119.940 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.820 4.000 124.020 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.580 4.000 128.780 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.940 4.000 11.140 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.660 4.000 132.860 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.420 4.000 137.620 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.700 4.000 15.900 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.780 4.000 19.980 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.860 4.000 24.060 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.620 4.000 28.820 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.700 4.000 32.900 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.460 4.000 37.660 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.500 4.000 141.700 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.020 4.000 185.220 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.100 4.000 189.300 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.860 4.000 194.060 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.940 4.000 198.140 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.700 4.000 202.900 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.780 4.000 206.980 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.860 4.000 211.060 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.620 4.000 215.820 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.700 4.000 219.900 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.780 4.000 223.980 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.580 4.000 145.780 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.540 4.000 228.740 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.620 4.000 232.820 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.380 4.000 237.580 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.460 4.000 241.660 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.540 4.000 245.740 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.300 4.000 250.500 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.380 4.000 254.580 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.140 4.000 259.340 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.220 4.000 263.420 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.300 4.000 267.500 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.340 4.000 150.540 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.060 4.000 272.260 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.140 4.000 276.340 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.420 4.000 154.620 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.180 4.000 159.380 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.260 4.000 163.460 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.340 4.000 167.540 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.100 4.000 172.300 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.180 4.000 176.380 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.940 4.000 181.140 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 1.100 300.000 2.300 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.460 300.000 37.660 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.860 300.000 41.060 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 43.940 300.000 45.140 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.340 300.000 48.540 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 50.740 300.000 51.940 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.140 300.000 55.340 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 58.220 300.000 59.420 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 61.620 300.000 62.820 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.020 300.000 66.220 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.420 300.000 69.620 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 4.500 300.000 5.700 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 72.500 300.000 73.700 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 75.900 300.000 77.100 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 79.300 300.000 80.500 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 82.700 300.000 83.900 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 86.780 300.000 87.980 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 90.180 300.000 91.380 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 93.580 300.000 94.780 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 96.980 300.000 98.180 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.060 300.000 102.260 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 104.460 300.000 105.660 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 7.900 300.000 9.100 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.860 300.000 109.060 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.260 300.000 112.460 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 11.300 300.000 12.500 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 15.380 300.000 16.580 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 18.780 300.000 19.980 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 22.180 300.000 23.380 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 25.580 300.000 26.780 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 29.660 300.000 30.860 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 33.060 300.000 34.260 ;
    END
  END la1_oenb[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 2.480 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 2.480 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 2.480 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 2.480 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 296.000 8.790 300.000 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 2.635 294.400 288.405 ;
      LAYER met1 ;
        RECT 2.830 2.080 297.090 289.300 ;
      LAYER met2 ;
        RECT 3.550 295.720 7.950 297.685 ;
        RECT 9.070 295.720 13.930 297.685 ;
        RECT 15.050 295.720 19.450 297.685 ;
        RECT 20.570 295.720 25.430 297.685 ;
        RECT 26.550 295.720 30.950 297.685 ;
        RECT 32.070 295.720 36.930 297.685 ;
        RECT 38.050 295.720 42.450 297.685 ;
        RECT 43.570 295.720 48.430 297.685 ;
        RECT 49.550 295.720 53.950 297.685 ;
        RECT 55.070 295.720 59.930 297.685 ;
        RECT 61.050 295.720 65.450 297.685 ;
        RECT 66.570 295.720 71.430 297.685 ;
        RECT 72.550 295.720 77.410 297.685 ;
        RECT 78.530 295.720 82.930 297.685 ;
        RECT 84.050 295.720 88.910 297.685 ;
        RECT 90.030 295.720 94.430 297.685 ;
        RECT 95.550 295.720 100.410 297.685 ;
        RECT 101.530 295.720 105.930 297.685 ;
        RECT 107.050 295.720 111.910 297.685 ;
        RECT 113.030 295.720 117.430 297.685 ;
        RECT 118.550 295.720 123.410 297.685 ;
        RECT 124.530 295.720 128.930 297.685 ;
        RECT 130.050 295.720 134.910 297.685 ;
        RECT 136.030 295.720 140.430 297.685 ;
        RECT 141.550 295.720 146.410 297.685 ;
        RECT 147.530 295.720 152.390 297.685 ;
        RECT 153.510 295.720 157.910 297.685 ;
        RECT 159.030 295.720 163.890 297.685 ;
        RECT 165.010 295.720 169.410 297.685 ;
        RECT 170.530 295.720 175.390 297.685 ;
        RECT 176.510 295.720 180.910 297.685 ;
        RECT 182.030 295.720 186.890 297.685 ;
        RECT 188.010 295.720 192.410 297.685 ;
        RECT 193.530 295.720 198.390 297.685 ;
        RECT 199.510 295.720 203.910 297.685 ;
        RECT 205.030 295.720 209.890 297.685 ;
        RECT 211.010 295.720 215.410 297.685 ;
        RECT 216.530 295.720 221.390 297.685 ;
        RECT 222.510 295.720 227.370 297.685 ;
        RECT 228.490 295.720 232.890 297.685 ;
        RECT 234.010 295.720 238.870 297.685 ;
        RECT 239.990 295.720 244.390 297.685 ;
        RECT 245.510 295.720 250.370 297.685 ;
        RECT 251.490 295.720 255.890 297.685 ;
        RECT 257.010 295.720 261.870 297.685 ;
        RECT 262.990 295.720 267.390 297.685 ;
        RECT 268.510 295.720 273.370 297.685 ;
        RECT 274.490 295.720 278.890 297.685 ;
        RECT 280.010 295.720 284.870 297.685 ;
        RECT 285.990 295.720 290.390 297.685 ;
        RECT 291.510 295.720 296.370 297.685 ;
        RECT 2.860 4.280 297.060 295.720 ;
        RECT 2.860 2.050 20.830 4.280 ;
        RECT 21.950 2.050 63.610 4.280 ;
        RECT 64.730 2.050 106.390 4.280 ;
        RECT 107.510 2.050 149.170 4.280 ;
        RECT 150.290 2.050 191.950 4.280 ;
        RECT 193.070 2.050 234.730 4.280 ;
        RECT 235.850 2.050 277.510 4.280 ;
        RECT 278.630 2.050 297.060 4.280 ;
      LAYER met3 ;
        RECT 4.400 296.500 295.600 297.665 ;
        RECT 4.000 295.100 296.000 296.500 ;
        RECT 4.000 294.420 295.600 295.100 ;
        RECT 4.400 293.100 295.600 294.420 ;
        RECT 4.400 292.420 296.000 293.100 ;
        RECT 4.000 291.700 296.000 292.420 ;
        RECT 4.000 289.700 295.600 291.700 ;
        RECT 4.000 289.660 296.000 289.700 ;
        RECT 4.400 288.300 296.000 289.660 ;
        RECT 4.400 287.660 295.600 288.300 ;
        RECT 4.000 286.300 295.600 287.660 ;
        RECT 4.000 285.580 296.000 286.300 ;
        RECT 4.400 284.220 296.000 285.580 ;
        RECT 4.400 283.580 295.600 284.220 ;
        RECT 4.000 282.220 295.600 283.580 ;
        RECT 4.000 281.500 296.000 282.220 ;
        RECT 4.400 280.820 296.000 281.500 ;
        RECT 4.400 279.500 295.600 280.820 ;
        RECT 4.000 278.820 295.600 279.500 ;
        RECT 4.000 277.420 296.000 278.820 ;
        RECT 4.000 276.740 295.600 277.420 ;
        RECT 4.400 275.420 295.600 276.740 ;
        RECT 4.400 274.740 296.000 275.420 ;
        RECT 4.000 274.020 296.000 274.740 ;
        RECT 4.000 272.660 295.600 274.020 ;
        RECT 4.400 272.020 295.600 272.660 ;
        RECT 4.400 270.660 296.000 272.020 ;
        RECT 4.000 269.940 296.000 270.660 ;
        RECT 4.000 267.940 295.600 269.940 ;
        RECT 4.000 267.900 296.000 267.940 ;
        RECT 4.400 266.540 296.000 267.900 ;
        RECT 4.400 265.900 295.600 266.540 ;
        RECT 4.000 264.540 295.600 265.900 ;
        RECT 4.000 263.820 296.000 264.540 ;
        RECT 4.400 263.140 296.000 263.820 ;
        RECT 4.400 261.820 295.600 263.140 ;
        RECT 4.000 261.140 295.600 261.820 ;
        RECT 4.000 259.740 296.000 261.140 ;
        RECT 4.400 257.740 295.600 259.740 ;
        RECT 4.000 255.660 296.000 257.740 ;
        RECT 4.000 254.980 295.600 255.660 ;
        RECT 4.400 253.660 295.600 254.980 ;
        RECT 4.400 252.980 296.000 253.660 ;
        RECT 4.000 252.260 296.000 252.980 ;
        RECT 4.000 250.900 295.600 252.260 ;
        RECT 4.400 250.260 295.600 250.900 ;
        RECT 4.400 248.900 296.000 250.260 ;
        RECT 4.000 248.860 296.000 248.900 ;
        RECT 4.000 246.860 295.600 248.860 ;
        RECT 4.000 246.140 296.000 246.860 ;
        RECT 4.400 245.460 296.000 246.140 ;
        RECT 4.400 244.140 295.600 245.460 ;
        RECT 4.000 243.460 295.600 244.140 ;
        RECT 4.000 242.060 296.000 243.460 ;
        RECT 4.400 241.380 296.000 242.060 ;
        RECT 4.400 240.060 295.600 241.380 ;
        RECT 4.000 239.380 295.600 240.060 ;
        RECT 4.000 237.980 296.000 239.380 ;
        RECT 4.400 235.980 295.600 237.980 ;
        RECT 4.000 234.580 296.000 235.980 ;
        RECT 4.000 233.220 295.600 234.580 ;
        RECT 4.400 232.580 295.600 233.220 ;
        RECT 4.400 231.220 296.000 232.580 ;
        RECT 4.000 231.180 296.000 231.220 ;
        RECT 4.000 229.180 295.600 231.180 ;
        RECT 4.000 229.140 296.000 229.180 ;
        RECT 4.400 227.140 296.000 229.140 ;
        RECT 4.000 227.100 296.000 227.140 ;
        RECT 4.000 225.100 295.600 227.100 ;
        RECT 4.000 224.380 296.000 225.100 ;
        RECT 4.400 223.700 296.000 224.380 ;
        RECT 4.400 222.380 295.600 223.700 ;
        RECT 4.000 221.700 295.600 222.380 ;
        RECT 4.000 220.300 296.000 221.700 ;
        RECT 4.400 218.300 295.600 220.300 ;
        RECT 4.000 216.900 296.000 218.300 ;
        RECT 4.000 216.220 295.600 216.900 ;
        RECT 4.400 214.900 295.600 216.220 ;
        RECT 4.400 214.220 296.000 214.900 ;
        RECT 4.000 212.820 296.000 214.220 ;
        RECT 4.000 211.460 295.600 212.820 ;
        RECT 4.400 210.820 295.600 211.460 ;
        RECT 4.400 209.460 296.000 210.820 ;
        RECT 4.000 209.420 296.000 209.460 ;
        RECT 4.000 207.420 295.600 209.420 ;
        RECT 4.000 207.380 296.000 207.420 ;
        RECT 4.400 206.020 296.000 207.380 ;
        RECT 4.400 205.380 295.600 206.020 ;
        RECT 4.000 204.020 295.600 205.380 ;
        RECT 4.000 203.300 296.000 204.020 ;
        RECT 4.400 202.620 296.000 203.300 ;
        RECT 4.400 201.300 295.600 202.620 ;
        RECT 4.000 200.620 295.600 201.300 ;
        RECT 4.000 198.540 296.000 200.620 ;
        RECT 4.400 196.540 295.600 198.540 ;
        RECT 4.000 195.140 296.000 196.540 ;
        RECT 4.000 194.460 295.600 195.140 ;
        RECT 4.400 193.140 295.600 194.460 ;
        RECT 4.400 192.460 296.000 193.140 ;
        RECT 4.000 191.740 296.000 192.460 ;
        RECT 4.000 189.740 295.600 191.740 ;
        RECT 4.000 189.700 296.000 189.740 ;
        RECT 4.400 188.340 296.000 189.700 ;
        RECT 4.400 187.700 295.600 188.340 ;
        RECT 4.000 186.340 295.600 187.700 ;
        RECT 4.000 185.620 296.000 186.340 ;
        RECT 4.400 184.260 296.000 185.620 ;
        RECT 4.400 183.620 295.600 184.260 ;
        RECT 4.000 182.260 295.600 183.620 ;
        RECT 4.000 181.540 296.000 182.260 ;
        RECT 4.400 180.860 296.000 181.540 ;
        RECT 4.400 179.540 295.600 180.860 ;
        RECT 4.000 178.860 295.600 179.540 ;
        RECT 4.000 177.460 296.000 178.860 ;
        RECT 4.000 176.780 295.600 177.460 ;
        RECT 4.400 175.460 295.600 176.780 ;
        RECT 4.400 174.780 296.000 175.460 ;
        RECT 4.000 174.060 296.000 174.780 ;
        RECT 4.000 172.700 295.600 174.060 ;
        RECT 4.400 172.060 295.600 172.700 ;
        RECT 4.400 170.700 296.000 172.060 ;
        RECT 4.000 169.980 296.000 170.700 ;
        RECT 4.000 167.980 295.600 169.980 ;
        RECT 4.000 167.940 296.000 167.980 ;
        RECT 4.400 166.580 296.000 167.940 ;
        RECT 4.400 165.940 295.600 166.580 ;
        RECT 4.000 164.580 295.600 165.940 ;
        RECT 4.000 163.860 296.000 164.580 ;
        RECT 4.400 163.180 296.000 163.860 ;
        RECT 4.400 161.860 295.600 163.180 ;
        RECT 4.000 161.180 295.600 161.860 ;
        RECT 4.000 159.780 296.000 161.180 ;
        RECT 4.400 157.780 295.600 159.780 ;
        RECT 4.000 155.700 296.000 157.780 ;
        RECT 4.000 155.020 295.600 155.700 ;
        RECT 4.400 153.700 295.600 155.020 ;
        RECT 4.400 153.020 296.000 153.700 ;
        RECT 4.000 152.300 296.000 153.020 ;
        RECT 4.000 150.940 295.600 152.300 ;
        RECT 4.400 150.300 295.600 150.940 ;
        RECT 4.400 148.940 296.000 150.300 ;
        RECT 4.000 148.900 296.000 148.940 ;
        RECT 4.000 146.900 295.600 148.900 ;
        RECT 4.000 146.180 296.000 146.900 ;
        RECT 4.400 145.500 296.000 146.180 ;
        RECT 4.400 144.180 295.600 145.500 ;
        RECT 4.000 143.500 295.600 144.180 ;
        RECT 4.000 142.100 296.000 143.500 ;
        RECT 4.400 141.420 296.000 142.100 ;
        RECT 4.400 140.100 295.600 141.420 ;
        RECT 4.000 139.420 295.600 140.100 ;
        RECT 4.000 138.020 296.000 139.420 ;
        RECT 4.400 136.020 295.600 138.020 ;
        RECT 4.000 134.620 296.000 136.020 ;
        RECT 4.000 133.260 295.600 134.620 ;
        RECT 4.400 132.620 295.600 133.260 ;
        RECT 4.400 131.260 296.000 132.620 ;
        RECT 4.000 131.220 296.000 131.260 ;
        RECT 4.000 129.220 295.600 131.220 ;
        RECT 4.000 129.180 296.000 129.220 ;
        RECT 4.400 127.180 296.000 129.180 ;
        RECT 4.000 127.140 296.000 127.180 ;
        RECT 4.000 125.140 295.600 127.140 ;
        RECT 4.000 124.420 296.000 125.140 ;
        RECT 4.400 123.740 296.000 124.420 ;
        RECT 4.400 122.420 295.600 123.740 ;
        RECT 4.000 121.740 295.600 122.420 ;
        RECT 4.000 120.340 296.000 121.740 ;
        RECT 4.400 118.340 295.600 120.340 ;
        RECT 4.000 116.940 296.000 118.340 ;
        RECT 4.000 116.260 295.600 116.940 ;
        RECT 4.400 114.940 295.600 116.260 ;
        RECT 4.400 114.260 296.000 114.940 ;
        RECT 4.000 112.860 296.000 114.260 ;
        RECT 4.000 111.500 295.600 112.860 ;
        RECT 4.400 110.860 295.600 111.500 ;
        RECT 4.400 109.500 296.000 110.860 ;
        RECT 4.000 109.460 296.000 109.500 ;
        RECT 4.000 107.460 295.600 109.460 ;
        RECT 4.000 107.420 296.000 107.460 ;
        RECT 4.400 106.060 296.000 107.420 ;
        RECT 4.400 105.420 295.600 106.060 ;
        RECT 4.000 104.060 295.600 105.420 ;
        RECT 4.000 103.340 296.000 104.060 ;
        RECT 4.400 102.660 296.000 103.340 ;
        RECT 4.400 101.340 295.600 102.660 ;
        RECT 4.000 100.660 295.600 101.340 ;
        RECT 4.000 98.580 296.000 100.660 ;
        RECT 4.400 96.580 295.600 98.580 ;
        RECT 4.000 95.180 296.000 96.580 ;
        RECT 4.000 94.500 295.600 95.180 ;
        RECT 4.400 93.180 295.600 94.500 ;
        RECT 4.400 92.500 296.000 93.180 ;
        RECT 4.000 91.780 296.000 92.500 ;
        RECT 4.000 89.780 295.600 91.780 ;
        RECT 4.000 89.740 296.000 89.780 ;
        RECT 4.400 88.380 296.000 89.740 ;
        RECT 4.400 87.740 295.600 88.380 ;
        RECT 4.000 86.380 295.600 87.740 ;
        RECT 4.000 85.660 296.000 86.380 ;
        RECT 4.400 84.300 296.000 85.660 ;
        RECT 4.400 83.660 295.600 84.300 ;
        RECT 4.000 82.300 295.600 83.660 ;
        RECT 4.000 81.580 296.000 82.300 ;
        RECT 4.400 80.900 296.000 81.580 ;
        RECT 4.400 79.580 295.600 80.900 ;
        RECT 4.000 78.900 295.600 79.580 ;
        RECT 4.000 77.500 296.000 78.900 ;
        RECT 4.000 76.820 295.600 77.500 ;
        RECT 4.400 75.500 295.600 76.820 ;
        RECT 4.400 74.820 296.000 75.500 ;
        RECT 4.000 74.100 296.000 74.820 ;
        RECT 4.000 72.740 295.600 74.100 ;
        RECT 4.400 72.100 295.600 72.740 ;
        RECT 4.400 70.740 296.000 72.100 ;
        RECT 4.000 70.020 296.000 70.740 ;
        RECT 4.000 68.020 295.600 70.020 ;
        RECT 4.000 67.980 296.000 68.020 ;
        RECT 4.400 66.620 296.000 67.980 ;
        RECT 4.400 65.980 295.600 66.620 ;
        RECT 4.000 64.620 295.600 65.980 ;
        RECT 4.000 63.900 296.000 64.620 ;
        RECT 4.400 63.220 296.000 63.900 ;
        RECT 4.400 61.900 295.600 63.220 ;
        RECT 4.000 61.220 295.600 61.900 ;
        RECT 4.000 59.820 296.000 61.220 ;
        RECT 4.400 57.820 295.600 59.820 ;
        RECT 4.000 55.740 296.000 57.820 ;
        RECT 4.000 55.060 295.600 55.740 ;
        RECT 4.400 53.740 295.600 55.060 ;
        RECT 4.400 53.060 296.000 53.740 ;
        RECT 4.000 52.340 296.000 53.060 ;
        RECT 4.000 50.980 295.600 52.340 ;
        RECT 4.400 50.340 295.600 50.980 ;
        RECT 4.400 48.980 296.000 50.340 ;
        RECT 4.000 48.940 296.000 48.980 ;
        RECT 4.000 46.940 295.600 48.940 ;
        RECT 4.000 46.220 296.000 46.940 ;
        RECT 4.400 45.540 296.000 46.220 ;
        RECT 4.400 44.220 295.600 45.540 ;
        RECT 4.000 43.540 295.600 44.220 ;
        RECT 4.000 42.140 296.000 43.540 ;
        RECT 4.400 41.460 296.000 42.140 ;
        RECT 4.400 40.140 295.600 41.460 ;
        RECT 4.000 39.460 295.600 40.140 ;
        RECT 4.000 38.060 296.000 39.460 ;
        RECT 4.400 36.060 295.600 38.060 ;
        RECT 4.000 34.660 296.000 36.060 ;
        RECT 4.000 33.300 295.600 34.660 ;
        RECT 4.400 32.660 295.600 33.300 ;
        RECT 4.400 31.300 296.000 32.660 ;
        RECT 4.000 31.260 296.000 31.300 ;
        RECT 4.000 29.260 295.600 31.260 ;
        RECT 4.000 29.220 296.000 29.260 ;
        RECT 4.400 27.220 296.000 29.220 ;
        RECT 4.000 27.180 296.000 27.220 ;
        RECT 4.000 25.180 295.600 27.180 ;
        RECT 4.000 24.460 296.000 25.180 ;
        RECT 4.400 23.780 296.000 24.460 ;
        RECT 4.400 22.460 295.600 23.780 ;
        RECT 4.000 21.780 295.600 22.460 ;
        RECT 4.000 20.380 296.000 21.780 ;
        RECT 4.400 18.380 295.600 20.380 ;
        RECT 4.000 16.980 296.000 18.380 ;
        RECT 4.000 16.300 295.600 16.980 ;
        RECT 4.400 14.980 295.600 16.300 ;
        RECT 4.400 14.300 296.000 14.980 ;
        RECT 4.000 12.900 296.000 14.300 ;
        RECT 4.000 11.540 295.600 12.900 ;
        RECT 4.400 10.900 295.600 11.540 ;
        RECT 4.400 9.540 296.000 10.900 ;
        RECT 4.000 9.500 296.000 9.540 ;
        RECT 4.000 7.500 295.600 9.500 ;
        RECT 4.000 7.460 296.000 7.500 ;
        RECT 4.400 6.100 296.000 7.460 ;
        RECT 4.400 5.460 295.600 6.100 ;
        RECT 4.000 4.100 295.600 5.460 ;
        RECT 4.000 3.380 296.000 4.100 ;
        RECT 4.400 2.700 296.000 3.380 ;
        RECT 4.400 2.555 295.600 2.700 ;
      LAYER met4 ;
        RECT 19.615 19.895 20.640 283.385 ;
        RECT 23.040 19.895 97.440 283.385 ;
        RECT 99.840 19.895 174.240 283.385 ;
        RECT 176.640 19.895 183.705 283.385 ;
  END
END wrapped_vgademo_on_fpga
END LIBRARY

