magic
tech sky130A
magscale 1 2
timestamp 1647805935
<< metal1 >>
rect 201494 703264 201500 703316
rect 201552 703304 201558 703316
rect 202782 703304 202788 703316
rect 201552 703276 202788 703304
rect 201552 703264 201558 703276
rect 202782 703264 202788 703276
rect 202840 703264 202846 703316
rect 82078 703196 82084 703248
rect 82136 703236 82142 703248
rect 267642 703236 267648 703248
rect 82136 703208 267648 703236
rect 82136 703196 82142 703208
rect 267642 703196 267648 703208
rect 267700 703196 267706 703248
rect 99282 703128 99288 703180
rect 99340 703168 99346 703180
rect 332502 703168 332508 703180
rect 99340 703140 332508 703168
rect 99340 703128 99346 703140
rect 332502 703128 332508 703140
rect 332560 703128 332566 703180
rect 115198 703060 115204 703112
rect 115256 703100 115262 703112
rect 348786 703100 348792 703112
rect 115256 703072 348792 703100
rect 115256 703060 115262 703072
rect 348786 703060 348792 703072
rect 348844 703060 348850 703112
rect 79318 702992 79324 703044
rect 79376 703032 79382 703044
rect 364334 703032 364340 703044
rect 79376 703004 364340 703032
rect 79376 702992 79382 703004
rect 364334 702992 364340 703004
rect 364392 703032 364398 703044
rect 364978 703032 364984 703044
rect 364392 703004 364984 703032
rect 364392 702992 364398 703004
rect 364978 702992 364984 703004
rect 365036 702992 365042 703044
rect 107562 702924 107568 702976
rect 107620 702964 107626 702976
rect 413646 702964 413652 702976
rect 107620 702936 413652 702964
rect 107620 702924 107626 702936
rect 413646 702924 413652 702936
rect 413704 702924 413710 702976
rect 116578 702856 116584 702908
rect 116636 702896 116642 702908
rect 462314 702896 462320 702908
rect 116636 702868 462320 702896
rect 116636 702856 116642 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 78582 702788 78588 702840
rect 78640 702828 78646 702840
rect 429194 702828 429200 702840
rect 78640 702800 429200 702828
rect 78640 702788 78646 702800
rect 429194 702788 429200 702800
rect 429252 702828 429258 702840
rect 429838 702828 429844 702840
rect 429252 702800 429844 702828
rect 429252 702788 429258 702800
rect 429838 702788 429844 702800
rect 429896 702788 429902 702840
rect 71774 702720 71780 702772
rect 71832 702760 71838 702772
rect 72970 702760 72976 702772
rect 71832 702732 72976 702760
rect 71832 702720 71838 702732
rect 72970 702720 72976 702732
rect 73028 702720 73034 702772
rect 113818 702720 113824 702772
rect 113876 702760 113882 702772
rect 478506 702760 478512 702772
rect 113876 702732 478512 702760
rect 113876 702720 113882 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 115290 702652 115296 702704
rect 115348 702692 115354 702704
rect 453942 702692 453948 702704
rect 115348 702664 453948 702692
rect 115348 702652 115354 702664
rect 453942 702652 453948 702664
rect 454000 702652 454006 702704
rect 492582 702652 492588 702704
rect 492640 702692 492646 702704
rect 494790 702692 494796 702704
rect 492640 702664 494796 702692
rect 492640 702652 492646 702664
rect 494790 702652 494796 702664
rect 494848 702652 494854 702704
rect 69198 702584 69204 702636
rect 69256 702624 69262 702636
rect 580902 702624 580908 702636
rect 69256 702596 580908 702624
rect 69256 702584 69262 702596
rect 580902 702584 580908 702596
rect 580960 702584 580966 702636
rect 113082 702516 113088 702568
rect 113140 702556 113146 702568
rect 521562 702556 521568 702568
rect 113140 702528 521568 702556
rect 113140 702516 113146 702528
rect 521562 702516 521568 702528
rect 521620 702516 521626 702568
rect 550542 702516 550548 702568
rect 550600 702556 550606 702568
rect 559650 702556 559656 702568
rect 550600 702528 559656 702556
rect 550600 702516 550606 702528
rect 559650 702516 559656 702528
rect 559708 702516 559714 702568
rect 80698 702448 80704 702500
rect 80756 702488 80762 702500
rect 527174 702488 527180 702500
rect 80756 702460 527180 702488
rect 80756 702448 80762 702460
rect 527174 702448 527180 702460
rect 527232 702448 527238 702500
rect 519538 700952 519544 701004
rect 519596 700992 519602 701004
rect 521562 700992 521568 701004
rect 519596 700964 521568 700992
rect 519596 700952 519602 700964
rect 521562 700952 521568 700964
rect 521620 700952 521626 701004
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 75178 700380 75184 700392
rect 40552 700352 75184 700380
rect 40552 700340 40558 700352
rect 75178 700340 75184 700352
rect 75236 700340 75242 700392
rect 128998 700340 129004 700392
rect 129056 700380 129062 700392
rect 154114 700380 154120 700392
rect 129056 700352 154120 700380
rect 129056 700340 129062 700352
rect 154114 700340 154120 700352
rect 154172 700340 154178 700392
rect 188338 700340 188344 700392
rect 188396 700380 188402 700392
rect 218974 700380 218980 700392
rect 188396 700352 218980 700380
rect 188396 700340 188402 700352
rect 218974 700340 218980 700352
rect 219032 700340 219038 700392
rect 62022 700272 62028 700324
rect 62080 700312 62086 700324
rect 235166 700312 235172 700324
rect 62080 700284 235172 700312
rect 62080 700272 62086 700284
rect 235166 700272 235172 700284
rect 235224 700272 235230 700324
rect 238018 700272 238024 700324
rect 238076 700312 238082 700324
rect 283834 700312 283840 700324
rect 238076 700284 283840 700312
rect 238076 700272 238082 700284
rect 283834 700272 283840 700284
rect 283892 700272 283898 700324
rect 450538 700272 450544 700324
rect 450596 700312 450602 700324
rect 453942 700312 453948 700324
rect 450596 700284 453948 700312
rect 450596 700272 450602 700284
rect 453942 700272 453948 700284
rect 454000 700312 454006 700324
rect 492582 700312 492588 700324
rect 454000 700284 492588 700312
rect 454000 700272 454006 700284
rect 492582 700272 492588 700284
rect 492640 700272 492646 700324
rect 521562 700272 521568 700324
rect 521620 700312 521626 700324
rect 550542 700312 550548 700324
rect 521620 700284 550548 700312
rect 521620 700272 521626 700284
rect 550542 700272 550548 700284
rect 550600 700272 550606 700324
rect 24302 697552 24308 697604
rect 24360 697592 24366 697604
rect 110598 697592 110604 697604
rect 24360 697564 110604 697592
rect 24360 697552 24366 697564
rect 110598 697552 110604 697564
rect 110656 697552 110662 697604
rect 71038 692044 71044 692096
rect 71096 692084 71102 692096
rect 136634 692084 136640 692096
rect 71096 692056 136640 692084
rect 71096 692044 71102 692056
rect 136634 692044 136640 692056
rect 136692 692044 136698 692096
rect 68922 690616 68928 690668
rect 68980 690656 68986 690668
rect 169754 690656 169760 690668
rect 68980 690628 169760 690656
rect 68980 690616 68986 690628
rect 169754 690616 169760 690628
rect 169812 690616 169818 690668
rect 68646 687896 68652 687948
rect 68704 687936 68710 687948
rect 128998 687936 129004 687948
rect 68704 687908 129004 687936
rect 68704 687896 68710 687908
rect 128998 687896 129004 687908
rect 129056 687896 129062 687948
rect 6914 686468 6920 686520
rect 6972 686508 6978 686520
rect 89714 686508 89720 686520
rect 6972 686480 89720 686508
rect 6972 686468 6978 686480
rect 89714 686468 89720 686480
rect 89772 686468 89778 686520
rect 75178 685788 75184 685840
rect 75236 685828 75242 685840
rect 77110 685828 77116 685840
rect 75236 685800 77116 685828
rect 75236 685788 75242 685800
rect 77110 685788 77116 685800
rect 77168 685788 77174 685840
rect 68830 685108 68836 685160
rect 68888 685148 68894 685160
rect 238018 685148 238024 685160
rect 68888 685120 238024 685148
rect 68888 685108 68894 685120
rect 238018 685108 238024 685120
rect 238076 685108 238082 685160
rect 102226 683748 102232 683800
rect 102284 683788 102290 683800
rect 188338 683788 188344 683800
rect 102284 683760 188344 683788
rect 102284 683748 102290 683760
rect 188338 683748 188344 683760
rect 188396 683748 188402 683800
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 75178 683176 75184 683188
rect 3476 683148 75184 683176
rect 3476 683136 3482 683148
rect 75178 683136 75184 683148
rect 75236 683136 75242 683188
rect 196618 683136 196624 683188
rect 196676 683176 196682 683188
rect 580166 683176 580172 683188
rect 196676 683148 580172 683176
rect 196676 683136 196682 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 90634 681952 90640 681964
rect 55186 681924 90640 681952
rect 55186 681760 55214 681924
rect 90634 681912 90640 681924
rect 90692 681912 90698 681964
rect 59262 681844 59268 681896
rect 59320 681884 59326 681896
rect 70026 681884 70032 681896
rect 59320 681856 70032 681884
rect 59320 681844 59326 681856
rect 70026 681844 70032 681856
rect 70084 681844 70090 681896
rect 57790 681776 57796 681828
rect 57848 681816 57854 681828
rect 80698 681816 80704 681828
rect 57848 681788 80704 681816
rect 57848 681776 57854 681788
rect 80698 681776 80704 681788
rect 80756 681776 80762 681828
rect 4798 681708 4804 681760
rect 4856 681748 4862 681760
rect 55122 681748 55128 681760
rect 4856 681720 55128 681748
rect 4856 681708 4862 681720
rect 55122 681708 55128 681720
rect 55180 681720 55214 681760
rect 55180 681708 55186 681720
rect 109310 681708 109316 681760
rect 109368 681748 109374 681760
rect 125686 681748 125692 681760
rect 109368 681720 125692 681748
rect 109368 681708 109374 681720
rect 125686 681708 125692 681720
rect 125744 681708 125750 681760
rect 53742 680960 53748 681012
rect 53800 681000 53806 681012
rect 71774 681000 71780 681012
rect 53800 680972 71780 681000
rect 53800 680960 53806 680972
rect 71774 680960 71780 680972
rect 71832 680960 71838 681012
rect 104894 680960 104900 681012
rect 104952 681000 104958 681012
rect 113174 681000 113180 681012
rect 104952 680972 113180 681000
rect 104952 680960 104958 680972
rect 113174 680960 113180 680972
rect 113232 680960 113238 681012
rect 69106 680348 69112 680400
rect 69164 680388 69170 680400
rect 72602 680388 72608 680400
rect 69164 680360 72608 680388
rect 69164 680348 69170 680360
rect 72602 680348 72608 680360
rect 72660 680348 72666 680400
rect 84838 680348 84844 680400
rect 84896 680388 84902 680400
rect 580258 680388 580264 680400
rect 84896 680360 580264 680388
rect 84896 680348 84902 680360
rect 580258 680348 580264 680360
rect 580316 680348 580322 680400
rect 69290 679328 69296 679380
rect 69348 679368 69354 679380
rect 71038 679368 71044 679380
rect 69348 679340 71044 679368
rect 69348 679328 69354 679340
rect 71038 679328 71044 679340
rect 71096 679328 71102 679380
rect 111794 677628 111800 677680
rect 111852 677668 111858 677680
rect 118694 677668 118700 677680
rect 111852 677640 118700 677668
rect 111852 677628 111858 677640
rect 118694 677628 118700 677640
rect 118752 677628 118758 677680
rect 64690 677560 64696 677612
rect 64748 677600 64754 677612
rect 67634 677600 67640 677612
rect 64748 677572 67640 677600
rect 64748 677560 64754 677572
rect 67634 677560 67640 677572
rect 67692 677560 67698 677612
rect 112346 677560 112352 677612
rect 112404 677600 112410 677612
rect 122926 677600 122932 677612
rect 112404 677572 122932 677600
rect 112404 677560 112410 677572
rect 122926 677560 122932 677572
rect 122984 677560 122990 677612
rect 111794 676268 111800 676320
rect 111852 676308 111858 676320
rect 120350 676308 120356 676320
rect 111852 676280 120356 676308
rect 111852 676268 111858 676280
rect 120350 676268 120356 676280
rect 120408 676268 120414 676320
rect 33042 676200 33048 676252
rect 33100 676240 33106 676252
rect 67634 676240 67640 676252
rect 33100 676212 67640 676240
rect 33100 676200 33106 676212
rect 67634 676200 67640 676212
rect 67692 676200 67698 676252
rect 112714 676200 112720 676252
rect 112772 676240 112778 676252
rect 121546 676240 121552 676252
rect 112772 676212 121552 676240
rect 112772 676200 112778 676212
rect 121546 676200 121552 676212
rect 121604 676200 121610 676252
rect 55030 674908 55036 674960
rect 55088 674948 55094 674960
rect 67634 674948 67640 674960
rect 55088 674920 67640 674948
rect 55088 674908 55094 674920
rect 67634 674908 67640 674920
rect 67692 674908 67698 674960
rect 111978 674840 111984 674892
rect 112036 674880 112042 674892
rect 125778 674880 125784 674892
rect 112036 674852 125784 674880
rect 112036 674840 112042 674852
rect 125778 674840 125784 674852
rect 125836 674840 125842 674892
rect 66070 673684 66076 673736
rect 66128 673724 66134 673736
rect 67726 673724 67732 673736
rect 66128 673696 67732 673724
rect 66128 673684 66134 673696
rect 67726 673684 67732 673696
rect 67784 673684 67790 673736
rect 48130 673480 48136 673532
rect 48188 673520 48194 673532
rect 67634 673520 67640 673532
rect 48188 673492 67640 673520
rect 48188 673480 48194 673492
rect 67634 673480 67640 673492
rect 67692 673480 67698 673532
rect 111794 671984 111800 672036
rect 111852 672024 111858 672036
rect 196618 672024 196624 672036
rect 111852 671996 196624 672024
rect 111852 671984 111858 671996
rect 196618 671984 196624 671996
rect 196676 671984 196682 672036
rect 65886 670760 65892 670812
rect 65944 670800 65950 670812
rect 68646 670800 68652 670812
rect 65944 670772 68652 670800
rect 65944 670760 65950 670772
rect 68646 670760 68652 670772
rect 68704 670760 68710 670812
rect 63218 670692 63224 670744
rect 63276 670732 63282 670744
rect 67634 670732 67640 670744
rect 63276 670704 67640 670732
rect 63276 670692 63282 670704
rect 67634 670692 67640 670704
rect 67692 670692 67698 670744
rect 111794 670692 111800 670744
rect 111852 670732 111858 670744
rect 114554 670732 114560 670744
rect 111852 670704 114560 670732
rect 111852 670692 111858 670704
rect 114554 670692 114560 670704
rect 114612 670692 114618 670744
rect 111794 669468 111800 669520
rect 111852 669508 111858 669520
rect 123018 669508 123024 669520
rect 111852 669480 123024 669508
rect 111852 669468 111858 669480
rect 123018 669468 123024 669480
rect 123076 669468 123082 669520
rect 66162 669400 66168 669452
rect 66220 669440 66226 669452
rect 67818 669440 67824 669452
rect 66220 669412 67824 669440
rect 66220 669400 66226 669412
rect 67818 669400 67824 669412
rect 67876 669400 67882 669452
rect 112714 669400 112720 669452
rect 112772 669440 112778 669452
rect 128446 669440 128452 669452
rect 112772 669412 128452 669440
rect 112772 669400 112778 669412
rect 128446 669400 128452 669412
rect 128504 669400 128510 669452
rect 64506 669332 64512 669384
rect 64564 669372 64570 669384
rect 67634 669372 67640 669384
rect 64564 669344 67640 669372
rect 64564 669332 64570 669344
rect 67634 669332 67640 669344
rect 67692 669332 67698 669384
rect 111794 669332 111800 669384
rect 111852 669372 111858 669384
rect 133966 669372 133972 669384
rect 111852 669344 133972 669372
rect 111852 669332 111858 669344
rect 133966 669332 133972 669344
rect 134024 669332 134030 669384
rect 67358 667904 67364 667956
rect 67416 667944 67422 667956
rect 67726 667944 67732 667956
rect 67416 667916 67732 667944
rect 67416 667904 67422 667916
rect 67726 667904 67732 667916
rect 67784 667904 67790 667956
rect 65978 666612 65984 666664
rect 66036 666652 66042 666664
rect 67818 666652 67824 666664
rect 66036 666624 67824 666652
rect 66036 666612 66042 666624
rect 67818 666612 67824 666624
rect 67876 666612 67882 666664
rect 61930 666544 61936 666596
rect 61988 666584 61994 666596
rect 67634 666584 67640 666596
rect 61988 666556 67640 666584
rect 61988 666544 61994 666556
rect 67634 666544 67640 666556
rect 67692 666544 67698 666596
rect 68554 666544 68560 666596
rect 68612 666584 68618 666596
rect 68830 666584 68836 666596
rect 68612 666556 68836 666584
rect 68612 666544 68618 666556
rect 68830 666544 68836 666556
rect 68888 666544 68894 666596
rect 111794 666544 111800 666596
rect 111852 666584 111858 666596
rect 118786 666584 118792 666596
rect 111852 666556 118792 666584
rect 111852 666544 111858 666556
rect 118786 666544 118792 666556
rect 118844 666544 118850 666596
rect 44082 665252 44088 665304
rect 44140 665292 44146 665304
rect 67726 665292 67732 665304
rect 44140 665264 67732 665292
rect 44140 665252 44146 665264
rect 67726 665252 67732 665264
rect 67784 665252 67790 665304
rect 42702 665184 42708 665236
rect 42760 665224 42766 665236
rect 67634 665224 67640 665236
rect 42760 665196 67640 665224
rect 42760 665184 42766 665196
rect 67634 665184 67640 665196
rect 67692 665184 67698 665236
rect 111794 665184 111800 665236
rect 111852 665224 111858 665236
rect 124398 665224 124404 665236
rect 111852 665196 124404 665224
rect 111852 665184 111858 665196
rect 124398 665184 124404 665196
rect 124456 665184 124462 665236
rect 61838 663824 61844 663876
rect 61896 663864 61902 663876
rect 67634 663864 67640 663876
rect 61896 663836 67640 663864
rect 61896 663824 61902 663836
rect 67634 663824 67640 663836
rect 67692 663824 67698 663876
rect 112346 663824 112352 663876
rect 112404 663864 112410 663876
rect 128538 663864 128544 663876
rect 112404 663836 128544 663864
rect 112404 663824 112410 663836
rect 128538 663824 128544 663836
rect 128596 663824 128602 663876
rect 52362 663756 52368 663808
rect 52420 663796 52426 663808
rect 67726 663796 67732 663808
rect 52420 663768 67732 663796
rect 52420 663756 52426 663768
rect 67726 663756 67732 663768
rect 67784 663756 67790 663808
rect 111794 663756 111800 663808
rect 111852 663796 111858 663808
rect 142154 663796 142160 663808
rect 111852 663768 142160 663796
rect 111852 663756 111858 663768
rect 142154 663756 142160 663768
rect 142212 663756 142218 663808
rect 62022 663008 62028 663060
rect 62080 663048 62086 663060
rect 67634 663048 67640 663060
rect 62080 663020 67640 663048
rect 62080 663008 62086 663020
rect 67634 663008 67640 663020
rect 67692 663008 67698 663060
rect 111794 662396 111800 662448
rect 111852 662436 111858 662448
rect 117406 662436 117412 662448
rect 111852 662408 117412 662436
rect 111852 662396 111858 662408
rect 117406 662396 117412 662408
rect 117464 662396 117470 662448
rect 53650 661648 53656 661700
rect 53708 661688 53714 661700
rect 62022 661688 62028 661700
rect 53708 661660 62028 661688
rect 53708 661648 53714 661660
rect 62022 661648 62028 661660
rect 62080 661648 62086 661700
rect 111150 661512 111156 661564
rect 111208 661552 111214 661564
rect 113818 661552 113824 661564
rect 111208 661524 113824 661552
rect 111208 661512 111214 661524
rect 113818 661512 113824 661524
rect 113876 661512 113882 661564
rect 60642 661036 60648 661088
rect 60700 661076 60706 661088
rect 67634 661076 67640 661088
rect 60700 661048 67640 661076
rect 60700 661036 60706 661048
rect 67634 661036 67640 661048
rect 67692 661036 67698 661088
rect 59078 659744 59084 659796
rect 59136 659784 59142 659796
rect 67634 659784 67640 659796
rect 59136 659756 67640 659784
rect 59136 659744 59142 659756
rect 67634 659744 67640 659756
rect 67692 659744 67698 659796
rect 112530 659744 112536 659796
rect 112588 659784 112594 659796
rect 136726 659784 136732 659796
rect 112588 659756 136732 659784
rect 112588 659744 112594 659756
rect 136726 659744 136732 659756
rect 136784 659744 136790 659796
rect 50798 659676 50804 659728
rect 50856 659716 50862 659728
rect 67726 659716 67732 659728
rect 50856 659688 67732 659716
rect 50856 659676 50862 659688
rect 67726 659676 67732 659688
rect 67784 659676 67790 659728
rect 112346 659676 112352 659728
rect 112404 659716 112410 659728
rect 146294 659716 146300 659728
rect 112404 659688 146300 659716
rect 112404 659676 112410 659688
rect 146294 659676 146300 659688
rect 146352 659676 146358 659728
rect 39942 658928 39948 658980
rect 40000 658968 40006 658980
rect 68554 658968 68560 658980
rect 40000 658940 68560 658968
rect 40000 658928 40006 658940
rect 68554 658928 68560 658940
rect 68612 658928 68618 658980
rect 109034 658384 109040 658436
rect 109092 658424 109098 658436
rect 110598 658424 110604 658436
rect 109092 658396 110604 658424
rect 109092 658384 109098 658396
rect 110598 658384 110604 658396
rect 110656 658384 110662 658436
rect 63402 658248 63408 658300
rect 63460 658288 63466 658300
rect 67634 658288 67640 658300
rect 63460 658260 67640 658288
rect 63460 658248 63466 658260
rect 67634 658248 67640 658260
rect 67692 658248 67698 658300
rect 2774 658180 2780 658232
rect 2832 658220 2838 658232
rect 4798 658220 4804 658232
rect 2832 658192 4804 658220
rect 2832 658180 2838 658192
rect 4798 658180 4804 658192
rect 4856 658180 4862 658232
rect 133782 657500 133788 657552
rect 133840 657540 133846 657552
rect 201494 657540 201500 657552
rect 133840 657512 201500 657540
rect 133840 657500 133846 657512
rect 201494 657500 201500 657512
rect 201552 657500 201558 657552
rect 56502 656956 56508 657008
rect 56560 656996 56566 657008
rect 68186 656996 68192 657008
rect 56560 656968 68192 656996
rect 56560 656956 56566 656968
rect 68186 656956 68192 656968
rect 68244 656956 68250 657008
rect 49602 656888 49608 656940
rect 49660 656928 49666 656940
rect 67726 656928 67732 656940
rect 49660 656900 67732 656928
rect 49660 656888 49666 656900
rect 67726 656888 67732 656900
rect 67784 656888 67790 656940
rect 112530 656888 112536 656940
rect 112588 656928 112594 656940
rect 132494 656928 132500 656940
rect 112588 656900 132500 656928
rect 112588 656888 112594 656900
rect 132494 656888 132500 656900
rect 132552 656928 132558 656940
rect 133782 656928 133788 656940
rect 132552 656900 133788 656928
rect 132552 656888 132558 656900
rect 133782 656888 133788 656900
rect 133840 656888 133846 656940
rect 112530 655596 112536 655648
rect 112588 655636 112594 655648
rect 121638 655636 121644 655648
rect 112588 655608 121644 655636
rect 112588 655596 112594 655608
rect 121638 655596 121644 655608
rect 121696 655596 121702 655648
rect 41230 655528 41236 655580
rect 41288 655568 41294 655580
rect 67634 655568 67640 655580
rect 41288 655540 67640 655568
rect 41288 655528 41294 655540
rect 67634 655528 67640 655540
rect 67692 655528 67698 655580
rect 112346 655528 112352 655580
rect 112404 655568 112410 655580
rect 139394 655568 139400 655580
rect 112404 655540 139400 655568
rect 112404 655528 112410 655540
rect 139394 655528 139400 655540
rect 139452 655528 139458 655580
rect 58618 654780 58624 654832
rect 58676 654820 58682 654832
rect 67634 654820 67640 654832
rect 58676 654792 67640 654820
rect 58676 654780 58682 654792
rect 67634 654780 67640 654792
rect 67692 654780 67698 654832
rect 57882 652808 57888 652860
rect 57940 652848 57946 652860
rect 67910 652848 67916 652860
rect 57940 652820 67916 652848
rect 57940 652808 57946 652820
rect 67910 652808 67916 652820
rect 67968 652808 67974 652860
rect 48038 652740 48044 652792
rect 48096 652780 48102 652792
rect 67726 652780 67732 652792
rect 48096 652752 67732 652780
rect 48096 652740 48102 652752
rect 67726 652740 67732 652752
rect 67784 652740 67790 652792
rect 64782 651380 64788 651432
rect 64840 651420 64846 651432
rect 67634 651420 67640 651432
rect 64840 651392 67640 651420
rect 64840 651380 64846 651392
rect 67634 651380 67640 651392
rect 67692 651380 67698 651432
rect 112530 651380 112536 651432
rect 112588 651420 112594 651432
rect 129826 651420 129832 651432
rect 112588 651392 129832 651420
rect 112588 651380 112594 651392
rect 129826 651380 129832 651392
rect 129884 651380 129890 651432
rect 112070 650088 112076 650140
rect 112128 650128 112134 650140
rect 119338 650128 119344 650140
rect 112128 650100 119344 650128
rect 112128 650088 112134 650100
rect 119338 650088 119344 650100
rect 119396 650088 119402 650140
rect 34422 650020 34428 650072
rect 34480 650060 34486 650072
rect 67634 650060 67640 650072
rect 34480 650032 67640 650060
rect 34480 650020 34486 650032
rect 67634 650020 67640 650032
rect 67692 650020 67698 650072
rect 111978 650020 111984 650072
rect 112036 650060 112042 650072
rect 143626 650060 143632 650072
rect 112036 650032 143632 650060
rect 112036 650020 112042 650032
rect 143626 650020 143632 650032
rect 143684 650020 143690 650072
rect 112990 648660 112996 648712
rect 113048 648700 113054 648712
rect 115934 648700 115940 648712
rect 113048 648672 115940 648700
rect 113048 648660 113054 648672
rect 115934 648660 115940 648672
rect 115992 648660 115998 648712
rect 64598 648592 64604 648644
rect 64656 648632 64662 648644
rect 67634 648632 67640 648644
rect 64656 648604 67640 648632
rect 64656 648592 64662 648604
rect 67634 648592 67640 648604
rect 67692 648592 67698 648644
rect 113082 648592 113088 648644
rect 113140 648632 113146 648644
rect 138014 648632 138020 648644
rect 113140 648604 138020 648632
rect 113140 648592 113146 648604
rect 138014 648592 138020 648604
rect 138072 648592 138078 648644
rect 63126 647300 63132 647352
rect 63184 647340 63190 647352
rect 67726 647340 67732 647352
rect 63184 647312 67732 647340
rect 63184 647300 63190 647312
rect 67726 647300 67732 647312
rect 67784 647300 67790 647352
rect 62022 647232 62028 647284
rect 62080 647272 62086 647284
rect 67634 647272 67640 647284
rect 62080 647244 67640 647272
rect 62080 647232 62086 647244
rect 67634 647232 67640 647244
rect 67692 647232 67698 647284
rect 109402 647232 109408 647284
rect 109460 647272 109466 647284
rect 112162 647272 112168 647284
rect 109460 647244 112168 647272
rect 109460 647232 109466 647244
rect 112162 647232 112168 647244
rect 112220 647232 112226 647284
rect 113082 647232 113088 647284
rect 113140 647272 113146 647284
rect 143534 647272 143540 647284
rect 113140 647244 143540 647272
rect 113140 647232 113146 647244
rect 143534 647232 143540 647244
rect 143592 647232 143598 647284
rect 37090 645872 37096 645924
rect 37148 645912 37154 645924
rect 67634 645912 67640 645924
rect 37148 645884 67640 645912
rect 37148 645872 37154 645884
rect 67634 645872 67640 645884
rect 67692 645872 67698 645924
rect 112990 644512 112996 644564
rect 113048 644552 113054 644564
rect 132862 644552 132868 644564
rect 113048 644524 132868 644552
rect 113048 644512 113054 644524
rect 132862 644512 132868 644524
rect 132920 644512 132926 644564
rect 113082 644444 113088 644496
rect 113140 644484 113146 644496
rect 135254 644484 135260 644496
rect 113140 644456 135260 644484
rect 113140 644444 113146 644456
rect 135254 644444 135260 644456
rect 135312 644444 135318 644496
rect 112806 644308 112812 644360
rect 112864 644348 112870 644360
rect 115290 644348 115296 644360
rect 112864 644320 115296 644348
rect 112864 644308 112870 644320
rect 115290 644308 115296 644320
rect 115348 644308 115354 644360
rect 57790 643696 57796 643748
rect 57848 643736 57854 643748
rect 69658 643736 69664 643748
rect 57848 643708 69664 643736
rect 57848 643696 57854 643708
rect 69658 643696 69664 643708
rect 69716 643696 69722 643748
rect 119338 643696 119344 643748
rect 119396 643736 119402 643748
rect 134058 643736 134064 643748
rect 119396 643708 134064 643736
rect 119396 643696 119402 643708
rect 134058 643696 134064 643708
rect 134116 643736 134122 643748
rect 135162 643736 135168 643748
rect 134116 643708 135168 643736
rect 134116 643696 134122 643708
rect 135162 643696 135168 643708
rect 135220 643696 135226 643748
rect 135162 643084 135168 643136
rect 135220 643124 135226 643136
rect 580166 643124 580172 643136
rect 135220 643096 580172 643124
rect 135220 643084 135226 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 116026 643016 116032 643068
rect 116084 643056 116090 643068
rect 116578 643056 116584 643068
rect 116084 643028 116584 643056
rect 116084 643016 116090 643028
rect 116578 643016 116584 643028
rect 116636 643016 116642 643068
rect 112622 642064 112628 642116
rect 112680 642104 112686 642116
rect 116026 642104 116032 642116
rect 112680 642076 116032 642104
rect 112680 642064 112686 642076
rect 116026 642064 116032 642076
rect 116084 642064 116090 642116
rect 61746 641792 61752 641844
rect 61804 641832 61810 641844
rect 67726 641832 67732 641844
rect 61804 641804 67732 641832
rect 61804 641792 61810 641804
rect 67726 641792 67732 641804
rect 67784 641792 67790 641844
rect 37182 641724 37188 641776
rect 37240 641764 37246 641776
rect 67634 641764 67640 641776
rect 37240 641736 67640 641764
rect 37240 641724 37246 641736
rect 67634 641724 67640 641736
rect 67692 641724 67698 641776
rect 113082 641724 113088 641776
rect 113140 641764 113146 641776
rect 140774 641764 140780 641776
rect 113140 641736 140780 641764
rect 113140 641724 113146 641736
rect 140774 641724 140780 641736
rect 140832 641724 140838 641776
rect 63310 640364 63316 640416
rect 63368 640404 63374 640416
rect 67634 640404 67640 640416
rect 63368 640376 67640 640404
rect 63368 640364 63374 640376
rect 67634 640364 67640 640376
rect 67692 640364 67698 640416
rect 34146 640296 34152 640348
rect 34204 640336 34210 640348
rect 67726 640336 67732 640348
rect 34204 640308 67732 640336
rect 34204 640296 34210 640308
rect 67726 640296 67732 640308
rect 67784 640296 67790 640348
rect 108850 639616 108856 639668
rect 108908 639656 108914 639668
rect 112254 639656 112260 639668
rect 108908 639628 112260 639656
rect 108908 639616 108914 639628
rect 112254 639616 112260 639628
rect 112312 639616 112318 639668
rect 124122 639548 124128 639600
rect 124180 639588 124186 639600
rect 299474 639588 299480 639600
rect 124180 639560 299480 639588
rect 124180 639548 124186 639560
rect 299474 639548 299480 639560
rect 299532 639548 299538 639600
rect 38562 638936 38568 638988
rect 38620 638976 38626 638988
rect 71314 638976 71320 638988
rect 38620 638948 71320 638976
rect 38620 638936 38626 638948
rect 71314 638936 71320 638948
rect 71372 638936 71378 638988
rect 112898 638936 112904 638988
rect 112956 638976 112962 638988
rect 129918 638976 129924 638988
rect 112956 638948 129924 638976
rect 112956 638936 112962 638948
rect 129918 638936 129924 638948
rect 129976 638936 129982 638988
rect 46842 638868 46848 638920
rect 46900 638908 46906 638920
rect 53742 638908 53748 638920
rect 46900 638880 53748 638908
rect 46900 638868 46906 638880
rect 53742 638868 53748 638880
rect 53800 638908 53806 638920
rect 73890 638908 73896 638920
rect 53800 638880 73896 638908
rect 53800 638868 53806 638880
rect 73890 638868 73896 638880
rect 73948 638868 73954 638920
rect 104158 638868 104164 638920
rect 104216 638908 104222 638920
rect 122834 638908 122840 638920
rect 104216 638880 122840 638908
rect 104216 638868 104222 638880
rect 122834 638868 122840 638880
rect 122892 638908 122898 638920
rect 124122 638908 124128 638920
rect 122892 638880 124128 638908
rect 122892 638868 122898 638880
rect 124122 638868 124128 638880
rect 124180 638868 124186 638920
rect 72694 638460 72700 638512
rect 72752 638500 72758 638512
rect 84194 638500 84200 638512
rect 72752 638472 84200 638500
rect 72752 638460 72758 638472
rect 84194 638460 84200 638472
rect 84252 638460 84258 638512
rect 95142 638460 95148 638512
rect 95200 638500 95206 638512
rect 105538 638500 105544 638512
rect 95200 638472 105544 638500
rect 95200 638460 95206 638472
rect 105538 638460 105544 638472
rect 105596 638460 105602 638512
rect 108942 638460 108948 638512
rect 109000 638500 109006 638512
rect 124306 638500 124312 638512
rect 109000 638472 124312 638500
rect 109000 638460 109006 638472
rect 124306 638460 124312 638472
rect 124364 638460 124370 638512
rect 57790 638392 57796 638444
rect 57848 638432 57854 638444
rect 82262 638432 82268 638444
rect 57848 638404 82268 638432
rect 57848 638392 57854 638404
rect 82262 638392 82268 638404
rect 82320 638392 82326 638444
rect 99006 638392 99012 638444
rect 99064 638432 99070 638444
rect 117314 638432 117320 638444
rect 99064 638404 117320 638432
rect 99064 638392 99070 638404
rect 117314 638392 117320 638404
rect 117372 638392 117378 638444
rect 54754 638324 54760 638376
rect 54812 638364 54818 638376
rect 82906 638364 82912 638376
rect 54812 638336 82912 638364
rect 54812 638324 54818 638336
rect 82906 638324 82912 638336
rect 82964 638324 82970 638376
rect 99650 638324 99656 638376
rect 99708 638364 99714 638376
rect 121454 638364 121460 638376
rect 99708 638336 121460 638364
rect 99708 638324 99714 638336
rect 121454 638324 121460 638336
rect 121512 638324 121518 638376
rect 48222 638256 48228 638308
rect 48280 638296 48286 638308
rect 79042 638296 79048 638308
rect 48280 638268 79048 638296
rect 48280 638256 48286 638268
rect 79042 638256 79048 638268
rect 79100 638256 79106 638308
rect 102870 638256 102876 638308
rect 102928 638296 102934 638308
rect 131114 638296 131120 638308
rect 102928 638268 131120 638296
rect 102928 638256 102934 638268
rect 131114 638256 131120 638268
rect 131172 638256 131178 638308
rect 3418 638188 3424 638240
rect 3476 638228 3482 638240
rect 59170 638228 59176 638240
rect 3476 638200 59176 638228
rect 3476 638188 3482 638200
rect 59170 638188 59176 638200
rect 59228 638228 59234 638240
rect 91922 638228 91928 638240
rect 59228 638200 91928 638228
rect 59228 638188 59234 638200
rect 91922 638188 91928 638200
rect 91980 638188 91986 638240
rect 96430 638188 96436 638240
rect 96488 638228 96494 638240
rect 124214 638228 124220 638240
rect 96488 638200 124220 638228
rect 96488 638188 96494 638200
rect 124214 638188 124220 638200
rect 124272 638188 124278 638240
rect 96522 637984 96528 638036
rect 96580 638024 96586 638036
rect 99650 638024 99656 638036
rect 96580 637996 99656 638024
rect 96580 637984 96586 637996
rect 99650 637984 99656 637996
rect 99708 637984 99714 638036
rect 74442 637576 74448 637628
rect 74500 637616 74506 637628
rect 74500 637588 74580 637616
rect 74500 637576 74506 637588
rect 74552 637548 74580 637588
rect 93854 637576 93860 637628
rect 93912 637616 93918 637628
rect 101398 637616 101404 637628
rect 93912 637588 101404 637616
rect 93912 637576 93918 637588
rect 101398 637576 101404 637588
rect 101456 637576 101462 637628
rect 75822 637548 75828 637560
rect 74552 637520 75828 637548
rect 75822 637508 75828 637520
rect 75880 637508 75886 637560
rect 75914 637440 75920 637492
rect 75972 637480 75978 637492
rect 77110 637480 77116 637492
rect 75972 637452 77116 637480
rect 75972 637440 75978 637452
rect 77110 637440 77116 637452
rect 77168 637440 77174 637492
rect 85574 637440 85580 637492
rect 85632 637480 85638 637492
rect 86770 637480 86776 637492
rect 85632 637452 86776 637480
rect 85632 637440 85638 637452
rect 86770 637440 86776 637452
rect 86828 637440 86834 637492
rect 86954 637440 86960 637492
rect 87012 637480 87018 637492
rect 88058 637480 88064 637492
rect 87012 637452 88064 637480
rect 87012 637440 87018 637452
rect 88058 637440 88064 637452
rect 88116 637440 88122 637492
rect 96614 637440 96620 637492
rect 96672 637480 96678 637492
rect 97718 637480 97724 637492
rect 96672 637452 97724 637480
rect 96672 637440 96678 637452
rect 97718 637440 97724 637452
rect 97776 637440 97782 637492
rect 103606 637440 103612 637492
rect 103664 637480 103670 637492
rect 104802 637480 104808 637492
rect 103664 637452 104808 637480
rect 103664 637440 103670 637452
rect 104802 637440 104808 637452
rect 104860 637440 104866 637492
rect 69198 637168 69204 637220
rect 69256 637208 69262 637220
rect 69750 637208 69756 637220
rect 69256 637180 69756 637208
rect 69256 637168 69262 637180
rect 69750 637168 69756 637180
rect 69808 637168 69814 637220
rect 52270 636964 52276 637016
rect 52328 637004 52334 637016
rect 78398 637004 78404 637016
rect 52328 636976 78404 637004
rect 52328 636964 52334 636976
rect 78398 636964 78404 636976
rect 78456 636964 78462 637016
rect 101582 636964 101588 637016
rect 101640 637004 101646 637016
rect 128354 637004 128360 637016
rect 101640 636976 128360 637004
rect 101640 636964 101646 636976
rect 128354 636964 128360 636976
rect 128412 636964 128418 637016
rect 45370 636896 45376 636948
rect 45428 636936 45434 636948
rect 74534 636936 74540 636948
rect 45428 636908 74540 636936
rect 45428 636896 45434 636908
rect 74534 636896 74540 636908
rect 74592 636896 74598 636948
rect 88702 636896 88708 636948
rect 88760 636936 88766 636948
rect 118878 636936 118884 636948
rect 88760 636908 118884 636936
rect 88760 636896 88766 636908
rect 118878 636896 118884 636908
rect 118936 636896 118942 636948
rect 50982 636828 50988 636880
rect 51040 636868 51046 636880
rect 84838 636868 84844 636880
rect 51040 636840 84844 636868
rect 51040 636828 51046 636840
rect 84838 636828 84844 636840
rect 84896 636828 84902 636880
rect 103514 636828 103520 636880
rect 103572 636868 103578 636880
rect 136634 636868 136640 636880
rect 103572 636840 136640 636868
rect 103572 636828 103578 636840
rect 136634 636828 136640 636840
rect 136692 636828 136698 636880
rect 60366 635740 60372 635792
rect 60424 635780 60430 635792
rect 71958 635780 71964 635792
rect 60424 635752 71964 635780
rect 60424 635740 60430 635752
rect 71958 635740 71964 635752
rect 72016 635740 72022 635792
rect 56318 635672 56324 635724
rect 56376 635712 56382 635724
rect 73246 635712 73252 635724
rect 56376 635684 73252 635712
rect 56376 635672 56382 635684
rect 73246 635672 73252 635684
rect 73304 635672 73310 635724
rect 73798 635672 73804 635724
rect 73856 635712 73862 635724
rect 92566 635712 92572 635724
rect 73856 635684 92572 635712
rect 73856 635672 73862 635684
rect 92566 635672 92572 635684
rect 92624 635672 92630 635724
rect 94498 635672 94504 635724
rect 94556 635712 94562 635724
rect 120074 635712 120080 635724
rect 94556 635684 120080 635712
rect 94556 635672 94562 635684
rect 120074 635672 120080 635684
rect 120132 635672 120138 635724
rect 55122 635604 55128 635656
rect 55180 635644 55186 635656
rect 80698 635644 80704 635656
rect 55180 635616 80704 635644
rect 55180 635604 55186 635616
rect 80698 635604 80704 635616
rect 80756 635604 80762 635656
rect 93210 635604 93216 635656
rect 93268 635644 93274 635656
rect 126974 635644 126980 635656
rect 93268 635616 126980 635644
rect 93268 635604 93274 635616
rect 126974 635604 126980 635616
rect 127032 635604 127038 635656
rect 50706 635536 50712 635588
rect 50764 635576 50770 635588
rect 80974 635576 80980 635588
rect 50764 635548 80980 635576
rect 50764 635536 50770 635548
rect 80974 635536 80980 635548
rect 81032 635536 81038 635588
rect 91278 635536 91284 635588
rect 91336 635576 91342 635588
rect 125594 635576 125600 635588
rect 91336 635548 125600 635576
rect 91336 635536 91342 635548
rect 125594 635536 125600 635548
rect 125652 635536 125658 635588
rect 4062 635468 4068 635520
rect 4120 635508 4126 635520
rect 96522 635508 96528 635520
rect 4120 635480 96528 635508
rect 4120 635468 4126 635480
rect 96522 635468 96528 635480
rect 96580 635468 96586 635520
rect 102226 635468 102232 635520
rect 102284 635508 102290 635520
rect 133874 635508 133880 635520
rect 102284 635480 133880 635508
rect 102284 635468 102290 635480
rect 133874 635468 133880 635480
rect 133932 635468 133938 635520
rect 133874 634788 133880 634840
rect 133932 634828 133938 634840
rect 579798 634828 579804 634840
rect 133932 634800 579804 634828
rect 133932 634788 133938 634800
rect 579798 634788 579804 634800
rect 579856 634788 579862 634840
rect 53742 634108 53748 634160
rect 53800 634148 53806 634160
rect 87414 634148 87420 634160
rect 53800 634120 87420 634148
rect 53800 634108 53806 634120
rect 87414 634108 87420 634120
rect 87472 634108 87478 634160
rect 99926 634108 99932 634160
rect 99984 634148 99990 634160
rect 132678 634148 132684 634160
rect 99984 634120 132684 634148
rect 99984 634108 99990 634120
rect 132678 634108 132684 634120
rect 132736 634108 132742 634160
rect 3418 634040 3424 634092
rect 3476 634080 3482 634092
rect 108022 634080 108028 634092
rect 3476 634052 108028 634080
rect 3476 634040 3482 634052
rect 108022 634040 108028 634052
rect 108080 634080 108086 634092
rect 127158 634080 127164 634092
rect 108080 634052 127164 634080
rect 108080 634040 108086 634052
rect 127158 634040 127164 634052
rect 127216 634040 127222 634092
rect 107562 632952 107568 633004
rect 107620 632992 107626 633004
rect 121546 632992 121552 633004
rect 107620 632964 121552 632992
rect 107620 632952 107626 632964
rect 121546 632952 121552 632964
rect 121604 632952 121610 633004
rect 54938 632884 54944 632936
rect 54996 632924 55002 632936
rect 83550 632924 83556 632936
rect 54996 632896 83556 632924
rect 54996 632884 55002 632896
rect 83550 632884 83556 632896
rect 83608 632884 83614 632936
rect 57698 632816 57704 632868
rect 57756 632856 57762 632868
rect 86126 632856 86132 632868
rect 57756 632828 86132 632856
rect 57756 632816 57762 632828
rect 86126 632816 86132 632828
rect 86184 632816 86190 632868
rect 89990 632816 89996 632868
rect 90048 632856 90054 632868
rect 121546 632856 121552 632868
rect 90048 632828 121552 632856
rect 90048 632816 90054 632828
rect 121546 632816 121552 632828
rect 121604 632816 121610 632868
rect 52086 632748 52092 632800
rect 52144 632788 52150 632800
rect 81618 632788 81624 632800
rect 52144 632760 81624 632788
rect 52144 632748 52150 632760
rect 81618 632748 81624 632760
rect 81676 632748 81682 632800
rect 97074 632748 97080 632800
rect 97132 632788 97138 632800
rect 129734 632788 129740 632800
rect 97132 632760 129740 632788
rect 97132 632748 97138 632760
rect 129734 632748 129740 632760
rect 129792 632748 129798 632800
rect 39758 632680 39764 632732
rect 39816 632720 39822 632732
rect 71774 632720 71780 632732
rect 39816 632692 71780 632720
rect 39816 632680 39822 632692
rect 71774 632680 71780 632692
rect 71832 632680 71838 632732
rect 96614 632680 96620 632732
rect 96672 632720 96678 632732
rect 131298 632720 131304 632732
rect 96672 632692 131304 632720
rect 96672 632680 96678 632692
rect 131298 632680 131304 632692
rect 131356 632680 131362 632732
rect 45278 629960 45284 630012
rect 45336 630000 45342 630012
rect 70670 630000 70676 630012
rect 45336 629972 70676 630000
rect 45336 629960 45342 629972
rect 70670 629960 70676 629972
rect 70728 629960 70734 630012
rect 42518 629892 42524 629944
rect 42576 629932 42582 629944
rect 76466 629932 76472 629944
rect 42576 629904 76472 629932
rect 42576 629892 42582 629904
rect 76466 629892 76472 629904
rect 76524 629892 76530 629944
rect 98362 629892 98368 629944
rect 98420 629932 98426 629944
rect 131758 629932 131764 629944
rect 98420 629904 131764 629932
rect 98420 629892 98426 629904
rect 131758 629892 131764 629904
rect 131816 629892 131822 629944
rect 46750 627308 46756 627360
rect 46808 627348 46814 627360
rect 75914 627348 75920 627360
rect 46808 627320 75920 627348
rect 46808 627308 46814 627320
rect 75914 627308 75920 627320
rect 75972 627308 75978 627360
rect 49326 627240 49332 627292
rect 49384 627280 49390 627292
rect 79686 627280 79692 627292
rect 49384 627252 79692 627280
rect 49384 627240 49390 627252
rect 79686 627240 79692 627252
rect 79744 627240 79750 627292
rect 43990 627172 43996 627224
rect 44048 627212 44054 627224
rect 74626 627212 74632 627224
rect 44048 627184 74632 627212
rect 44048 627172 44054 627184
rect 74626 627172 74632 627184
rect 74684 627172 74690 627224
rect 3510 618604 3516 618656
rect 3568 618644 3574 618656
rect 7558 618644 7564 618656
rect 3568 618616 7564 618644
rect 3568 618604 3574 618616
rect 7558 618604 7564 618616
rect 7616 618604 7622 618656
rect 115842 618196 115848 618248
rect 115900 618236 115906 618248
rect 118878 618236 118884 618248
rect 115900 618208 118884 618236
rect 115900 618196 115906 618208
rect 118878 618196 118884 618208
rect 118936 618236 118942 618248
rect 580166 618236 580172 618248
rect 118936 618208 580172 618236
rect 118936 618196 118942 618208
rect 580166 618196 580172 618208
rect 580224 618196 580230 618248
rect 80790 591880 80796 591932
rect 80848 591920 80854 591932
rect 84286 591920 84292 591932
rect 80848 591892 84292 591920
rect 80848 591880 80854 591892
rect 84286 591880 84292 591892
rect 84344 591880 84350 591932
rect 385678 590656 385684 590708
rect 385736 590696 385742 590708
rect 579798 590696 579804 590708
rect 385736 590668 579804 590696
rect 385736 590656 385742 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 7558 589908 7564 589960
rect 7616 589948 7622 589960
rect 96154 589948 96160 589960
rect 7616 589920 96160 589948
rect 7616 589908 7622 589920
rect 96154 589908 96160 589920
rect 96212 589948 96218 589960
rect 96430 589948 96436 589960
rect 96212 589920 96436 589948
rect 96212 589908 96218 589920
rect 96430 589908 96436 589920
rect 96488 589908 96494 589960
rect 96062 588548 96068 588600
rect 96120 588588 96126 588600
rect 121730 588588 121736 588600
rect 96120 588560 121736 588588
rect 96120 588548 96126 588560
rect 121730 588548 121736 588560
rect 121788 588548 121794 588600
rect 92290 587868 92296 587920
rect 92348 587908 92354 587920
rect 96062 587908 96068 587920
rect 92348 587880 96068 587908
rect 92348 587868 92354 587880
rect 96062 587868 96068 587880
rect 96120 587868 96126 587920
rect 97166 586576 97172 586628
rect 97224 586616 97230 586628
rect 125962 586616 125968 586628
rect 97224 586588 125968 586616
rect 97224 586576 97230 586588
rect 125962 586576 125968 586588
rect 126020 586576 126026 586628
rect 106918 586508 106924 586560
rect 106976 586548 106982 586560
rect 136818 586548 136824 586560
rect 106976 586520 136824 586548
rect 106976 586508 106982 586520
rect 136818 586508 136824 586520
rect 136876 586508 136882 586560
rect 47946 585760 47952 585812
rect 48004 585800 48010 585812
rect 80790 585800 80796 585812
rect 48004 585772 80796 585800
rect 48004 585760 48010 585772
rect 80790 585760 80796 585772
rect 80848 585760 80854 585812
rect 47946 585216 47952 585268
rect 48004 585256 48010 585268
rect 76006 585256 76012 585268
rect 48004 585228 76012 585256
rect 48004 585216 48010 585228
rect 76006 585216 76012 585228
rect 76064 585216 76070 585268
rect 85390 585216 85396 585268
rect 85448 585256 85454 585268
rect 107010 585256 107016 585268
rect 85448 585228 107016 585256
rect 85448 585216 85454 585228
rect 107010 585216 107016 585228
rect 107068 585216 107074 585268
rect 34330 585148 34336 585200
rect 34388 585188 34394 585200
rect 71958 585188 71964 585200
rect 34388 585160 71964 585188
rect 34388 585148 34394 585160
rect 71958 585148 71964 585160
rect 72016 585148 72022 585200
rect 75638 585148 75644 585200
rect 75696 585188 75702 585200
rect 77386 585188 77392 585200
rect 75696 585160 77392 585188
rect 75696 585148 75702 585160
rect 77386 585148 77392 585160
rect 77444 585148 77450 585200
rect 113450 585188 113456 585200
rect 106200 585160 113456 585188
rect 101858 585080 101864 585132
rect 101916 585120 101922 585132
rect 105538 585120 105544 585132
rect 101916 585092 105544 585120
rect 101916 585080 101922 585092
rect 105538 585080 105544 585092
rect 105596 585120 105602 585132
rect 106200 585120 106228 585160
rect 113450 585148 113456 585160
rect 113508 585148 113514 585200
rect 105596 585092 106228 585120
rect 105596 585080 105602 585092
rect 103882 584468 103888 584520
rect 103940 584508 103946 584520
rect 106918 584508 106924 584520
rect 103940 584480 106924 584508
rect 103940 584468 103946 584480
rect 106918 584468 106924 584480
rect 106976 584468 106982 584520
rect 53558 584400 53564 584452
rect 53616 584440 53622 584452
rect 81434 584440 81440 584452
rect 53616 584412 81440 584440
rect 53616 584400 53622 584412
rect 81434 584400 81440 584412
rect 81492 584400 81498 584452
rect 69658 584332 69664 584384
rect 69716 584372 69722 584384
rect 70302 584372 70308 584384
rect 69716 584344 70308 584372
rect 69716 584332 69722 584344
rect 70302 584332 70308 584344
rect 70360 584332 70366 584384
rect 94866 584196 94872 584248
rect 94924 584236 94930 584248
rect 97166 584236 97172 584248
rect 94924 584208 97172 584236
rect 94924 584196 94930 584208
rect 97166 584196 97172 584208
rect 97224 584196 97230 584248
rect 89622 583992 89628 584044
rect 89680 584032 89686 584044
rect 123110 584032 123116 584044
rect 89680 584004 123116 584032
rect 89680 583992 89686 584004
rect 123110 583992 123116 584004
rect 123168 583992 123174 584044
rect 105722 583924 105728 583976
rect 105780 583964 105786 583976
rect 118694 583964 118700 583976
rect 105780 583936 118700 583964
rect 105780 583924 105786 583936
rect 118694 583924 118700 583936
rect 118752 583924 118758 583976
rect 70302 583856 70308 583908
rect 70360 583896 70366 583908
rect 77386 583896 77392 583908
rect 70360 583868 77392 583896
rect 70360 583856 70366 583868
rect 77386 583856 77392 583868
rect 77444 583856 77450 583908
rect 96522 583856 96528 583908
rect 96580 583896 96586 583908
rect 114646 583896 114652 583908
rect 96580 583868 114652 583896
rect 96580 583856 96586 583868
rect 114646 583856 114652 583868
rect 114704 583856 114710 583908
rect 56410 583788 56416 583840
rect 56468 583828 56474 583840
rect 83366 583828 83372 583840
rect 56468 583800 83372 583828
rect 56468 583788 56474 583800
rect 83366 583788 83372 583800
rect 83424 583828 83430 583840
rect 84102 583828 84108 583840
rect 83424 583800 84108 583828
rect 83424 583788 83430 583800
rect 84102 583788 84108 583800
rect 84160 583788 84166 583840
rect 96154 583788 96160 583840
rect 96212 583828 96218 583840
rect 128630 583828 128636 583840
rect 96212 583800 128636 583828
rect 96212 583788 96218 583800
rect 128630 583788 128636 583800
rect 128688 583788 128694 583840
rect 49418 583720 49424 583772
rect 49476 583760 49482 583772
rect 76742 583760 76748 583772
rect 49476 583732 76748 583760
rect 49476 583720 49482 583732
rect 76742 583720 76748 583732
rect 76800 583720 76806 583772
rect 102594 583720 102600 583772
rect 102652 583760 102658 583772
rect 103422 583760 103428 583772
rect 102652 583732 103428 583760
rect 102652 583720 102658 583732
rect 103422 583720 103428 583732
rect 103480 583760 103486 583772
rect 106918 583760 106924 583772
rect 103480 583732 106924 583760
rect 103480 583720 103486 583732
rect 106918 583720 106924 583732
rect 106976 583720 106982 583772
rect 118694 583652 118700 583704
rect 118752 583692 118758 583704
rect 119522 583692 119528 583704
rect 118752 583664 119528 583692
rect 118752 583652 118758 583664
rect 119522 583652 119528 583664
rect 119580 583692 119586 583704
rect 125686 583692 125692 583704
rect 119580 583664 125692 583692
rect 119580 583652 119586 583664
rect 125686 583652 125692 583664
rect 125744 583652 125750 583704
rect 80698 582972 80704 583024
rect 80756 583012 80762 583024
rect 87690 583012 87696 583024
rect 80756 582984 87696 583012
rect 80756 582972 80762 582984
rect 87690 582972 87696 582984
rect 87748 582972 87754 583024
rect 56226 582564 56232 582616
rect 56284 582604 56290 582616
rect 85114 582604 85120 582616
rect 56284 582576 85120 582604
rect 56284 582564 56290 582576
rect 85114 582564 85120 582576
rect 85172 582564 85178 582616
rect 53466 582496 53472 582548
rect 53524 582536 53530 582548
rect 86218 582536 86224 582548
rect 53524 582508 86224 582536
rect 53524 582496 53530 582508
rect 86218 582496 86224 582508
rect 86276 582496 86282 582548
rect 91002 582496 91008 582548
rect 91060 582536 91066 582548
rect 107102 582536 107108 582548
rect 91060 582508 107108 582536
rect 91060 582496 91066 582508
rect 107102 582496 107108 582508
rect 107160 582496 107166 582548
rect 39666 582428 39672 582480
rect 39724 582468 39730 582480
rect 75730 582468 75736 582480
rect 39724 582440 75736 582468
rect 39724 582428 39730 582440
rect 75730 582428 75736 582440
rect 75788 582428 75794 582480
rect 87690 582428 87696 582480
rect 87748 582468 87754 582480
rect 113358 582468 113364 582480
rect 87748 582440 113364 582468
rect 87748 582428 87754 582440
rect 113358 582428 113364 582440
rect 113416 582428 113422 582480
rect 41046 582360 41052 582412
rect 41104 582400 41110 582412
rect 79962 582400 79968 582412
rect 41104 582372 79968 582400
rect 41104 582360 41110 582372
rect 79962 582360 79968 582372
rect 80020 582360 80026 582412
rect 92842 582360 92848 582412
rect 92900 582400 92906 582412
rect 93762 582400 93768 582412
rect 92900 582372 93768 582400
rect 92900 582360 92906 582372
rect 93762 582360 93768 582372
rect 93820 582400 93826 582412
rect 124490 582400 124496 582412
rect 93820 582372 124496 582400
rect 93820 582360 93826 582372
rect 124490 582360 124496 582372
rect 124548 582360 124554 582412
rect 103698 581952 103704 582004
rect 103756 581992 103762 582004
rect 103756 581964 113174 581992
rect 103756 581952 103762 581964
rect 69106 581884 69112 581936
rect 69164 581924 69170 581936
rect 69750 581924 69756 581936
rect 69164 581896 69756 581924
rect 69164 581884 69170 581896
rect 69750 581884 69756 581896
rect 69808 581884 69814 581936
rect 70486 581816 70492 581868
rect 70544 581856 70550 581868
rect 71774 581856 71780 581868
rect 70544 581828 71780 581856
rect 70544 581816 70550 581828
rect 71774 581816 71780 581828
rect 71832 581816 71838 581868
rect 72418 581788 72424 581800
rect 64846 581760 72424 581788
rect 57606 581612 57612 581664
rect 57664 581652 57670 581664
rect 64846 581652 64874 581760
rect 72418 581748 72424 581760
rect 72476 581748 72482 581800
rect 101398 581748 101404 581800
rect 101456 581788 101462 581800
rect 101456 581760 103514 581788
rect 101456 581748 101462 581760
rect 70210 581680 70216 581732
rect 70268 581720 70274 581732
rect 73798 581720 73804 581732
rect 70268 581692 73804 581720
rect 70268 581680 70274 581692
rect 73798 581680 73804 581692
rect 73856 581680 73862 581732
rect 57664 581624 64874 581652
rect 57664 581612 57670 581624
rect 103486 581516 103514 581760
rect 104434 581680 104440 581732
rect 104492 581720 104498 581732
rect 105630 581720 105636 581732
rect 104492 581692 105636 581720
rect 104492 581680 104498 581692
rect 105630 581680 105636 581692
rect 105688 581680 105694 581732
rect 113146 581720 113174 581964
rect 120166 581720 120172 581732
rect 113146 581692 120172 581720
rect 120166 581680 120172 581692
rect 120224 581680 120230 581732
rect 121730 581516 121736 581528
rect 103486 581488 121736 581516
rect 121730 581476 121736 581488
rect 121788 581476 121794 581528
rect 36998 581068 37004 581120
rect 37056 581108 37062 581120
rect 70394 581108 70400 581120
rect 37056 581080 70400 581108
rect 37056 581068 37062 581080
rect 70394 581068 70400 581080
rect 70452 581068 70458 581120
rect 53558 581000 53564 581052
rect 53616 581040 53622 581052
rect 70486 581040 70492 581052
rect 53616 581012 70492 581040
rect 53616 581000 53622 581012
rect 70486 581000 70492 581012
rect 70544 581000 70550 581052
rect 105630 581000 105636 581052
rect 105688 581040 105694 581052
rect 114738 581040 114744 581052
rect 105688 581012 114744 581040
rect 105688 581000 105694 581012
rect 114738 581000 114744 581012
rect 114796 581000 114802 581052
rect 108022 580932 108028 580984
rect 108080 580972 108086 580984
rect 122926 580972 122932 580984
rect 108080 580944 122932 580972
rect 108080 580932 108086 580944
rect 122926 580932 122932 580944
rect 122984 580972 122990 580984
rect 125870 580972 125876 580984
rect 122984 580944 125876 580972
rect 122984 580932 122990 580944
rect 125870 580932 125876 580944
rect 125928 580932 125934 580984
rect 108942 580864 108948 580916
rect 109000 580904 109006 580916
rect 118694 580904 118700 580916
rect 109000 580876 118700 580904
rect 109000 580864 109006 580876
rect 118694 580864 118700 580876
rect 118752 580864 118758 580916
rect 105814 580252 105820 580304
rect 105872 580292 105878 580304
rect 119338 580292 119344 580304
rect 105872 580264 119344 580292
rect 105872 580252 105878 580264
rect 119338 580252 119344 580264
rect 119396 580252 119402 580304
rect 35618 579640 35624 579692
rect 35676 579680 35682 579692
rect 69658 579680 69664 579692
rect 35676 579652 69664 579680
rect 35676 579640 35682 579652
rect 69658 579640 69664 579652
rect 69716 579640 69722 579692
rect 59262 579572 59268 579624
rect 59320 579612 59326 579624
rect 67634 579612 67640 579624
rect 59320 579584 67640 579612
rect 59320 579572 59326 579584
rect 67634 579572 67640 579584
rect 67692 579572 67698 579624
rect 108942 579572 108948 579624
rect 109000 579612 109006 579624
rect 120350 579612 120356 579624
rect 109000 579584 120356 579612
rect 109000 579572 109006 579584
rect 120350 579572 120356 579584
rect 120408 579612 120414 579624
rect 121086 579612 121092 579624
rect 120408 579584 121092 579612
rect 120408 579572 120414 579584
rect 121086 579572 121092 579584
rect 121144 579572 121150 579624
rect 50890 578892 50896 578944
rect 50948 578932 50954 578944
rect 59262 578932 59268 578944
rect 50948 578904 59268 578932
rect 50948 578892 50954 578904
rect 59262 578892 59268 578904
rect 59320 578892 59326 578944
rect 121086 578280 121092 578332
rect 121144 578320 121150 578332
rect 123570 578320 123576 578332
rect 121144 578292 123576 578320
rect 121144 578280 121150 578292
rect 123570 578280 123576 578292
rect 123628 578280 123634 578332
rect 108666 578212 108672 578264
rect 108724 578252 108730 578264
rect 140866 578252 140872 578264
rect 108724 578224 140872 578252
rect 108724 578212 108730 578224
rect 140866 578212 140872 578224
rect 140924 578212 140930 578264
rect 108114 578144 108120 578196
rect 108172 578184 108178 578196
rect 125778 578184 125784 578196
rect 108172 578156 125784 578184
rect 108172 578144 108178 578156
rect 125778 578144 125784 578156
rect 125836 578144 125842 578196
rect 108942 577464 108948 577516
rect 109000 577504 109006 577516
rect 116394 577504 116400 577516
rect 109000 577476 116400 577504
rect 109000 577464 109006 577476
rect 116394 577464 116400 577476
rect 116452 577464 116458 577516
rect 108666 576172 108672 576224
rect 108724 576212 108730 576224
rect 116302 576212 116308 576224
rect 108724 576184 116308 576212
rect 108724 576172 108730 576184
rect 116302 576172 116308 576184
rect 116360 576172 116366 576224
rect 108758 576104 108764 576156
rect 108816 576144 108822 576156
rect 142246 576144 142252 576156
rect 108816 576116 142252 576144
rect 108816 576104 108822 576116
rect 142246 576104 142252 576116
rect 142304 576104 142310 576156
rect 35802 575492 35808 575544
rect 35860 575532 35866 575544
rect 67634 575532 67640 575544
rect 35860 575504 67640 575532
rect 35860 575492 35866 575504
rect 67634 575492 67640 575504
rect 67692 575492 67698 575544
rect 117130 575492 117136 575544
rect 117188 575532 117194 575544
rect 126238 575532 126244 575544
rect 117188 575504 126244 575532
rect 117188 575492 117194 575504
rect 126238 575492 126244 575504
rect 126296 575492 126302 575544
rect 53834 574744 53840 574796
rect 53892 574784 53898 574796
rect 55030 574784 55036 574796
rect 53892 574756 55036 574784
rect 53892 574744 53898 574756
rect 55030 574744 55036 574756
rect 55088 574784 55094 574796
rect 67634 574784 67640 574796
rect 55088 574756 67640 574784
rect 55088 574744 55094 574756
rect 67634 574744 67640 574756
rect 67692 574744 67698 574796
rect 105630 574472 105636 574524
rect 105688 574512 105694 574524
rect 110414 574512 110420 574524
rect 105688 574484 110420 574512
rect 105688 574472 105694 574484
rect 110414 574472 110420 574484
rect 110472 574472 110478 574524
rect 48130 573996 48136 574048
rect 48188 574036 48194 574048
rect 67634 574036 67640 574048
rect 48188 574008 67640 574036
rect 48188 573996 48194 574008
rect 67634 573996 67640 574008
rect 67692 573996 67698 574048
rect 108574 573996 108580 574048
rect 108632 574036 108638 574048
rect 123018 574036 123024 574048
rect 108632 574008 123024 574036
rect 108632 573996 108638 574008
rect 123018 573996 123024 574008
rect 123076 573996 123082 574048
rect 108942 573928 108948 573980
rect 109000 573968 109006 573980
rect 109678 573968 109684 573980
rect 109000 573940 109684 573968
rect 109000 573928 109006 573940
rect 109678 573928 109684 573940
rect 109736 573928 109742 573980
rect 43898 573384 43904 573436
rect 43956 573424 43962 573436
rect 53834 573424 53840 573436
rect 43956 573396 53840 573424
rect 43956 573384 43962 573396
rect 53834 573384 53840 573396
rect 53892 573384 53898 573436
rect 32950 573316 32956 573368
rect 33008 573356 33014 573368
rect 48130 573356 48136 573368
rect 33008 573328 48136 573356
rect 33008 573316 33014 573328
rect 48130 573316 48136 573328
rect 48188 573316 48194 573368
rect 109678 573316 109684 573368
rect 109736 573356 109742 573368
rect 140958 573356 140964 573368
rect 109736 573328 140964 573356
rect 109736 573316 109742 573328
rect 140958 573316 140964 573328
rect 141016 573316 141022 573368
rect 108942 573180 108948 573232
rect 109000 573220 109006 573232
rect 114554 573220 114560 573232
rect 109000 573192 114560 573220
rect 109000 573180 109006 573192
rect 114554 573180 114560 573192
rect 114612 573180 114618 573232
rect 108022 571956 108028 572008
rect 108080 571996 108086 572008
rect 133966 571996 133972 572008
rect 108080 571968 133972 571996
rect 108080 571956 108086 571968
rect 133966 571956 133972 571968
rect 134024 571996 134030 572008
rect 134150 571996 134156 572008
rect 134024 571968 134156 571996
rect 134024 571956 134030 571968
rect 134150 571956 134156 571968
rect 134208 571956 134214 572008
rect 65886 571752 65892 571804
rect 65944 571792 65950 571804
rect 66070 571792 66076 571804
rect 65944 571764 66076 571792
rect 65944 571752 65950 571764
rect 66070 571752 66076 571764
rect 66128 571792 66134 571804
rect 67634 571792 67640 571804
rect 66128 571764 67640 571792
rect 66128 571752 66134 571764
rect 67634 571752 67640 571764
rect 67692 571752 67698 571804
rect 64506 571276 64512 571328
rect 64564 571316 64570 571328
rect 65886 571316 65892 571328
rect 64564 571288 65892 571316
rect 64564 571276 64570 571288
rect 65886 571276 65892 571288
rect 65944 571316 65950 571328
rect 67726 571316 67732 571328
rect 65944 571288 67732 571316
rect 65944 571276 65950 571288
rect 67726 571276 67732 571288
rect 67784 571276 67790 571328
rect 108298 571276 108304 571328
rect 108356 571316 108362 571328
rect 128446 571316 128452 571328
rect 108356 571288 128452 571316
rect 108356 571276 108362 571288
rect 128446 571276 128452 571288
rect 128504 571276 128510 571328
rect 63218 571208 63224 571260
rect 63276 571248 63282 571260
rect 67634 571248 67640 571260
rect 63276 571220 67640 571248
rect 63276 571208 63282 571220
rect 67634 571208 67640 571220
rect 67692 571208 67698 571260
rect 66162 569848 66168 569900
rect 66220 569888 66226 569900
rect 66990 569888 66996 569900
rect 66220 569860 66996 569888
rect 66220 569848 66226 569860
rect 66990 569848 66996 569860
rect 67048 569848 67054 569900
rect 66990 568896 66996 568948
rect 67048 568936 67054 568948
rect 67818 568936 67824 568948
rect 67048 568908 67824 568936
rect 67048 568896 67054 568908
rect 67818 568896 67824 568908
rect 67876 568896 67882 568948
rect 63218 568624 63224 568676
rect 63276 568664 63282 568676
rect 67358 568664 67364 568676
rect 63276 568636 67364 568664
rect 63276 568624 63282 568636
rect 67358 568624 67364 568636
rect 67416 568664 67422 568676
rect 67634 568664 67640 568676
rect 67416 568636 67640 568664
rect 67416 568624 67422 568636
rect 67634 568624 67640 568636
rect 67692 568624 67698 568676
rect 108942 568556 108948 568608
rect 109000 568596 109006 568608
rect 118602 568596 118608 568608
rect 109000 568568 118608 568596
rect 109000 568556 109006 568568
rect 118602 568556 118608 568568
rect 118660 568556 118666 568608
rect 108850 568488 108856 568540
rect 108908 568528 108914 568540
rect 124398 568528 124404 568540
rect 108908 568500 124404 568528
rect 108908 568488 108914 568500
rect 124398 568488 124404 568500
rect 124456 568528 124462 568540
rect 125502 568528 125508 568540
rect 124456 568500 125508 568528
rect 124456 568488 124462 568500
rect 125502 568488 125508 568500
rect 125560 568488 125566 568540
rect 65978 568216 65984 568268
rect 66036 568256 66042 568268
rect 67634 568256 67640 568268
rect 66036 568228 67640 568256
rect 66036 568216 66042 568228
rect 67634 568216 67640 568228
rect 67692 568216 67698 568268
rect 42794 567808 42800 567860
rect 42852 567848 42858 567860
rect 43714 567848 43720 567860
rect 42852 567820 43720 567848
rect 42852 567808 42858 567820
rect 43714 567808 43720 567820
rect 43772 567848 43778 567860
rect 67634 567848 67640 567860
rect 43772 567820 67640 567848
rect 43772 567808 43778 567820
rect 67634 567808 67640 567820
rect 67692 567808 67698 567860
rect 125502 567808 125508 567860
rect 125560 567848 125566 567860
rect 132586 567848 132592 567860
rect 125560 567820 132592 567848
rect 125560 567808 125566 567820
rect 132586 567808 132592 567820
rect 132644 567808 132650 567860
rect 30282 567196 30288 567248
rect 30340 567236 30346 567248
rect 42794 567236 42800 567248
rect 30340 567208 42800 567236
rect 30340 567196 30346 567208
rect 42794 567196 42800 567208
rect 42852 567196 42858 567248
rect 60458 567196 60464 567248
rect 60516 567236 60522 567248
rect 65978 567236 65984 567248
rect 60516 567208 65984 567236
rect 60516 567196 60522 567208
rect 65978 567196 65984 567208
rect 66036 567196 66042 567248
rect 108942 567196 108948 567248
rect 109000 567236 109006 567248
rect 110506 567236 110512 567248
rect 109000 567208 110512 567236
rect 109000 567196 109006 567208
rect 110506 567196 110512 567208
rect 110564 567236 110570 567248
rect 113542 567236 113548 567248
rect 110564 567208 113548 567236
rect 110564 567196 110570 567208
rect 113542 567196 113548 567208
rect 113600 567196 113606 567248
rect 61930 566448 61936 566500
rect 61988 566488 61994 566500
rect 67634 566488 67640 566500
rect 61988 566460 67640 566488
rect 61988 566448 61994 566460
rect 67634 566448 67640 566460
rect 67692 566448 67698 566500
rect 108942 566448 108948 566500
rect 109000 566488 109006 566500
rect 128538 566488 128544 566500
rect 109000 566460 128544 566488
rect 109000 566448 109006 566460
rect 128538 566448 128544 566460
rect 128596 566448 128602 566500
rect 135162 566448 135168 566500
rect 135220 566488 135226 566500
rect 142154 566488 142160 566500
rect 135220 566460 142160 566488
rect 135220 566448 135226 566460
rect 142154 566448 142160 566460
rect 142212 566448 142218 566500
rect 3234 565836 3240 565888
rect 3292 565876 3298 565888
rect 25498 565876 25504 565888
rect 3292 565848 25504 565876
rect 3292 565836 3298 565848
rect 25498 565836 25504 565848
rect 25556 565836 25562 565888
rect 108942 565836 108948 565888
rect 109000 565876 109006 565888
rect 134518 565876 134524 565888
rect 109000 565848 134524 565876
rect 109000 565836 109006 565848
rect 134518 565836 134524 565848
rect 134576 565876 134582 565888
rect 135162 565876 135168 565888
rect 134576 565848 135168 565876
rect 134576 565836 134582 565848
rect 135162 565836 135168 565848
rect 135220 565836 135226 565888
rect 108850 565768 108856 565820
rect 108908 565808 108914 565820
rect 117406 565808 117412 565820
rect 108908 565780 117412 565808
rect 108908 565768 108914 565780
rect 117406 565768 117412 565780
rect 117464 565768 117470 565820
rect 44082 565088 44088 565140
rect 44140 565128 44146 565140
rect 66898 565128 66904 565140
rect 44140 565100 66904 565128
rect 44140 565088 44146 565100
rect 66898 565088 66904 565100
rect 66956 565128 66962 565140
rect 67634 565128 67640 565140
rect 66956 565100 67640 565128
rect 66956 565088 66962 565100
rect 67634 565088 67640 565100
rect 67692 565088 67698 565140
rect 126238 565088 126244 565140
rect 126296 565128 126302 565140
rect 497458 565128 497464 565140
rect 126296 565100 497464 565128
rect 126296 565088 126302 565100
rect 497458 565088 497464 565100
rect 497516 565128 497522 565140
rect 504358 565128 504364 565140
rect 497516 565100 504364 565128
rect 497516 565088 497522 565100
rect 504358 565088 504364 565100
rect 504416 565088 504422 565140
rect 67634 564448 67640 564460
rect 64846 564420 67640 564448
rect 42702 564340 42708 564392
rect 42760 564380 42766 564392
rect 63494 564380 63500 564392
rect 42760 564352 63500 564380
rect 42760 564340 42766 564352
rect 63494 564340 63500 564352
rect 63552 564380 63558 564392
rect 64846 564380 64874 564420
rect 67634 564408 67640 564420
rect 67692 564408 67698 564460
rect 117406 564408 117412 564460
rect 117464 564448 117470 564460
rect 119430 564448 119436 564460
rect 117464 564420 119436 564448
rect 117464 564408 117470 564420
rect 119430 564408 119436 564420
rect 119488 564408 119494 564460
rect 63552 564352 64874 564380
rect 63552 564340 63558 564352
rect 52362 564272 52368 564324
rect 52420 564312 52426 564324
rect 67634 564312 67640 564324
rect 52420 564284 67640 564312
rect 52420 564272 52426 564284
rect 67634 564272 67640 564284
rect 67692 564272 67698 564324
rect 61838 564204 61844 564256
rect 61896 564244 61902 564256
rect 67726 564244 67732 564256
rect 61896 564216 67732 564244
rect 61896 564204 61902 564216
rect 67726 564204 67732 564216
rect 67784 564204 67790 564256
rect 111702 564136 111708 564188
rect 111760 564176 111766 564188
rect 113358 564176 113364 564188
rect 111760 564148 113364 564176
rect 111760 564136 111766 564148
rect 113358 564136 113364 564148
rect 113416 564136 113422 564188
rect 111150 563796 111156 563848
rect 111208 563836 111214 563848
rect 114738 563836 114744 563848
rect 111208 563808 114744 563836
rect 111208 563796 111214 563808
rect 114738 563796 114744 563808
rect 114796 563796 114802 563848
rect 111242 563660 111248 563712
rect 111300 563700 111306 563712
rect 116210 563700 116216 563712
rect 111300 563672 116216 563700
rect 111300 563660 111306 563672
rect 116210 563660 116216 563672
rect 116268 563660 116274 563712
rect 504358 563660 504364 563712
rect 504416 563700 504422 563712
rect 580166 563700 580172 563712
rect 504416 563672 580172 563700
rect 504416 563660 504422 563672
rect 580166 563660 580172 563672
rect 580224 563660 580230 563712
rect 108942 563456 108948 563508
rect 109000 563496 109006 563508
rect 111058 563496 111064 563508
rect 109000 563468 111064 563496
rect 109000 563456 109006 563468
rect 111058 563456 111064 563468
rect 111116 563496 111122 563508
rect 113818 563496 113824 563508
rect 111116 563468 113824 563496
rect 111116 563456 111122 563468
rect 113818 563456 113824 563468
rect 113876 563456 113882 563508
rect 60274 563184 60280 563236
rect 60332 563224 60338 563236
rect 60642 563224 60648 563236
rect 60332 563196 60648 563224
rect 60332 563184 60338 563196
rect 60642 563184 60648 563196
rect 60700 563184 60706 563236
rect 60550 563116 60556 563168
rect 60608 563156 60614 563168
rect 61378 563156 61384 563168
rect 60608 563128 61384 563156
rect 60608 563116 60614 563128
rect 61378 563116 61384 563128
rect 61436 563116 61442 563168
rect 49510 563048 49516 563100
rect 49568 563088 49574 563100
rect 52362 563088 52368 563100
rect 49568 563060 52368 563088
rect 49568 563048 49574 563060
rect 52362 563048 52368 563060
rect 52420 563048 52426 563100
rect 60642 563048 60648 563100
rect 60700 563088 60706 563100
rect 61838 563088 61844 563100
rect 60700 563060 61844 563088
rect 60700 563048 60706 563060
rect 61838 563048 61844 563060
rect 61896 563048 61902 563100
rect 53650 562300 53656 562352
rect 53708 562340 53714 562352
rect 54478 562340 54484 562352
rect 53708 562312 54484 562340
rect 53708 562300 53714 562312
rect 54478 562300 54484 562312
rect 54536 562340 54542 562352
rect 67634 562340 67640 562352
rect 54536 562312 67640 562340
rect 54536 562300 54542 562312
rect 67634 562300 67640 562312
rect 67692 562300 67698 562352
rect 108942 562300 108948 562352
rect 109000 562340 109006 562352
rect 142154 562340 142160 562352
rect 109000 562312 142160 562340
rect 109000 562300 109006 562312
rect 142154 562300 142160 562312
rect 142212 562340 142218 562352
rect 146294 562340 146300 562352
rect 142212 562312 146300 562340
rect 142212 562300 142218 562312
rect 146294 562300 146300 562312
rect 146352 562300 146358 562352
rect 48130 561620 48136 561672
rect 48188 561660 48194 561672
rect 50798 561660 50804 561672
rect 48188 561632 50804 561660
rect 48188 561620 48194 561632
rect 50798 561620 50804 561632
rect 50856 561660 50862 561672
rect 67726 561660 67732 561672
rect 50856 561632 67732 561660
rect 50856 561620 50862 561632
rect 67726 561620 67732 561632
rect 67784 561620 67790 561672
rect 135898 561620 135904 561672
rect 135956 561660 135962 561672
rect 136726 561660 136732 561672
rect 135956 561632 136732 561660
rect 135956 561620 135962 561632
rect 136726 561620 136732 561632
rect 136784 561620 136790 561672
rect 58986 561552 58992 561604
rect 59044 561592 59050 561604
rect 60274 561592 60280 561604
rect 59044 561564 60280 561592
rect 59044 561552 59050 561564
rect 60274 561552 60280 561564
rect 60332 561592 60338 561604
rect 67634 561592 67640 561604
rect 60332 561564 67640 561592
rect 60332 561552 60338 561564
rect 67634 561552 67640 561564
rect 67692 561552 67698 561604
rect 108942 561008 108948 561060
rect 109000 561048 109006 561060
rect 111794 561048 111800 561060
rect 109000 561020 111800 561048
rect 109000 561008 109006 561020
rect 111794 561008 111800 561020
rect 111852 561048 111858 561060
rect 117498 561048 117504 561060
rect 111852 561020 117504 561048
rect 111852 561008 111858 561020
rect 117498 561008 117504 561020
rect 117556 561008 117562 561060
rect 108850 560940 108856 560992
rect 108908 560980 108914 560992
rect 135898 560980 135904 560992
rect 108908 560952 135904 560980
rect 108908 560940 108914 560952
rect 135898 560940 135904 560952
rect 135956 560940 135962 560992
rect 59078 560192 59084 560244
rect 59136 560232 59142 560244
rect 59262 560232 59268 560244
rect 59136 560204 59268 560232
rect 59136 560192 59142 560204
rect 59262 560192 59268 560204
rect 59320 560232 59326 560244
rect 67634 560232 67640 560244
rect 59320 560204 67640 560232
rect 59320 560192 59326 560204
rect 67634 560192 67640 560204
rect 67692 560192 67698 560244
rect 112898 559580 112904 559632
rect 112956 559620 112962 559632
rect 131298 559620 131304 559632
rect 112956 559592 131304 559620
rect 112956 559580 112962 559592
rect 131298 559580 131304 559592
rect 131356 559580 131362 559632
rect 42610 559512 42616 559564
rect 42668 559552 42674 559564
rect 59262 559552 59268 559564
rect 42668 559524 59268 559552
rect 42668 559512 42674 559524
rect 59262 559512 59268 559524
rect 59320 559512 59326 559564
rect 108942 559512 108948 559564
rect 109000 559552 109006 559564
rect 132494 559552 132500 559564
rect 109000 559524 132500 559552
rect 109000 559512 109006 559524
rect 132494 559512 132500 559524
rect 132552 559552 132558 559564
rect 132770 559552 132776 559564
rect 132552 559524 132776 559552
rect 132552 559512 132558 559524
rect 132770 559512 132776 559524
rect 132828 559512 132834 559564
rect 56410 558832 56416 558884
rect 56468 558872 56474 558884
rect 58710 558872 58716 558884
rect 56468 558844 58716 558872
rect 56468 558832 56474 558844
rect 58710 558832 58716 558844
rect 58768 558832 58774 558884
rect 63402 558832 63408 558884
rect 63460 558872 63466 558884
rect 64138 558872 64144 558884
rect 63460 558844 64144 558872
rect 63460 558832 63466 558844
rect 64138 558832 64144 558844
rect 64196 558832 64202 558884
rect 108022 558832 108028 558884
rect 108080 558872 108086 558884
rect 139394 558872 139400 558884
rect 108080 558844 139400 558872
rect 108080 558832 108086 558844
rect 139394 558832 139400 558844
rect 139452 558832 139458 558884
rect 107746 558764 107752 558816
rect 107804 558804 107810 558816
rect 111886 558804 111892 558816
rect 107804 558776 111892 558804
rect 107804 558764 107810 558776
rect 111886 558764 111892 558776
rect 111944 558764 111950 558816
rect 108942 558152 108948 558204
rect 109000 558192 109006 558204
rect 121638 558192 121644 558204
rect 109000 558164 121644 558192
rect 109000 558152 109006 558164
rect 121638 558152 121644 558164
rect 121696 558152 121702 558204
rect 64138 557608 64144 557660
rect 64196 557648 64202 557660
rect 67634 557648 67640 557660
rect 64196 557620 67640 557648
rect 64196 557608 64202 557620
rect 67634 557608 67640 557620
rect 67692 557608 67698 557660
rect 50338 557580 50344 557592
rect 49528 557552 50344 557580
rect 39942 557404 39948 557456
rect 40000 557444 40006 557456
rect 49528 557444 49556 557552
rect 50338 557540 50344 557552
rect 50396 557580 50402 557592
rect 67726 557580 67732 557592
rect 50396 557552 67732 557580
rect 50396 557540 50402 557552
rect 67726 557540 67732 557552
rect 67784 557540 67790 557592
rect 49602 557472 49608 557524
rect 49660 557512 49666 557524
rect 67818 557512 67824 557524
rect 49660 557484 67824 557512
rect 49660 557472 49666 557484
rect 67818 557472 67824 557484
rect 67876 557472 67882 557524
rect 40000 557416 49556 557444
rect 40000 557404 40006 557416
rect 56502 557404 56508 557456
rect 56560 557444 56566 557456
rect 67634 557444 67640 557456
rect 56560 557416 67640 557444
rect 56560 557404 56566 557416
rect 67634 557404 67640 557416
rect 67692 557404 67698 557456
rect 108942 557132 108948 557184
rect 109000 557172 109006 557184
rect 110598 557172 110604 557184
rect 109000 557144 110604 557172
rect 109000 557132 109006 557144
rect 110598 557132 110604 557144
rect 110656 557132 110662 557184
rect 34238 556860 34244 556912
rect 34296 556900 34302 556912
rect 49602 556900 49608 556912
rect 34296 556872 49608 556900
rect 34296 556860 34302 556872
rect 49602 556860 49608 556872
rect 49660 556860 49666 556912
rect 39850 556792 39856 556844
rect 39908 556832 39914 556844
rect 56502 556832 56508 556844
rect 39908 556804 56508 556832
rect 39908 556792 39914 556804
rect 56502 556792 56508 556804
rect 56560 556792 56566 556844
rect 110598 556792 110604 556844
rect 110656 556832 110662 556844
rect 141050 556832 141056 556844
rect 110656 556804 141056 556832
rect 110656 556792 110662 556804
rect 141050 556792 141056 556804
rect 141108 556792 141114 556844
rect 56502 556180 56508 556232
rect 56560 556220 56566 556232
rect 58618 556220 58624 556232
rect 56560 556192 58624 556220
rect 56560 556180 56566 556192
rect 58618 556180 58624 556192
rect 58676 556180 58682 556232
rect 58636 556152 58664 556180
rect 67726 556152 67732 556164
rect 58636 556124 67732 556152
rect 67726 556112 67732 556124
rect 67784 556112 67790 556164
rect 112990 555500 112996 555552
rect 113048 555540 113054 555552
rect 119522 555540 119528 555552
rect 113048 555512 119528 555540
rect 113048 555500 113054 555512
rect 119522 555500 119528 555512
rect 119580 555500 119586 555552
rect 113082 555432 113088 555484
rect 113140 555472 113146 555484
rect 113542 555472 113548 555484
rect 113140 555444 113548 555472
rect 113140 555432 113146 555444
rect 113542 555432 113548 555444
rect 113600 555432 113606 555484
rect 109770 555364 109776 555416
rect 109828 555404 109834 555416
rect 121730 555404 121736 555416
rect 109828 555376 121736 555404
rect 109828 555364 109834 555376
rect 121730 555364 121736 555376
rect 121788 555364 121794 555416
rect 105630 555092 105636 555144
rect 105688 555132 105694 555144
rect 105814 555132 105820 555144
rect 105688 555104 105820 555132
rect 105688 555092 105694 555104
rect 105814 555092 105820 555104
rect 105872 555092 105878 555144
rect 67634 554792 67640 554804
rect 62132 554764 67640 554792
rect 62132 554736 62160 554764
rect 67634 554752 67640 554764
rect 67692 554752 67698 554804
rect 108850 554752 108856 554804
rect 108908 554792 108914 554804
rect 113266 554792 113272 554804
rect 108908 554764 113272 554792
rect 108908 554752 108914 554764
rect 113266 554752 113272 554764
rect 113324 554792 113330 554804
rect 114094 554792 114100 554804
rect 113324 554764 114100 554792
rect 113324 554752 113330 554764
rect 114094 554752 114100 554764
rect 114152 554752 114158 554804
rect 41230 554684 41236 554736
rect 41288 554724 41294 554736
rect 62114 554724 62120 554736
rect 41288 554696 62120 554724
rect 41288 554684 41294 554696
rect 62114 554684 62120 554696
rect 62172 554684 62178 554736
rect 108942 554684 108948 554736
rect 109000 554724 109006 554736
rect 129826 554724 129832 554736
rect 109000 554696 129832 554724
rect 109000 554684 109006 554696
rect 129826 554684 129832 554696
rect 129884 554684 129890 554736
rect 45462 554616 45468 554668
rect 45520 554656 45526 554668
rect 48038 554656 48044 554668
rect 45520 554628 48044 554656
rect 45520 554616 45526 554628
rect 48038 554616 48044 554628
rect 48096 554656 48102 554668
rect 67634 554656 67640 554668
rect 48096 554628 67640 554656
rect 48096 554616 48102 554628
rect 67634 554616 67640 554628
rect 67692 554616 67698 554668
rect 129826 554072 129832 554124
rect 129884 554112 129890 554124
rect 136726 554112 136732 554124
rect 129884 554084 136732 554112
rect 129884 554072 129890 554084
rect 136726 554072 136732 554084
rect 136784 554072 136790 554124
rect 108942 554004 108948 554056
rect 109000 554044 109006 554056
rect 133966 554044 133972 554056
rect 109000 554016 133972 554044
rect 109000 554004 109006 554016
rect 133966 554004 133972 554016
rect 134024 554004 134030 554056
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 40678 553432 40684 553444
rect 3384 553404 40684 553432
rect 3384 553392 3390 553404
rect 40678 553392 40684 553404
rect 40736 553392 40742 553444
rect 67910 553432 67916 553444
rect 57624 553404 67916 553432
rect 57624 553376 57652 553404
rect 67910 553392 67916 553404
rect 67968 553392 67974 553444
rect 114094 553392 114100 553444
rect 114152 553432 114158 553444
rect 116578 553432 116584 553444
rect 114152 553404 116584 553432
rect 114152 553392 114158 553404
rect 116578 553392 116584 553404
rect 116636 553392 116642 553444
rect 57606 553324 57612 553376
rect 57664 553324 57670 553376
rect 57238 552644 57244 552696
rect 57296 552684 57302 552696
rect 57882 552684 57888 552696
rect 57296 552656 57888 552684
rect 57296 552644 57302 552656
rect 57882 552644 57888 552656
rect 57940 552684 57946 552696
rect 67634 552684 67640 552696
rect 57940 552656 67640 552684
rect 57940 552644 57946 552656
rect 67634 552644 67640 552656
rect 67692 552644 67698 552696
rect 130194 552644 130200 552696
rect 130252 552684 130258 552696
rect 138014 552684 138020 552696
rect 130252 552656 138020 552684
rect 130252 552644 130258 552656
rect 138014 552644 138020 552656
rect 138072 552644 138078 552696
rect 108942 552032 108948 552084
rect 109000 552072 109006 552084
rect 130010 552072 130016 552084
rect 109000 552044 130016 552072
rect 109000 552032 109006 552044
rect 130010 552032 130016 552044
rect 130068 552072 130074 552084
rect 130194 552072 130200 552084
rect 130068 552044 130200 552072
rect 130068 552032 130074 552044
rect 130194 552032 130200 552044
rect 130252 552032 130258 552084
rect 64782 551964 64788 552016
rect 64840 552004 64846 552016
rect 65610 552004 65616 552016
rect 64840 551976 65616 552004
rect 64840 551964 64846 551976
rect 65610 551964 65616 551976
rect 65668 552004 65674 552016
rect 67634 552004 67640 552016
rect 65668 551976 67640 552004
rect 65668 551964 65674 551976
rect 67634 551964 67640 551976
rect 67692 551964 67698 552016
rect 108298 551964 108304 552016
rect 108356 552004 108362 552016
rect 143626 552004 143632 552016
rect 108356 551976 143632 552004
rect 108356 551964 108362 551976
rect 143626 551964 143632 551976
rect 143684 551964 143690 552016
rect 112622 551352 112628 551404
rect 112680 551392 112686 551404
rect 116118 551392 116124 551404
rect 112680 551364 116124 551392
rect 112680 551352 112686 551364
rect 116118 551352 116124 551364
rect 116176 551352 116182 551404
rect 109678 551284 109684 551336
rect 109736 551324 109742 551336
rect 117590 551324 117596 551336
rect 109736 551296 117596 551324
rect 109736 551284 109742 551296
rect 117590 551284 117596 551296
rect 117648 551284 117654 551336
rect 106734 551216 106740 551268
rect 106792 551256 106798 551268
rect 111978 551256 111984 551268
rect 106792 551228 111984 551256
rect 106792 551216 106798 551228
rect 111978 551216 111984 551228
rect 112036 551216 112042 551268
rect 108942 550604 108948 550656
rect 109000 550644 109006 550656
rect 109000 550616 110460 550644
rect 109000 550604 109006 550616
rect 59262 550536 59268 550588
rect 59320 550576 59326 550588
rect 64598 550576 64604 550588
rect 59320 550548 64604 550576
rect 59320 550536 59326 550548
rect 64598 550536 64604 550548
rect 64656 550576 64662 550588
rect 67634 550576 67640 550588
rect 64656 550548 67640 550576
rect 64656 550536 64662 550548
rect 67634 550536 67640 550548
rect 67692 550536 67698 550588
rect 110432 550576 110460 550616
rect 111058 550576 111064 550588
rect 110432 550548 111064 550576
rect 111058 550536 111064 550548
rect 111116 550576 111122 550588
rect 115934 550576 115940 550588
rect 111116 550548 115940 550576
rect 111116 550536 111122 550548
rect 115934 550536 115940 550548
rect 115992 550536 115998 550588
rect 63126 549176 63132 549228
rect 63184 549216 63190 549228
rect 63402 549216 63408 549228
rect 63184 549188 63408 549216
rect 63184 549176 63190 549188
rect 63402 549176 63408 549188
rect 63460 549176 63466 549228
rect 108942 549176 108948 549228
rect 109000 549216 109006 549228
rect 132862 549216 132868 549228
rect 109000 549188 132868 549216
rect 109000 549176 109006 549188
rect 132862 549176 132868 549188
rect 132920 549216 132926 549228
rect 133782 549216 133788 549228
rect 132920 549188 133788 549216
rect 132920 549176 132926 549188
rect 133782 549176 133788 549188
rect 133840 549176 133846 549228
rect 109862 549108 109868 549160
rect 109920 549148 109926 549160
rect 111150 549148 111156 549160
rect 109920 549120 111156 549148
rect 109920 549108 109926 549120
rect 111150 549108 111156 549120
rect 111208 549108 111214 549160
rect 63402 548564 63408 548616
rect 63460 548604 63466 548616
rect 67634 548604 67640 548616
rect 63460 548576 67640 548604
rect 63460 548564 63466 548576
rect 67634 548564 67640 548576
rect 67692 548564 67698 548616
rect 133782 548564 133788 548616
rect 133840 548604 133846 548616
rect 142338 548604 142344 548616
rect 133840 548576 142344 548604
rect 133840 548564 133846 548576
rect 142338 548564 142344 548576
rect 142396 548564 142402 548616
rect 108850 548496 108856 548548
rect 108908 548536 108914 548548
rect 138658 548536 138664 548548
rect 108908 548508 138664 548536
rect 108908 548496 108914 548508
rect 138658 548496 138664 548508
rect 138716 548536 138722 548548
rect 143534 548536 143540 548548
rect 138716 548508 143540 548536
rect 138716 548496 138722 548508
rect 143534 548496 143540 548508
rect 143592 548496 143598 548548
rect 41138 547884 41144 547936
rect 41196 547924 41202 547936
rect 67726 547924 67732 547936
rect 41196 547896 67732 547924
rect 41196 547884 41202 547896
rect 67726 547884 67732 547896
rect 67784 547884 67790 547936
rect 108942 547136 108948 547188
rect 109000 547176 109006 547188
rect 135254 547176 135260 547188
rect 109000 547148 135260 547176
rect 109000 547136 109006 547148
rect 135254 547136 135260 547148
rect 135312 547136 135318 547188
rect 62022 546592 62028 546644
rect 62080 546632 62086 546644
rect 64782 546632 64788 546644
rect 62080 546604 64788 546632
rect 62080 546592 62086 546604
rect 64782 546592 64788 546604
rect 64840 546632 64846 546644
rect 67634 546632 67640 546644
rect 64840 546604 67640 546632
rect 64840 546592 64846 546604
rect 67634 546592 67640 546604
rect 67692 546592 67698 546644
rect 60734 546456 60740 546508
rect 60792 546496 60798 546508
rect 67634 546496 67640 546508
rect 60792 546468 67640 546496
rect 60792 546456 60798 546468
rect 67634 546456 67640 546468
rect 67692 546456 67698 546508
rect 108942 545640 108948 545692
rect 109000 545680 109006 545692
rect 115198 545680 115204 545692
rect 109000 545652 115204 545680
rect 109000 545640 109006 545652
rect 115198 545640 115204 545652
rect 115256 545640 115262 545692
rect 38378 545096 38384 545148
rect 38436 545136 38442 545148
rect 65978 545136 65984 545148
rect 38436 545108 65984 545136
rect 38436 545096 38442 545108
rect 65978 545096 65984 545108
rect 66036 545136 66042 545148
rect 67634 545136 67640 545148
rect 66036 545108 67640 545136
rect 66036 545096 66042 545108
rect 67634 545096 67640 545108
rect 67692 545096 67698 545148
rect 25498 545028 25504 545080
rect 25556 545068 25562 545080
rect 68554 545068 68560 545080
rect 25556 545040 68560 545068
rect 25556 545028 25562 545040
rect 68554 545028 68560 545040
rect 68612 545028 68618 545080
rect 108942 544416 108948 544468
rect 109000 544456 109006 544468
rect 116026 544456 116032 544468
rect 109000 544428 116032 544456
rect 109000 544416 109006 544428
rect 116026 544416 116032 544428
rect 116084 544416 116090 544468
rect 108850 544348 108856 544400
rect 108908 544388 108914 544400
rect 139578 544388 139584 544400
rect 108908 544360 139584 544388
rect 108908 544348 108914 544360
rect 139578 544348 139584 544360
rect 139636 544348 139642 544400
rect 108850 543736 108856 543788
rect 108908 543776 108914 543788
rect 109402 543776 109408 543788
rect 108908 543748 109408 543776
rect 108908 543736 108914 543748
rect 109402 543736 109408 543748
rect 109460 543776 109466 543788
rect 113266 543776 113272 543788
rect 109460 543748 113272 543776
rect 109460 543736 109466 543748
rect 113266 543736 113272 543748
rect 113324 543736 113330 543788
rect 139578 543736 139584 543788
rect 139636 543776 139642 543788
rect 140774 543776 140780 543788
rect 139636 543748 140780 543776
rect 139636 543736 139642 543748
rect 140774 543736 140780 543748
rect 140832 543736 140838 543788
rect 60642 543668 60648 543720
rect 60700 543708 60706 543720
rect 61746 543708 61752 543720
rect 60700 543680 61752 543708
rect 60700 543668 60706 543680
rect 61746 543668 61752 543680
rect 61804 543708 61810 543720
rect 67726 543708 67732 543720
rect 61804 543680 67732 543708
rect 61804 543668 61810 543680
rect 67726 543668 67732 543680
rect 67784 543668 67790 543720
rect 108942 543668 108948 543720
rect 109000 543708 109006 543720
rect 129918 543708 129924 543720
rect 109000 543680 129924 543708
rect 109000 543668 109006 543680
rect 129918 543668 129924 543680
rect 129976 543708 129982 543720
rect 130746 543708 130752 543720
rect 129976 543680 130752 543708
rect 129976 543668 129982 543680
rect 130746 543668 130752 543680
rect 130804 543668 130810 543720
rect 60734 542988 60740 543040
rect 60792 543028 60798 543040
rect 67634 543028 67640 543040
rect 60792 543000 67640 543028
rect 60792 542988 60798 543000
rect 67634 542988 67640 543000
rect 67692 542988 67698 543040
rect 130746 542988 130752 543040
rect 130804 543028 130810 543040
rect 139394 543028 139400 543040
rect 130804 543000 139400 543028
rect 130804 542988 130810 543000
rect 139394 542988 139400 543000
rect 139452 542988 139458 543040
rect 34146 541628 34152 541680
rect 34204 541668 34210 541680
rect 65518 541668 65524 541680
rect 34204 541640 65524 541668
rect 34204 541628 34210 541640
rect 65518 541628 65524 541640
rect 65576 541668 65582 541680
rect 67634 541668 67640 541680
rect 65576 541640 67640 541668
rect 65576 541628 65582 541640
rect 67634 541628 67640 541640
rect 67692 541628 67698 541680
rect 108850 540948 108856 541000
rect 108908 540988 108914 541000
rect 110414 540988 110420 541000
rect 108908 540960 110420 540988
rect 108908 540948 108914 540960
rect 110414 540948 110420 540960
rect 110472 540948 110478 541000
rect 62022 540880 62028 540932
rect 62080 540920 62086 540932
rect 63310 540920 63316 540932
rect 62080 540892 63316 540920
rect 62080 540880 62086 540892
rect 63310 540880 63316 540892
rect 63368 540920 63374 540932
rect 67634 540920 67640 540932
rect 63368 540892 67640 540920
rect 63368 540880 63374 540892
rect 67634 540880 67640 540892
rect 67692 540880 67698 540932
rect 108942 540880 108948 540932
rect 109000 540920 109006 540932
rect 127158 540920 127164 540932
rect 109000 540892 127164 540920
rect 109000 540880 109006 540892
rect 127158 540880 127164 540892
rect 127216 540920 127222 540932
rect 131298 540920 131304 540932
rect 127216 540892 131304 540920
rect 127216 540880 127222 540892
rect 131298 540880 131304 540892
rect 131356 540880 131362 540932
rect 110414 540812 110420 540864
rect 110472 540852 110478 540864
rect 111150 540852 111156 540864
rect 110472 540824 111156 540852
rect 110472 540812 110478 540824
rect 111150 540812 111156 540824
rect 111208 540852 111214 540864
rect 124306 540852 124312 540864
rect 111208 540824 124312 540852
rect 111208 540812 111214 540824
rect 124306 540812 124312 540824
rect 124364 540812 124370 540864
rect 37090 540336 37096 540388
rect 37148 540376 37154 540388
rect 38562 540376 38568 540388
rect 37148 540348 38568 540376
rect 37148 540336 37154 540348
rect 38562 540336 38568 540348
rect 38620 540336 38626 540388
rect 48038 540200 48044 540252
rect 48096 540240 48102 540252
rect 60090 540240 60096 540252
rect 48096 540212 60096 540240
rect 48096 540200 48102 540212
rect 60090 540200 60096 540212
rect 60148 540240 60154 540252
rect 60366 540240 60372 540252
rect 60148 540212 60372 540240
rect 60148 540200 60154 540212
rect 60366 540200 60372 540212
rect 60424 540200 60430 540252
rect 122926 540240 122932 540252
rect 113146 540212 122932 540240
rect 103698 539928 103704 539980
rect 103756 539968 103762 539980
rect 113146 539968 113174 540212
rect 122926 540200 122932 540212
rect 122984 540200 122990 540252
rect 103756 539940 113174 539968
rect 103756 539928 103762 539940
rect 105538 539860 105544 539912
rect 105596 539900 105602 539912
rect 105814 539900 105820 539912
rect 105596 539872 105820 539900
rect 105596 539860 105602 539872
rect 105814 539860 105820 539872
rect 105872 539860 105878 539912
rect 38470 539724 38476 539776
rect 38528 539764 38534 539776
rect 45278 539764 45284 539776
rect 38528 539736 45284 539764
rect 38528 539724 38534 539736
rect 45278 539724 45284 539736
rect 45336 539764 45342 539776
rect 70486 539764 70492 539776
rect 45336 539736 70492 539764
rect 45336 539724 45342 539736
rect 70486 539724 70492 539736
rect 70544 539724 70550 539776
rect 60090 539656 60096 539708
rect 60148 539696 60154 539708
rect 71958 539696 71964 539708
rect 60148 539668 71964 539696
rect 60148 539656 60154 539668
rect 71958 539656 71964 539668
rect 72016 539656 72022 539708
rect 38562 539588 38568 539640
rect 38620 539628 38626 539640
rect 71314 539628 71320 539640
rect 38620 539600 71320 539628
rect 38620 539588 38626 539600
rect 71314 539588 71320 539600
rect 71372 539588 71378 539640
rect 108022 539588 108028 539640
rect 108080 539628 108086 539640
rect 113174 539628 113180 539640
rect 108080 539600 113180 539628
rect 108080 539588 108086 539600
rect 113174 539588 113180 539600
rect 113232 539588 113238 539640
rect 132862 539628 132868 539640
rect 132466 539600 132868 539628
rect 40678 539520 40684 539572
rect 40736 539560 40742 539572
rect 114554 539560 114560 539572
rect 40736 539532 114560 539560
rect 40736 539520 40742 539532
rect 114554 539520 114560 539532
rect 114612 539560 114618 539572
rect 115198 539560 115204 539572
rect 114612 539532 115204 539560
rect 114612 539520 114618 539532
rect 115198 539520 115204 539532
rect 115256 539520 115262 539572
rect 42702 539452 42708 539504
rect 42760 539492 42766 539504
rect 45370 539492 45376 539504
rect 42760 539464 45376 539492
rect 42760 539452 42766 539464
rect 45370 539452 45376 539464
rect 45428 539492 45434 539504
rect 75178 539492 75184 539504
rect 45428 539464 75184 539492
rect 45428 539452 45434 539464
rect 75178 539452 75184 539464
rect 75236 539452 75242 539504
rect 97718 539452 97724 539504
rect 97776 539492 97782 539504
rect 131758 539492 131764 539504
rect 97776 539464 131764 539492
rect 97776 539452 97782 539464
rect 131758 539452 131764 539464
rect 131816 539492 131822 539504
rect 132466 539492 132494 539600
rect 132862 539588 132868 539600
rect 132920 539588 132926 539640
rect 131816 539464 132494 539492
rect 131816 539452 131822 539464
rect 52362 539384 52368 539436
rect 52420 539424 52426 539436
rect 77754 539424 77760 539436
rect 52420 539396 77760 539424
rect 52420 539384 52426 539396
rect 77754 539384 77760 539396
rect 77812 539384 77818 539436
rect 132678 539424 132684 539436
rect 103486 539396 132684 539424
rect 99650 539248 99656 539300
rect 99708 539288 99714 539300
rect 100570 539288 100576 539300
rect 99708 539260 100576 539288
rect 99708 539248 99714 539260
rect 100570 539248 100576 539260
rect 100628 539288 100634 539300
rect 103486 539288 103514 539396
rect 132678 539384 132684 539396
rect 132736 539384 132742 539436
rect 104158 539316 104164 539368
rect 104216 539356 104222 539368
rect 104710 539356 104716 539368
rect 104216 539328 104716 539356
rect 104216 539316 104222 539328
rect 104710 539316 104716 539328
rect 104768 539356 104774 539368
rect 120166 539356 120172 539368
rect 104768 539328 120172 539356
rect 104768 539316 104774 539328
rect 120166 539316 120172 539328
rect 120224 539316 120230 539368
rect 100628 539260 103514 539288
rect 100628 539248 100634 539260
rect 105630 538976 105636 539028
rect 105688 539016 105694 539028
rect 105814 539016 105820 539028
rect 105688 538988 105820 539016
rect 105688 538976 105694 538988
rect 105814 538976 105820 538988
rect 105872 538976 105878 539028
rect 52086 538908 52092 538960
rect 52144 538948 52150 538960
rect 73338 538948 73344 538960
rect 52144 538920 73344 538948
rect 52144 538908 52150 538920
rect 73338 538908 73344 538920
rect 73396 538908 73402 538960
rect 103238 538908 103244 538960
rect 103296 538948 103302 538960
rect 106366 538948 106372 538960
rect 103296 538920 106372 538948
rect 103296 538908 103302 538920
rect 106366 538908 106372 538920
rect 106424 538908 106430 538960
rect 3418 538840 3424 538892
rect 3476 538880 3482 538892
rect 93854 538880 93860 538892
rect 3476 538852 93860 538880
rect 3476 538840 3482 538852
rect 93854 538840 93860 538852
rect 93912 538840 93918 538892
rect 99282 538840 99288 538892
rect 99340 538880 99346 538892
rect 111242 538880 111248 538892
rect 99340 538852 111248 538880
rect 99340 538840 99346 538852
rect 111242 538840 111248 538852
rect 111300 538840 111306 538892
rect 119338 538228 119344 538280
rect 119396 538268 119402 538280
rect 125686 538268 125692 538280
rect 119396 538240 125692 538268
rect 119396 538228 119402 538240
rect 125686 538228 125692 538240
rect 125744 538228 125750 538280
rect 70118 538160 70124 538212
rect 70176 538200 70182 538212
rect 86126 538200 86132 538212
rect 70176 538172 86132 538200
rect 70176 538160 70182 538172
rect 86126 538160 86132 538172
rect 86184 538160 86190 538212
rect 93854 538160 93860 538212
rect 93912 538200 93918 538212
rect 98362 538200 98368 538212
rect 93912 538172 98368 538200
rect 93912 538160 93918 538172
rect 98362 538160 98368 538172
rect 98420 538160 98426 538212
rect 100294 538160 100300 538212
rect 100352 538200 100358 538212
rect 128354 538200 128360 538212
rect 100352 538172 128360 538200
rect 100352 538160 100358 538172
rect 128354 538160 128360 538172
rect 128412 538160 128418 538212
rect 50706 538092 50712 538144
rect 50764 538132 50770 538144
rect 80330 538132 80336 538144
rect 50764 538104 80336 538132
rect 50764 538092 50770 538104
rect 80330 538092 80336 538104
rect 80388 538092 80394 538144
rect 102226 538092 102232 538144
rect 102284 538132 102290 538144
rect 131114 538132 131120 538144
rect 102284 538104 131120 538132
rect 102284 538092 102290 538104
rect 131114 538092 131120 538104
rect 131172 538092 131178 538144
rect 54938 538024 54944 538076
rect 54996 538064 55002 538076
rect 83550 538064 83556 538076
rect 54996 538036 83556 538064
rect 54996 538024 55002 538036
rect 83550 538024 83556 538036
rect 83608 538024 83614 538076
rect 94498 538024 94504 538076
rect 94556 538064 94562 538076
rect 119338 538064 119344 538076
rect 94556 538036 119344 538064
rect 94556 538024 94562 538036
rect 119338 538024 119344 538036
rect 119396 538024 119402 538076
rect 52270 537956 52276 538008
rect 52328 537996 52334 538008
rect 78398 537996 78404 538008
rect 52328 537968 78404 537996
rect 52328 537956 52334 537968
rect 78398 537956 78404 537968
rect 78456 537956 78462 538008
rect 99006 537956 99012 538008
rect 99064 537996 99070 538008
rect 121454 537996 121460 538008
rect 99064 537968 121460 537996
rect 99064 537956 99070 537968
rect 121454 537956 121460 537968
rect 121512 537956 121518 538008
rect 56318 537888 56324 537940
rect 56376 537928 56382 537940
rect 73246 537928 73252 537940
rect 56376 537900 73252 537928
rect 56376 537888 56382 537900
rect 73246 537888 73252 537900
rect 73304 537888 73310 537940
rect 73338 537888 73344 537940
rect 73396 537928 73402 537940
rect 80974 537928 80980 537940
rect 73396 537900 80980 537928
rect 73396 537888 73402 537900
rect 80974 537888 80980 537900
rect 81032 537888 81038 537940
rect 103514 537888 103520 537940
rect 103572 537928 103578 537940
rect 122834 537928 122840 537940
rect 103572 537900 122840 537928
rect 103572 537888 103578 537900
rect 122834 537888 122840 537900
rect 122892 537888 122898 537940
rect 44082 537820 44088 537872
rect 44140 537860 44146 537872
rect 74534 537860 74540 537872
rect 44140 537832 74540 537860
rect 44140 537820 44146 537832
rect 74534 537820 74540 537832
rect 74592 537820 74598 537872
rect 93210 537820 93216 537872
rect 93268 537860 93274 537872
rect 93762 537860 93768 537872
rect 93268 537832 93768 537860
rect 93268 537820 93274 537832
rect 93762 537820 93768 537832
rect 93820 537860 93826 537872
rect 109770 537860 109776 537872
rect 93820 537832 109776 537860
rect 93820 537820 93826 537832
rect 109770 537820 109776 537832
rect 109828 537820 109834 537872
rect 43990 537548 43996 537600
rect 44048 537588 44054 537600
rect 52270 537588 52276 537600
rect 44048 537560 52276 537588
rect 44048 537548 44054 537560
rect 52270 537548 52276 537560
rect 52328 537548 52334 537600
rect 89346 537548 89352 537600
rect 89404 537588 89410 537600
rect 97902 537588 97908 537600
rect 89404 537560 97908 537588
rect 89404 537548 89410 537560
rect 97902 537548 97908 537560
rect 97960 537588 97966 537600
rect 103698 537588 103704 537600
rect 97960 537560 103704 537588
rect 97960 537548 97966 537560
rect 103698 537548 103704 537560
rect 103756 537548 103762 537600
rect 45370 537480 45376 537532
rect 45428 537520 45434 537532
rect 56318 537520 56324 537532
rect 45428 537492 56324 537520
rect 45428 537480 45434 537492
rect 56318 537480 56324 537492
rect 56376 537480 56382 537532
rect 87414 537480 87420 537532
rect 87472 537520 87478 537532
rect 99374 537520 99380 537532
rect 87472 537492 99380 537520
rect 87472 537480 87478 537492
rect 99374 537480 99380 537492
rect 99432 537480 99438 537532
rect 119430 537480 119436 537532
rect 119488 537520 119494 537532
rect 142430 537520 142436 537532
rect 119488 537492 142436 537520
rect 119488 537480 119494 537492
rect 142430 537480 142436 537492
rect 142488 537480 142494 537532
rect 46474 536868 46480 536920
rect 46532 536908 46538 536920
rect 50706 536908 50712 536920
rect 46532 536880 50712 536908
rect 46532 536868 46538 536880
rect 50706 536868 50712 536880
rect 50764 536868 50770 536920
rect 99466 536868 99472 536920
rect 99524 536908 99530 536920
rect 100294 536908 100300 536920
rect 99524 536880 100300 536908
rect 99524 536868 99530 536880
rect 100294 536868 100300 536880
rect 100352 536868 100358 536920
rect 121454 536868 121460 536920
rect 121512 536908 121518 536920
rect 124858 536908 124864 536920
rect 121512 536880 124864 536908
rect 121512 536868 121518 536880
rect 124858 536868 124864 536880
rect 124916 536868 124922 536920
rect 49602 536800 49608 536852
rect 49660 536840 49666 536852
rect 54938 536840 54944 536852
rect 49660 536812 54944 536840
rect 49660 536800 49666 536812
rect 54938 536800 54944 536812
rect 54996 536800 55002 536852
rect 73338 536800 73344 536852
rect 73396 536840 73402 536852
rect 73798 536840 73804 536852
rect 73396 536812 73804 536840
rect 73396 536800 73402 536812
rect 73798 536800 73804 536812
rect 73856 536800 73862 536852
rect 82814 536800 82820 536852
rect 82872 536840 82878 536852
rect 83458 536840 83464 536852
rect 82872 536812 83464 536840
rect 82872 536800 82878 536812
rect 83458 536800 83464 536812
rect 83516 536840 83522 536852
rect 85482 536840 85488 536852
rect 83516 536812 85488 536840
rect 83516 536800 83522 536812
rect 85482 536800 85488 536812
rect 85540 536800 85546 536852
rect 97074 536800 97080 536852
rect 97132 536840 97138 536852
rect 97132 536812 103514 536840
rect 97132 536800 97138 536812
rect 59170 536732 59176 536784
rect 59228 536772 59234 536784
rect 91002 536772 91008 536784
rect 59228 536744 91008 536772
rect 59228 536732 59234 536744
rect 91002 536732 91008 536744
rect 91060 536732 91066 536784
rect 103486 536772 103514 536812
rect 115842 536800 115848 536852
rect 115900 536840 115906 536852
rect 121730 536840 121736 536852
rect 115900 536812 121736 536840
rect 115900 536800 115906 536812
rect 121730 536800 121736 536812
rect 121788 536800 121794 536852
rect 122834 536800 122840 536852
rect 122892 536840 122898 536852
rect 123478 536840 123484 536852
rect 122892 536812 123484 536840
rect 122892 536800 122898 536812
rect 123478 536800 123484 536812
rect 123536 536800 123542 536852
rect 142430 536800 142436 536852
rect 142488 536840 142494 536852
rect 580166 536840 580172 536852
rect 142488 536812 580172 536840
rect 142488 536800 142494 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 112254 536772 112260 536784
rect 103486 536744 112260 536772
rect 112254 536732 112260 536744
rect 112312 536732 112318 536784
rect 50614 536664 50620 536716
rect 50672 536704 50678 536716
rect 54754 536704 54760 536716
rect 50672 536676 54760 536704
rect 50672 536664 50678 536676
rect 54754 536664 54760 536676
rect 54812 536704 54818 536716
rect 82906 536704 82912 536716
rect 54812 536676 82912 536704
rect 54812 536664 54818 536676
rect 82906 536664 82912 536676
rect 82964 536664 82970 536716
rect 88058 536664 88064 536716
rect 88116 536704 88122 536716
rect 115860 536704 115888 536800
rect 88116 536676 115888 536704
rect 88116 536664 88122 536676
rect 57698 536596 57704 536648
rect 57756 536636 57762 536648
rect 82814 536636 82820 536648
rect 57756 536608 82820 536636
rect 57756 536596 57762 536608
rect 82814 536596 82820 536608
rect 82872 536596 82878 536648
rect 93946 536596 93952 536648
rect 94004 536636 94010 536648
rect 120074 536636 120080 536648
rect 94004 536608 120080 536636
rect 94004 536596 94010 536608
rect 120074 536596 120080 536608
rect 120132 536596 120138 536648
rect 98362 536528 98368 536580
rect 98420 536568 98426 536580
rect 117314 536568 117320 536580
rect 98420 536540 117320 536568
rect 98420 536528 98426 536540
rect 117314 536528 117320 536540
rect 117372 536528 117378 536580
rect 95786 536460 95792 536512
rect 95844 536500 95850 536512
rect 124214 536500 124220 536512
rect 95844 536472 124220 536500
rect 95844 536460 95850 536472
rect 124214 536460 124220 536472
rect 124272 536460 124278 536512
rect 112254 536324 112260 536376
rect 112312 536364 112318 536376
rect 112898 536364 112904 536376
rect 112312 536336 112904 536364
rect 112312 536324 112318 536336
rect 112898 536324 112904 536336
rect 112956 536364 112962 536376
rect 113174 536364 113180 536376
rect 112956 536336 113180 536364
rect 112956 536324 112962 536336
rect 113174 536324 113180 536336
rect 113232 536324 113238 536376
rect 46842 536052 46848 536104
rect 46900 536092 46906 536104
rect 51718 536092 51724 536104
rect 46900 536064 51724 536092
rect 46900 536052 46906 536064
rect 51718 536052 51724 536064
rect 51776 536092 51782 536104
rect 73890 536092 73896 536104
rect 51776 536064 73896 536092
rect 51776 536052 51782 536064
rect 73890 536052 73896 536064
rect 73948 536052 73954 536104
rect 120074 536052 120080 536104
rect 120132 536092 120138 536104
rect 128446 536092 128452 536104
rect 120132 536064 128452 536092
rect 120132 536052 120138 536064
rect 128446 536052 128452 536064
rect 128504 536052 128510 536104
rect 117314 535440 117320 535492
rect 117372 535480 117378 535492
rect 119338 535480 119344 535492
rect 117372 535452 119344 535480
rect 117372 535440 117378 535452
rect 119338 535440 119344 535452
rect 119396 535440 119402 535492
rect 124214 535440 124220 535492
rect 124272 535480 124278 535492
rect 125778 535480 125784 535492
rect 124272 535452 125784 535480
rect 124272 535440 124278 535452
rect 125778 535440 125784 535452
rect 125836 535440 125842 535492
rect 39758 535372 39764 535424
rect 39816 535412 39822 535424
rect 72602 535412 72608 535424
rect 39816 535384 72608 535412
rect 39816 535372 39822 535384
rect 72602 535372 72608 535384
rect 72660 535372 72666 535424
rect 92566 535372 92572 535424
rect 92624 535412 92630 535424
rect 126974 535412 126980 535424
rect 92624 535384 126980 535412
rect 92624 535372 92630 535384
rect 126974 535372 126980 535384
rect 127032 535372 127038 535424
rect 130378 535372 130384 535424
rect 130436 535412 130442 535424
rect 131114 535412 131120 535424
rect 130436 535384 131120 535412
rect 130436 535372 130442 535384
rect 131114 535372 131120 535384
rect 131172 535372 131178 535424
rect 53742 535304 53748 535356
rect 53800 535344 53806 535356
rect 86770 535344 86776 535356
rect 53800 535316 86776 535344
rect 53800 535304 53806 535316
rect 86770 535304 86776 535316
rect 86828 535304 86834 535356
rect 100938 535304 100944 535356
rect 100996 535344 101002 535356
rect 102042 535344 102048 535356
rect 100996 535316 102048 535344
rect 100996 535304 101002 535316
rect 102042 535304 102048 535316
rect 102100 535344 102106 535356
rect 133874 535344 133880 535356
rect 102100 535316 133880 535344
rect 102100 535304 102106 535316
rect 133874 535304 133880 535316
rect 133932 535304 133938 535356
rect 48222 535236 48228 535288
rect 48280 535276 48286 535288
rect 79042 535276 79048 535288
rect 48280 535248 79048 535276
rect 48280 535236 48286 535248
rect 79042 535236 79048 535248
rect 79100 535236 79106 535288
rect 49326 535168 49332 535220
rect 49384 535208 49390 535220
rect 79686 535208 79692 535220
rect 49384 535180 79692 535208
rect 49384 535168 49390 535180
rect 79686 535168 79692 535180
rect 79744 535168 79750 535220
rect 89990 534760 89996 534812
rect 90048 534800 90054 534812
rect 114738 534800 114744 534812
rect 90048 534772 114744 534800
rect 90048 534760 90054 534772
rect 114738 534760 114744 534772
rect 114796 534800 114802 534812
rect 121546 534800 121552 534812
rect 114796 534772 121552 534800
rect 114796 534760 114802 534772
rect 121546 534760 121552 534772
rect 121604 534760 121610 534812
rect 96430 534692 96436 534744
rect 96488 534732 96494 534744
rect 127158 534732 127164 534744
rect 96488 534704 127164 534732
rect 96488 534692 96494 534704
rect 127158 534692 127164 534704
rect 127216 534732 127222 534744
rect 129734 534732 129740 534744
rect 127216 534704 129740 534732
rect 127216 534692 127222 534704
rect 129734 534692 129740 534704
rect 129792 534692 129798 534744
rect 46658 534080 46664 534132
rect 46716 534120 46722 534132
rect 48222 534120 48228 534132
rect 46716 534092 48228 534120
rect 46716 534080 46722 534092
rect 48222 534080 48228 534092
rect 48280 534080 48286 534132
rect 126974 534080 126980 534132
rect 127032 534120 127038 534132
rect 131114 534120 131120 534132
rect 127032 534092 131120 534120
rect 127032 534080 127038 534092
rect 131114 534080 131120 534092
rect 131172 534080 131178 534132
rect 50982 534012 50988 534064
rect 51040 534052 51046 534064
rect 55030 534052 55036 534064
rect 51040 534024 55036 534052
rect 51040 534012 51046 534024
rect 55030 534012 55036 534024
rect 55088 534052 55094 534064
rect 84838 534052 84844 534064
rect 55088 534024 84844 534052
rect 55088 534012 55094 534024
rect 84838 534012 84844 534024
rect 84896 534012 84902 534064
rect 102870 534012 102876 534064
rect 102928 534052 102934 534064
rect 136634 534052 136640 534064
rect 102928 534024 136640 534052
rect 102928 534012 102934 534024
rect 136634 534012 136640 534024
rect 136692 534012 136698 534064
rect 57882 533944 57888 533996
rect 57940 533984 57946 533996
rect 84194 533984 84200 533996
rect 57940 533956 84200 533984
rect 57940 533944 57946 533956
rect 84194 533944 84200 533956
rect 84252 533944 84258 533996
rect 89622 533468 89628 533520
rect 89680 533508 89686 533520
rect 118878 533508 118884 533520
rect 89680 533480 118884 533508
rect 89680 533468 89686 533480
rect 118878 533468 118884 533480
rect 118936 533468 118942 533520
rect 56226 533400 56232 533452
rect 56284 533440 56290 533452
rect 83550 533440 83556 533452
rect 56284 533412 83556 533440
rect 56284 533400 56290 533412
rect 83550 533400 83556 533412
rect 83608 533400 83614 533452
rect 95142 533400 95148 533452
rect 95200 533440 95206 533452
rect 127250 533440 127256 533452
rect 95200 533412 127256 533440
rect 95200 533400 95206 533412
rect 127250 533400 127256 533412
rect 127308 533400 127314 533452
rect 42518 533332 42524 533384
rect 42576 533372 42582 533384
rect 45278 533372 45284 533384
rect 42576 533344 45284 533372
rect 42576 533332 42582 533344
rect 45278 533332 45284 533344
rect 45336 533372 45342 533384
rect 76466 533372 76472 533384
rect 45336 533344 76472 533372
rect 45336 533332 45342 533344
rect 76466 533332 76472 533344
rect 76524 533332 76530 533384
rect 90634 533332 90640 533384
rect 90692 533372 90698 533384
rect 124214 533372 124220 533384
rect 90692 533344 124220 533372
rect 90692 533332 90698 533344
rect 124214 533332 124220 533344
rect 124272 533372 124278 533384
rect 125594 533372 125600 533384
rect 124272 533344 125600 533372
rect 124272 533332 124278 533344
rect 125594 533332 125600 533344
rect 125652 533332 125658 533384
rect 91002 530680 91008 530732
rect 91060 530680 91066 530732
rect 91922 530680 91928 530732
rect 91980 530720 91986 530732
rect 109034 530720 109040 530732
rect 91980 530692 109040 530720
rect 91980 530680 91986 530692
rect 109034 530680 109040 530692
rect 109092 530680 109098 530732
rect 57330 530612 57336 530664
rect 57388 530652 57394 530664
rect 77110 530652 77116 530664
rect 57388 530624 77116 530652
rect 57388 530612 57394 530624
rect 77110 530612 77116 530624
rect 77168 530612 77174 530664
rect 91020 530652 91048 530680
rect 120718 530652 120724 530664
rect 91020 530624 120724 530652
rect 120718 530612 120724 530624
rect 120776 530612 120782 530664
rect 45186 530544 45192 530596
rect 45244 530584 45250 530596
rect 79318 530584 79324 530596
rect 45244 530556 79324 530584
rect 45244 530544 45250 530556
rect 79318 530544 79324 530556
rect 79376 530544 79382 530596
rect 91002 530544 91008 530596
rect 91060 530584 91066 530596
rect 124490 530584 124496 530596
rect 91060 530556 124496 530584
rect 91060 530544 91066 530556
rect 124490 530544 124496 530556
rect 124548 530544 124554 530596
rect 46750 529864 46756 529916
rect 46808 529904 46814 529916
rect 57330 529904 57336 529916
rect 46808 529876 57336 529904
rect 46808 529864 46814 529876
rect 57330 529864 57336 529876
rect 57388 529864 57394 529916
rect 111058 528612 111064 528624
rect 106246 528584 111064 528612
rect 3142 528504 3148 528556
rect 3200 528544 3206 528556
rect 106246 528544 106274 528584
rect 111058 528572 111064 528584
rect 111116 528572 111122 528624
rect 3200 528516 106274 528544
rect 3200 528504 3206 528516
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 11698 514808 11704 514820
rect 3476 514780 11704 514808
rect 3476 514768 3482 514780
rect 11698 514768 11704 514780
rect 11756 514768 11762 514820
rect 431218 510620 431224 510672
rect 431276 510660 431282 510672
rect 580166 510660 580172 510672
rect 431276 510632 580172 510660
rect 431276 510620 431282 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 11698 498788 11704 498840
rect 11756 498828 11762 498840
rect 91094 498828 91100 498840
rect 11756 498800 91100 498828
rect 11756 498788 11762 498800
rect 91094 498788 91100 498800
rect 91152 498788 91158 498840
rect 86126 498176 86132 498228
rect 86184 498216 86190 498228
rect 121454 498216 121460 498228
rect 86184 498188 121460 498216
rect 86184 498176 86190 498188
rect 121454 498176 121460 498188
rect 121512 498176 121518 498228
rect 3142 497428 3148 497480
rect 3200 497468 3206 497480
rect 82906 497468 82912 497480
rect 3200 497440 82912 497468
rect 3200 497428 3206 497440
rect 82906 497428 82912 497440
rect 82964 497428 82970 497480
rect 96522 496068 96528 496120
rect 96580 496108 96586 496120
rect 128630 496108 128636 496120
rect 96580 496080 128636 496108
rect 96580 496068 96586 496080
rect 128630 496068 128636 496080
rect 128688 496108 128694 496120
rect 132494 496108 132500 496120
rect 128688 496080 132500 496108
rect 128688 496068 128694 496080
rect 132494 496068 132500 496080
rect 132552 496068 132558 496120
rect 82814 495524 82820 495576
rect 82872 495564 82878 495576
rect 83550 495564 83556 495576
rect 82872 495536 83556 495564
rect 82872 495524 82878 495536
rect 83550 495524 83556 495536
rect 83608 495564 83614 495576
rect 114554 495564 114560 495576
rect 83608 495536 114560 495564
rect 83608 495524 83614 495536
rect 114554 495524 114560 495536
rect 114612 495524 114618 495576
rect 124306 495496 124312 495508
rect 89732 495468 124312 495496
rect 85482 495388 85488 495440
rect 85540 495428 85546 495440
rect 89732 495428 89760 495468
rect 124306 495456 124312 495468
rect 124364 495496 124370 495508
rect 128354 495496 128360 495508
rect 124364 495468 128360 495496
rect 124364 495456 124370 495468
rect 128354 495456 128360 495468
rect 128412 495456 128418 495508
rect 85540 495400 89760 495428
rect 85540 495388 85546 495400
rect 90634 494776 90640 494828
rect 90692 494816 90698 494828
rect 114646 494816 114652 494828
rect 90692 494788 114652 494816
rect 90692 494776 90698 494788
rect 114646 494776 114652 494788
rect 114704 494816 114710 494828
rect 124306 494816 124312 494828
rect 114704 494788 124312 494816
rect 114704 494776 114710 494788
rect 124306 494776 124312 494788
rect 124364 494776 124370 494828
rect 56318 494708 56324 494760
rect 56376 494748 56382 494760
rect 73798 494748 73804 494760
rect 56376 494720 73804 494748
rect 56376 494708 56382 494720
rect 73798 494708 73804 494720
rect 73856 494708 73862 494760
rect 95142 494708 95148 494760
rect 95200 494748 95206 494760
rect 130102 494748 130108 494760
rect 95200 494720 130108 494748
rect 95200 494708 95206 494720
rect 130102 494708 130108 494720
rect 130160 494748 130166 494760
rect 134058 494748 134064 494760
rect 130160 494720 134064 494748
rect 130160 494708 130166 494720
rect 134058 494708 134064 494720
rect 134116 494708 134122 494760
rect 89990 494232 89996 494284
rect 90048 494272 90054 494284
rect 96522 494272 96528 494284
rect 90048 494244 96528 494272
rect 90048 494232 90054 494244
rect 96522 494232 96528 494244
rect 96580 494232 96586 494284
rect 92474 494028 92480 494080
rect 92532 494068 92538 494080
rect 93670 494068 93676 494080
rect 92532 494040 93676 494068
rect 92532 494028 92538 494040
rect 93670 494028 93676 494040
rect 93728 494068 93734 494080
rect 111794 494068 111800 494080
rect 93728 494040 111800 494068
rect 93728 494028 93734 494040
rect 111794 494028 111800 494040
rect 111852 494028 111858 494080
rect 82906 493960 82912 494012
rect 82964 494000 82970 494012
rect 83550 494000 83556 494012
rect 82964 493972 83556 494000
rect 82964 493960 82970 493972
rect 83550 493960 83556 493972
rect 83608 494000 83614 494012
rect 120074 494000 120080 494012
rect 83608 493972 120080 494000
rect 83608 493960 83614 493972
rect 120074 493960 120080 493972
rect 120132 493960 120138 494012
rect 110414 493892 110420 493944
rect 110472 493932 110478 493944
rect 111702 493932 111708 493944
rect 110472 493904 111708 493932
rect 110472 493892 110478 493904
rect 111702 493892 111708 493904
rect 111760 493932 111766 493944
rect 113910 493932 113916 493944
rect 111760 493904 113916 493932
rect 111760 493892 111766 493904
rect 113910 493892 113916 493904
rect 113968 493892 113974 493944
rect 88702 493824 88708 493876
rect 88760 493864 88766 493876
rect 89622 493864 89628 493876
rect 88760 493836 89628 493864
rect 88760 493824 88766 493836
rect 89622 493824 89628 493836
rect 89680 493824 89686 493876
rect 80974 493348 80980 493400
rect 81032 493388 81038 493400
rect 110414 493388 110420 493400
rect 81032 493360 110420 493388
rect 81032 493348 81038 493360
rect 110414 493348 110420 493360
rect 110472 493348 110478 493400
rect 120074 493348 120080 493400
rect 120132 493388 120138 493400
rect 129918 493388 129924 493400
rect 120132 493360 129924 493388
rect 120132 493348 120138 493360
rect 129918 493348 129924 493360
rect 129976 493348 129982 493400
rect 82906 493280 82912 493332
rect 82964 493320 82970 493332
rect 123110 493320 123116 493332
rect 82964 493292 123116 493320
rect 82964 493280 82970 493292
rect 123110 493280 123116 493292
rect 123168 493320 123174 493332
rect 127342 493320 127348 493332
rect 123168 493292 127348 493320
rect 123168 493280 123174 493292
rect 127342 493280 127348 493292
rect 127400 493280 127406 493332
rect 114646 492844 114652 492856
rect 84166 492816 114652 492844
rect 54846 492736 54852 492788
rect 54904 492776 54910 492788
rect 55122 492776 55128 492788
rect 54904 492748 55128 492776
rect 54904 492736 54910 492748
rect 55122 492736 55128 492748
rect 55180 492776 55186 492788
rect 81894 492776 81900 492788
rect 55180 492748 81900 492776
rect 55180 492736 55186 492748
rect 81894 492736 81900 492748
rect 81952 492736 81958 492788
rect 79318 492708 79324 492720
rect 78324 492680 79324 492708
rect 47946 492600 47952 492652
rect 48004 492640 48010 492652
rect 48222 492640 48228 492652
rect 48004 492612 48228 492640
rect 48004 492600 48010 492612
rect 48222 492600 48228 492612
rect 48280 492600 48286 492652
rect 53466 492600 53472 492652
rect 53524 492640 53530 492652
rect 53650 492640 53656 492652
rect 53524 492612 53656 492640
rect 53524 492600 53530 492612
rect 53650 492600 53656 492612
rect 53708 492600 53714 492652
rect 58710 492600 58716 492652
rect 58768 492640 58774 492652
rect 59170 492640 59176 492652
rect 58768 492612 59176 492640
rect 58768 492600 58774 492612
rect 59170 492600 59176 492612
rect 59228 492600 59234 492652
rect 77754 492600 77760 492652
rect 77812 492640 77818 492652
rect 78324 492640 78352 492680
rect 79318 492668 79324 492680
rect 79376 492708 79382 492720
rect 84166 492708 84194 492816
rect 114646 492804 114652 492816
rect 114704 492804 114710 492856
rect 88702 492736 88708 492788
rect 88760 492776 88766 492788
rect 110414 492776 110420 492788
rect 88760 492748 110420 492776
rect 88760 492736 88766 492748
rect 110414 492736 110420 492748
rect 110472 492736 110478 492788
rect 79376 492680 84194 492708
rect 79376 492668 79382 492680
rect 114462 492668 114468 492720
rect 114520 492708 114526 492720
rect 129826 492708 129832 492720
rect 114520 492680 129832 492708
rect 114520 492668 114526 492680
rect 129826 492668 129832 492680
rect 129884 492668 129890 492720
rect 77812 492612 78352 492640
rect 77812 492600 77818 492612
rect 78398 492600 78404 492652
rect 78456 492640 78462 492652
rect 82814 492640 82820 492652
rect 78456 492612 82820 492640
rect 78456 492600 78462 492612
rect 82814 492600 82820 492612
rect 82872 492600 82878 492652
rect 97810 492600 97816 492652
rect 97868 492640 97874 492652
rect 98178 492640 98184 492652
rect 97868 492612 98184 492640
rect 97868 492600 97874 492612
rect 98178 492600 98184 492612
rect 98236 492600 98242 492652
rect 91094 492192 91100 492244
rect 91152 492232 91158 492244
rect 131206 492232 131212 492244
rect 91152 492204 131212 492232
rect 91152 492192 91158 492204
rect 131206 492192 131212 492204
rect 131264 492192 131270 492244
rect 47854 492056 47860 492108
rect 47912 492096 47918 492108
rect 49418 492096 49424 492108
rect 47912 492068 49424 492096
rect 47912 492056 47918 492068
rect 49418 492056 49424 492068
rect 49476 492096 49482 492108
rect 49476 492068 55214 492096
rect 49476 492056 49482 492068
rect 55186 492028 55214 492068
rect 81618 492056 81624 492108
rect 81676 492096 81682 492108
rect 92474 492096 92480 492108
rect 81676 492068 92480 492096
rect 81676 492056 81682 492068
rect 92474 492056 92480 492068
rect 92532 492056 92538 492108
rect 99650 492056 99656 492108
rect 99708 492096 99714 492108
rect 112990 492096 112996 492108
rect 99708 492068 112996 492096
rect 99708 492056 99714 492068
rect 112990 492056 112996 492068
rect 113048 492096 113054 492108
rect 120166 492096 120172 492108
rect 113048 492068 120172 492096
rect 113048 492056 113054 492068
rect 120166 492056 120172 492068
rect 120224 492056 120230 492108
rect 70394 492028 70400 492040
rect 55186 492000 70400 492028
rect 70394 491988 70400 492000
rect 70452 491988 70458 492040
rect 88058 491988 88064 492040
rect 88116 492028 88122 492040
rect 99190 492028 99196 492040
rect 88116 492000 99196 492028
rect 88116 491988 88122 492000
rect 99190 491988 99196 492000
rect 99248 492028 99254 492040
rect 115934 492028 115940 492040
rect 99248 492000 115940 492028
rect 99248 491988 99254 492000
rect 115934 491988 115940 492000
rect 115992 491988 115998 492040
rect 41230 491920 41236 491972
rect 41288 491960 41294 491972
rect 43806 491960 43812 491972
rect 41288 491932 43812 491960
rect 41288 491920 41294 491932
rect 43806 491920 43812 491932
rect 43864 491960 43870 491972
rect 71774 491960 71780 491972
rect 43864 491932 71780 491960
rect 43864 491920 43870 491932
rect 71774 491920 71780 491932
rect 71832 491920 71838 491972
rect 92566 491580 92572 491632
rect 92624 491620 92630 491632
rect 99282 491620 99288 491632
rect 92624 491592 99288 491620
rect 92624 491580 92630 491592
rect 99282 491580 99288 491592
rect 99340 491580 99346 491632
rect 59170 491512 59176 491564
rect 59228 491552 59234 491564
rect 76742 491552 76748 491564
rect 59228 491524 76748 491552
rect 59228 491512 59234 491524
rect 76742 491512 76748 491524
rect 76800 491512 76806 491564
rect 93210 491512 93216 491564
rect 93268 491552 93274 491564
rect 100662 491552 100668 491564
rect 93268 491524 100668 491552
rect 93268 491512 93274 491524
rect 100662 491512 100668 491524
rect 100720 491512 100726 491564
rect 48222 491444 48228 491496
rect 48280 491484 48286 491496
rect 70026 491484 70032 491496
rect 48280 491456 70032 491484
rect 48280 491444 48286 491456
rect 70026 491444 70032 491456
rect 70084 491444 70090 491496
rect 91922 491444 91928 491496
rect 91980 491484 91986 491496
rect 95050 491484 95056 491496
rect 91980 491456 95056 491484
rect 91980 491444 91986 491456
rect 95050 491444 95056 491456
rect 95108 491444 95114 491496
rect 99190 491444 99196 491496
rect 99248 491484 99254 491496
rect 109770 491484 109776 491496
rect 99248 491456 109776 491484
rect 99248 491444 99254 491456
rect 109770 491444 109776 491456
rect 109828 491444 109834 491496
rect 52270 491376 52276 491428
rect 52328 491416 52334 491428
rect 74534 491416 74540 491428
rect 52328 491388 74540 491416
rect 52328 491376 52334 491388
rect 74534 491376 74540 491388
rect 74592 491416 74598 491428
rect 75454 491416 75460 491428
rect 74592 491388 75460 491416
rect 74592 491376 74598 491388
rect 75454 491376 75460 491388
rect 75512 491376 75518 491428
rect 97718 491376 97724 491428
rect 97776 491416 97782 491428
rect 97776 491388 98316 491416
rect 97776 491376 97782 491388
rect 53650 491308 53656 491360
rect 53708 491348 53714 491360
rect 80054 491348 80060 491360
rect 53708 491320 80060 491348
rect 53708 491308 53714 491320
rect 80054 491308 80060 491320
rect 80112 491308 80118 491360
rect 86770 491308 86776 491360
rect 86828 491348 86834 491360
rect 91002 491348 91008 491360
rect 86828 491320 91008 491348
rect 86828 491308 86834 491320
rect 91002 491308 91008 491320
rect 91060 491348 91066 491360
rect 91738 491348 91744 491360
rect 91060 491320 91744 491348
rect 91060 491308 91066 491320
rect 91738 491308 91744 491320
rect 91796 491308 91802 491360
rect 96430 491308 96436 491360
rect 96488 491348 96494 491360
rect 98178 491348 98184 491360
rect 96488 491320 98184 491348
rect 96488 491308 96494 491320
rect 98178 491308 98184 491320
rect 98236 491308 98242 491360
rect 98288 491348 98316 491388
rect 98362 491376 98368 491428
rect 98420 491416 98426 491428
rect 109862 491416 109868 491428
rect 98420 491388 109868 491416
rect 98420 491376 98426 491388
rect 109862 491376 109868 491388
rect 109920 491376 109926 491428
rect 110506 491348 110512 491360
rect 98288 491320 110512 491348
rect 110506 491308 110512 491320
rect 110564 491308 110570 491360
rect 97902 491240 97908 491292
rect 97960 491280 97966 491292
rect 102686 491280 102692 491292
rect 97960 491252 102692 491280
rect 97960 491240 97966 491252
rect 102686 491240 102692 491252
rect 102744 491240 102750 491292
rect 127066 491280 127072 491292
rect 109006 491252 127072 491280
rect 100662 491172 100668 491224
rect 100720 491212 100726 491224
rect 109006 491212 109034 491252
rect 127066 491240 127072 491252
rect 127124 491240 127130 491292
rect 100720 491184 109034 491212
rect 100720 491172 100726 491184
rect 109126 491172 109132 491224
rect 109184 491212 109190 491224
rect 109678 491212 109684 491224
rect 109184 491184 109684 491212
rect 109184 491172 109190 491184
rect 109678 491172 109684 491184
rect 109736 491212 109742 491224
rect 112530 491212 112536 491224
rect 109736 491184 112536 491212
rect 109736 491172 109742 491184
rect 112530 491172 112536 491184
rect 112588 491172 112594 491224
rect 91738 490628 91744 490680
rect 91796 490668 91802 490680
rect 101398 490668 101404 490680
rect 91796 490640 101404 490668
rect 91796 490628 91802 490640
rect 101398 490628 101404 490640
rect 101456 490628 101462 490680
rect 39942 490560 39948 490612
rect 40000 490600 40006 490612
rect 46566 490600 46572 490612
rect 40000 490572 46572 490600
rect 40000 490560 40006 490572
rect 46566 490560 46572 490572
rect 46624 490600 46630 490612
rect 72234 490600 72240 490612
rect 46624 490572 72240 490600
rect 46624 490560 46630 490572
rect 72234 490560 72240 490572
rect 72292 490560 72298 490612
rect 93762 490560 93768 490612
rect 93820 490600 93826 490612
rect 103514 490600 103520 490612
rect 93820 490572 103520 490600
rect 93820 490560 93826 490572
rect 103514 490560 103520 490572
rect 103572 490560 103578 490612
rect 48958 489948 48964 490000
rect 49016 489988 49022 490000
rect 74350 489988 74356 490000
rect 49016 489960 74356 489988
rect 49016 489948 49022 489960
rect 74350 489948 74356 489960
rect 74408 489948 74414 490000
rect 41046 489880 41052 489932
rect 41104 489920 41110 489932
rect 73062 489920 73068 489932
rect 41104 489892 73068 489920
rect 41104 489880 41110 489892
rect 73062 489880 73068 489892
rect 73120 489880 73126 489932
rect 98178 489812 98184 489864
rect 98236 489852 98242 489864
rect 99190 489852 99196 489864
rect 98236 489824 99196 489852
rect 98236 489812 98242 489824
rect 99190 489812 99196 489824
rect 99248 489812 99254 489864
rect 99282 489200 99288 489252
rect 99340 489240 99346 489252
rect 107286 489240 107292 489252
rect 99340 489212 107292 489240
rect 99340 489200 99346 489212
rect 107286 489200 107292 489212
rect 107344 489240 107350 489252
rect 112622 489240 112628 489252
rect 107344 489212 112628 489240
rect 107344 489200 107350 489212
rect 112622 489200 112628 489212
rect 112680 489200 112686 489252
rect 99190 489132 99196 489184
rect 99248 489172 99254 489184
rect 112438 489172 112444 489184
rect 99248 489144 112444 489172
rect 99248 489132 99254 489144
rect 112438 489132 112444 489144
rect 112496 489132 112502 489184
rect 67726 488560 67732 488572
rect 42812 488532 67732 488560
rect 42812 488504 42840 488532
rect 67726 488520 67732 488532
rect 67784 488520 67790 488572
rect 103422 488520 103428 488572
rect 103480 488560 103486 488572
rect 117222 488560 117228 488572
rect 103480 488532 117228 488560
rect 103480 488520 103486 488532
rect 117222 488520 117228 488532
rect 117280 488520 117286 488572
rect 123570 488560 123576 488572
rect 122806 488532 123576 488560
rect 39666 488452 39672 488504
rect 39724 488492 39730 488504
rect 42794 488492 42800 488504
rect 39724 488464 42800 488492
rect 39724 488452 39730 488464
rect 42794 488452 42800 488464
rect 42852 488452 42858 488504
rect 52178 488452 52184 488504
rect 52236 488492 52242 488504
rect 67634 488492 67640 488504
rect 52236 488464 67640 488492
rect 52236 488452 52242 488464
rect 67634 488452 67640 488464
rect 67692 488452 67698 488504
rect 103330 488452 103336 488504
rect 103388 488492 103394 488504
rect 122806 488492 122834 488532
rect 123570 488520 123576 488532
rect 123628 488560 123634 488572
rect 126974 488560 126980 488572
rect 123628 488532 126980 488560
rect 123628 488520 123634 488532
rect 126974 488520 126980 488532
rect 127032 488520 127038 488572
rect 103388 488464 122834 488492
rect 103388 488452 103394 488464
rect 52362 487772 52368 487824
rect 52420 487812 52426 487824
rect 67634 487812 67640 487824
rect 52420 487784 67640 487812
rect 52420 487772 52426 487784
rect 67634 487772 67640 487784
rect 67692 487772 67698 487824
rect 103422 487228 103428 487280
rect 103480 487268 103486 487280
rect 124122 487268 124128 487280
rect 103480 487240 124128 487268
rect 103480 487228 103486 487240
rect 124122 487228 124128 487240
rect 124180 487228 124186 487280
rect 104894 487160 104900 487212
rect 104952 487200 104958 487212
rect 105722 487200 105728 487212
rect 104952 487172 105728 487200
rect 104952 487160 104958 487172
rect 105722 487160 105728 487172
rect 105780 487200 105786 487212
rect 147766 487200 147772 487212
rect 105780 487172 147772 487200
rect 105780 487160 105786 487172
rect 147766 487160 147772 487172
rect 147824 487160 147830 487212
rect 102778 487092 102784 487144
rect 102836 487132 102842 487144
rect 140774 487132 140780 487144
rect 102836 487104 140780 487132
rect 102836 487092 102842 487104
rect 140774 487092 140780 487104
rect 140832 487092 140838 487144
rect 103330 487024 103336 487076
rect 103388 487064 103394 487076
rect 104894 487064 104900 487076
rect 103388 487036 104900 487064
rect 103388 487024 103394 487036
rect 104894 487024 104900 487036
rect 104952 487024 104958 487076
rect 124122 487024 124128 487076
rect 124180 487064 124186 487076
rect 125870 487064 125876 487076
rect 124180 487036 125876 487064
rect 124180 487024 124186 487036
rect 125870 487024 125876 487036
rect 125928 487024 125934 487076
rect 140774 486412 140780 486464
rect 140832 486452 140838 486464
rect 152090 486452 152096 486464
rect 140832 486424 152096 486452
rect 140832 486412 140838 486424
rect 152090 486412 152096 486424
rect 152148 486412 152154 486464
rect 53834 485868 53840 485920
rect 53892 485908 53898 485920
rect 67726 485908 67732 485920
rect 53892 485880 67732 485908
rect 53892 485868 53898 485880
rect 67726 485868 67732 485880
rect 67784 485868 67790 485920
rect 36630 485840 36636 485852
rect 35866 485812 36636 485840
rect 34330 485732 34336 485784
rect 34388 485772 34394 485784
rect 35866 485772 35894 485812
rect 36630 485800 36636 485812
rect 36688 485840 36694 485852
rect 67634 485840 67640 485852
rect 36688 485812 67640 485840
rect 36688 485800 36694 485812
rect 67634 485800 67640 485812
rect 67692 485800 67698 485852
rect 34388 485744 35894 485772
rect 34388 485732 34394 485744
rect 41322 485732 41328 485784
rect 41380 485772 41386 485784
rect 53834 485772 53840 485784
rect 41380 485744 53840 485772
rect 41380 485732 41386 485744
rect 53834 485732 53840 485744
rect 53892 485732 53898 485784
rect 102134 485120 102140 485172
rect 102192 485160 102198 485172
rect 114462 485160 114468 485172
rect 102192 485132 114468 485160
rect 102192 485120 102198 485132
rect 114462 485120 114468 485132
rect 114520 485120 114526 485172
rect 53558 485052 53564 485104
rect 53616 485092 53622 485104
rect 67634 485092 67640 485104
rect 53616 485064 67640 485092
rect 53616 485052 53622 485064
rect 67634 485052 67640 485064
rect 67692 485052 67698 485104
rect 102410 485052 102416 485104
rect 102468 485092 102474 485104
rect 117222 485092 117228 485104
rect 102468 485064 117228 485092
rect 102468 485052 102474 485064
rect 117222 485052 117228 485064
rect 117280 485052 117286 485104
rect 64690 484372 64696 484424
rect 64748 484412 64754 484424
rect 68462 484412 68468 484424
rect 64748 484384 68468 484412
rect 64748 484372 64754 484384
rect 68462 484372 68468 484384
rect 68520 484372 68526 484424
rect 117222 484372 117228 484424
rect 117280 484412 117286 484424
rect 125594 484412 125600 484424
rect 117280 484384 125600 484412
rect 117280 484372 117286 484384
rect 125594 484372 125600 484384
rect 125652 484372 125658 484424
rect 286318 484372 286324 484424
rect 286376 484412 286382 484424
rect 580166 484412 580172 484424
rect 286376 484384 580172 484412
rect 286376 484372 286382 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 35526 483624 35532 483676
rect 35584 483664 35590 483676
rect 35710 483664 35716 483676
rect 35584 483636 35716 483664
rect 35584 483624 35590 483636
rect 35710 483624 35716 483636
rect 35768 483664 35774 483676
rect 67634 483664 67640 483676
rect 35768 483636 67640 483664
rect 35768 483624 35774 483636
rect 67634 483624 67640 483636
rect 67692 483624 67698 483676
rect 36998 482944 37004 482996
rect 37056 482984 37062 482996
rect 68002 482984 68008 482996
rect 37056 482956 68008 482984
rect 37056 482944 37062 482956
rect 68002 482944 68008 482956
rect 68060 482944 68066 482996
rect 102134 482740 102140 482792
rect 102192 482780 102198 482792
rect 105538 482780 105544 482792
rect 102192 482752 105544 482780
rect 102192 482740 102198 482752
rect 105538 482740 105544 482752
rect 105596 482780 105602 482792
rect 110598 482780 110604 482792
rect 105596 482752 110604 482780
rect 105596 482740 105602 482752
rect 110598 482740 110604 482752
rect 110656 482740 110662 482792
rect 115842 481720 115848 481772
rect 115900 481760 115906 481772
rect 143718 481760 143724 481772
rect 115900 481732 143724 481760
rect 115900 481720 115906 481732
rect 143718 481720 143724 481732
rect 143776 481720 143782 481772
rect 40954 481652 40960 481704
rect 41012 481692 41018 481704
rect 68922 481692 68928 481704
rect 41012 481664 68928 481692
rect 41012 481652 41018 481664
rect 68922 481652 68928 481664
rect 68980 481652 68986 481704
rect 102686 481652 102692 481704
rect 102744 481692 102750 481704
rect 104894 481692 104900 481704
rect 102744 481664 104900 481692
rect 102744 481652 102750 481664
rect 104894 481652 104900 481664
rect 104952 481652 104958 481704
rect 107562 481652 107568 481704
rect 107620 481692 107626 481704
rect 143534 481692 143540 481704
rect 107620 481664 143540 481692
rect 107620 481652 107626 481664
rect 143534 481652 143540 481664
rect 143592 481652 143598 481704
rect 102134 481584 102140 481636
rect 102192 481624 102198 481636
rect 115198 481624 115204 481636
rect 102192 481596 115204 481624
rect 102192 481584 102198 481596
rect 115198 481584 115204 481596
rect 115256 481624 115262 481636
rect 115842 481624 115848 481636
rect 115256 481596 115848 481624
rect 115256 481584 115262 481596
rect 115842 481584 115848 481596
rect 115900 481584 115906 481636
rect 102226 481516 102232 481568
rect 102284 481556 102290 481568
rect 107378 481556 107384 481568
rect 102284 481528 107384 481556
rect 102284 481516 102290 481528
rect 107378 481516 107384 481528
rect 107436 481556 107442 481568
rect 107562 481556 107568 481568
rect 107436 481528 107568 481556
rect 107436 481516 107442 481528
rect 107562 481516 107568 481528
rect 107620 481516 107626 481568
rect 66254 480836 66260 480888
rect 66312 480876 66318 480888
rect 67634 480876 67640 480888
rect 66312 480848 67640 480876
rect 66312 480836 66318 480848
rect 67634 480836 67640 480848
rect 67692 480836 67698 480888
rect 61838 480156 61844 480208
rect 61896 480196 61902 480208
rect 67542 480196 67548 480208
rect 61896 480168 67548 480196
rect 61896 480156 61902 480168
rect 67542 480156 67548 480168
rect 67600 480156 67606 480208
rect 102134 480156 102140 480208
rect 102192 480196 102198 480208
rect 134150 480196 134156 480208
rect 102192 480168 134156 480196
rect 102192 480156 102198 480168
rect 134150 480156 134156 480168
rect 134208 480156 134214 480208
rect 35618 479476 35624 479528
rect 35676 479516 35682 479528
rect 39666 479516 39672 479528
rect 35676 479488 39672 479516
rect 35676 479476 35682 479488
rect 39666 479476 39672 479488
rect 39724 479516 39730 479528
rect 66254 479516 66260 479528
rect 39724 479488 66260 479516
rect 39724 479476 39730 479488
rect 66254 479476 66260 479488
rect 66312 479476 66318 479528
rect 50890 478932 50896 478984
rect 50948 478972 50954 478984
rect 52178 478972 52184 478984
rect 50948 478944 52184 478972
rect 50948 478932 50954 478944
rect 52178 478932 52184 478944
rect 52236 478972 52242 478984
rect 52236 478944 55214 478972
rect 52236 478932 52242 478944
rect 55186 478904 55214 478944
rect 105538 478932 105544 478984
rect 105596 478972 105602 478984
rect 115290 478972 115296 478984
rect 105596 478944 115296 478972
rect 105596 478932 105602 478944
rect 115290 478932 115296 478944
rect 115348 478932 115354 478984
rect 67634 478904 67640 478916
rect 55186 478876 67640 478904
rect 67634 478864 67640 478876
rect 67692 478864 67698 478916
rect 107378 478864 107384 478916
rect 107436 478904 107442 478916
rect 111150 478904 111156 478916
rect 107436 478876 111156 478904
rect 107436 478864 107442 478876
rect 111150 478864 111156 478876
rect 111208 478864 111214 478916
rect 134150 478864 134156 478916
rect 134208 478904 134214 478916
rect 140866 478904 140872 478916
rect 134208 478876 140872 478904
rect 134208 478864 134214 478876
rect 140866 478864 140872 478876
rect 140924 478864 140930 478916
rect 118602 477572 118608 477624
rect 118660 477612 118666 477624
rect 120074 477612 120080 477624
rect 118660 477584 120080 477612
rect 118660 477572 118666 477584
rect 120074 477572 120080 477584
rect 120132 477572 120138 477624
rect 61746 477504 61752 477556
rect 61804 477544 61810 477556
rect 63034 477544 63040 477556
rect 61804 477516 63040 477544
rect 61804 477504 61810 477516
rect 63034 477504 63040 477516
rect 63092 477544 63098 477556
rect 67634 477544 67640 477556
rect 63092 477516 67640 477544
rect 63092 477504 63098 477516
rect 67634 477504 67640 477516
rect 67692 477504 67698 477556
rect 111886 477504 111892 477556
rect 111944 477544 111950 477556
rect 113082 477544 113088 477556
rect 111944 477516 113088 477544
rect 111944 477504 111950 477516
rect 113082 477504 113088 477516
rect 113140 477544 113146 477556
rect 118694 477544 118700 477556
rect 113140 477516 118700 477544
rect 113140 477504 113146 477516
rect 118694 477504 118700 477516
rect 118752 477504 118758 477556
rect 103422 477436 103428 477488
rect 103480 477476 103486 477488
rect 136910 477476 136916 477488
rect 103480 477448 136916 477476
rect 103480 477436 103486 477448
rect 136910 477436 136916 477448
rect 136968 477436 136974 477488
rect 102134 477368 102140 477420
rect 102192 477408 102198 477420
rect 118602 477408 118608 477420
rect 102192 477380 118608 477408
rect 102192 477368 102198 477380
rect 118602 477368 118608 477380
rect 118660 477368 118666 477420
rect 102226 477300 102232 477352
rect 102284 477340 102290 477352
rect 111886 477340 111892 477352
rect 102284 477312 111892 477340
rect 102284 477300 102290 477312
rect 111886 477300 111892 477312
rect 111944 477300 111950 477352
rect 38562 476076 38568 476128
rect 38620 476116 38626 476128
rect 67634 476116 67640 476128
rect 38620 476088 67640 476116
rect 38620 476076 38626 476088
rect 67634 476076 67640 476088
rect 67692 476076 67698 476128
rect 102318 476008 102324 476060
rect 102376 476048 102382 476060
rect 103330 476048 103336 476060
rect 102376 476020 103336 476048
rect 102376 476008 102382 476020
rect 103330 476008 103336 476020
rect 103388 476048 103394 476060
rect 139486 476048 139492 476060
rect 103388 476020 139492 476048
rect 103388 476008 103394 476020
rect 139486 476008 139492 476020
rect 139544 476008 139550 476060
rect 43898 475396 43904 475448
rect 43956 475436 43962 475448
rect 67634 475436 67640 475448
rect 43956 475408 67640 475436
rect 43956 475396 43962 475408
rect 67634 475396 67640 475408
rect 67692 475396 67698 475448
rect 32950 475328 32956 475380
rect 33008 475368 33014 475380
rect 67726 475368 67732 475380
rect 33008 475340 67732 475368
rect 33008 475328 33014 475340
rect 67726 475328 67732 475340
rect 67784 475328 67790 475380
rect 102134 475328 102140 475380
rect 102192 475368 102198 475380
rect 132586 475368 132592 475380
rect 102192 475340 132592 475368
rect 102192 475328 102198 475340
rect 132586 475328 132592 475340
rect 132644 475328 132650 475380
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 11698 474756 11704 474768
rect 3476 474728 11704 474756
rect 3476 474716 3482 474728
rect 11698 474716 11704 474728
rect 11756 474716 11762 474768
rect 102134 474716 102140 474768
rect 102192 474756 102198 474768
rect 121454 474756 121460 474768
rect 102192 474728 121460 474756
rect 102192 474716 102198 474728
rect 121454 474716 121460 474728
rect 121512 474716 121518 474768
rect 102226 474648 102232 474700
rect 102284 474688 102290 474700
rect 134518 474688 134524 474700
rect 102284 474660 134524 474688
rect 102284 474648 102290 474660
rect 134518 474648 134524 474660
rect 134576 474688 134582 474700
rect 135438 474688 135444 474700
rect 134576 474660 135444 474688
rect 134576 474648 134582 474660
rect 135438 474648 135444 474660
rect 135496 474648 135502 474700
rect 121454 474580 121460 474632
rect 121512 474620 121518 474632
rect 122742 474620 122748 474632
rect 121512 474592 122748 474620
rect 121512 474580 121518 474592
rect 122742 474580 122748 474592
rect 122800 474620 122806 474632
rect 128538 474620 128544 474632
rect 122800 474592 128544 474620
rect 122800 474580 122806 474592
rect 128538 474580 128544 474592
rect 128596 474580 128602 474632
rect 66070 473288 66076 473340
rect 66128 473328 66134 473340
rect 67634 473328 67640 473340
rect 66128 473300 67640 473328
rect 66128 473288 66134 473300
rect 67634 473288 67640 473300
rect 67692 473288 67698 473340
rect 34330 472608 34336 472660
rect 34388 472648 34394 472660
rect 66070 472648 66076 472660
rect 34388 472620 66076 472648
rect 34388 472608 34394 472620
rect 66070 472608 66076 472620
rect 66128 472608 66134 472660
rect 102134 472608 102140 472660
rect 102192 472648 102198 472660
rect 142246 472648 142252 472660
rect 102192 472620 142252 472648
rect 102192 472608 102198 472620
rect 142246 472608 142252 472620
rect 142304 472648 142310 472660
rect 142430 472648 142436 472660
rect 142304 472620 142436 472648
rect 142304 472608 142310 472620
rect 142430 472608 142436 472620
rect 142488 472608 142494 472660
rect 102134 472064 102140 472116
rect 102192 472104 102198 472116
rect 121454 472104 121460 472116
rect 102192 472076 121460 472104
rect 102192 472064 102198 472076
rect 121454 472064 121460 472076
rect 121512 472064 121518 472116
rect 113818 472036 113824 472048
rect 113146 472008 113824 472036
rect 102134 471928 102140 471980
rect 102192 471968 102198 471980
rect 113146 471968 113174 472008
rect 113818 471996 113824 472008
rect 113876 472036 113882 472048
rect 133874 472036 133880 472048
rect 113876 472008 133880 472036
rect 113876 471996 113882 472008
rect 133874 471996 133880 472008
rect 133932 471996 133938 472048
rect 102192 471940 113174 471968
rect 102192 471928 102198 471940
rect 121454 471928 121460 471980
rect 121512 471968 121518 471980
rect 138014 471968 138020 471980
rect 121512 471940 138020 471968
rect 121512 471928 121518 471940
rect 138014 471928 138020 471940
rect 138072 471928 138078 471980
rect 104066 471452 104072 471504
rect 104124 471492 104130 471504
rect 107746 471492 107752 471504
rect 104124 471464 107752 471492
rect 104124 471452 104130 471464
rect 107746 471452 107752 471464
rect 107804 471452 107810 471504
rect 138014 471316 138020 471368
rect 138072 471356 138078 471368
rect 148962 471356 148968 471368
rect 138072 471328 148968 471356
rect 138072 471316 138078 471328
rect 148962 471316 148968 471328
rect 149020 471316 149026 471368
rect 101950 471248 101956 471300
rect 102008 471288 102014 471300
rect 135898 471288 135904 471300
rect 102008 471260 135904 471288
rect 102008 471248 102014 471260
rect 135898 471248 135904 471260
rect 135956 471288 135962 471300
rect 149238 471288 149244 471300
rect 135956 471260 149244 471288
rect 135956 471248 135962 471260
rect 149238 471248 149244 471260
rect 149296 471248 149302 471300
rect 65886 471044 65892 471096
rect 65944 471084 65950 471096
rect 67082 471084 67088 471096
rect 65944 471056 67088 471084
rect 65944 471044 65950 471056
rect 67082 471044 67088 471056
rect 67140 471084 67146 471096
rect 67726 471084 67732 471096
rect 67140 471056 67732 471084
rect 67140 471044 67146 471056
rect 67726 471044 67732 471056
rect 67784 471044 67790 471096
rect 102134 470568 102140 470620
rect 102192 470608 102198 470620
rect 102192 470580 138888 470608
rect 102192 470568 102198 470580
rect 138860 470540 138888 470580
rect 148962 470568 148968 470620
rect 149020 470608 149026 470620
rect 579982 470608 579988 470620
rect 149020 470580 579988 470608
rect 149020 470568 149026 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 139302 470540 139308 470552
rect 138860 470512 139308 470540
rect 139302 470500 139308 470512
rect 139360 470540 139366 470552
rect 142154 470540 142160 470552
rect 139360 470512 142160 470540
rect 139360 470500 139366 470512
rect 142154 470500 142160 470512
rect 142212 470500 142218 470552
rect 66162 470432 66168 470484
rect 66220 470472 66226 470484
rect 66990 470472 66996 470484
rect 66220 470444 66996 470472
rect 66220 470432 66226 470444
rect 66990 470432 66996 470444
rect 67048 470472 67054 470484
rect 67726 470472 67732 470484
rect 67048 470444 67732 470472
rect 67048 470432 67054 470444
rect 67726 470432 67732 470444
rect 67784 470432 67790 470484
rect 63310 470160 63316 470212
rect 63368 470200 63374 470212
rect 67634 470200 67640 470212
rect 63368 470172 67640 470200
rect 63368 470160 63374 470172
rect 67634 470160 67640 470172
rect 67692 470160 67698 470212
rect 102134 469820 102140 469872
rect 102192 469860 102198 469872
rect 117498 469860 117504 469872
rect 102192 469832 117504 469860
rect 102192 469820 102198 469832
rect 117498 469820 117504 469832
rect 117556 469820 117562 469872
rect 117498 469276 117504 469328
rect 117556 469316 117562 469328
rect 117682 469316 117688 469328
rect 117556 469288 117688 469316
rect 117556 469276 117562 469288
rect 117682 469276 117688 469288
rect 117740 469276 117746 469328
rect 107470 469208 107476 469260
rect 107528 469248 107534 469260
rect 145098 469248 145104 469260
rect 107528 469220 145104 469248
rect 107528 469208 107534 469220
rect 145098 469208 145104 469220
rect 145156 469208 145162 469260
rect 102134 469140 102140 469192
rect 102192 469180 102198 469192
rect 107488 469180 107516 469208
rect 102192 469152 107516 469180
rect 102192 469140 102198 469152
rect 60458 468460 60464 468512
rect 60516 468500 60522 468512
rect 67634 468500 67640 468512
rect 60516 468472 67640 468500
rect 60516 468460 60522 468472
rect 67634 468460 67640 468472
rect 67692 468460 67698 468512
rect 64230 467916 64236 467968
rect 64288 467956 64294 467968
rect 67634 467956 67640 467968
rect 64288 467928 67640 467956
rect 64288 467916 64294 467928
rect 67634 467916 67640 467928
rect 67692 467916 67698 467968
rect 106182 467848 106188 467900
rect 106240 467888 106246 467900
rect 146478 467888 146484 467900
rect 106240 467860 146484 467888
rect 106240 467848 106246 467860
rect 146478 467848 146484 467860
rect 146536 467848 146542 467900
rect 61930 467780 61936 467832
rect 61988 467820 61994 467832
rect 67450 467820 67456 467832
rect 61988 467792 67456 467820
rect 61988 467780 61994 467792
rect 67450 467780 67456 467792
rect 67508 467780 67514 467832
rect 102134 467780 102140 467832
rect 102192 467820 102198 467832
rect 132770 467820 132776 467832
rect 102192 467792 132776 467820
rect 102192 467780 102198 467792
rect 132770 467780 132776 467792
rect 132828 467820 132834 467832
rect 137002 467820 137008 467832
rect 132828 467792 137008 467820
rect 132828 467780 132834 467792
rect 137002 467780 137008 467792
rect 137060 467780 137066 467832
rect 102226 467712 102232 467764
rect 102284 467752 102290 467764
rect 106182 467752 106188 467764
rect 102284 467724 106188 467752
rect 102284 467712 102290 467724
rect 106182 467712 106188 467724
rect 106240 467712 106246 467764
rect 113910 467100 113916 467152
rect 113968 467140 113974 467152
rect 128538 467140 128544 467152
rect 113968 467112 128544 467140
rect 113968 467100 113974 467112
rect 128538 467100 128544 467112
rect 128596 467100 128602 467152
rect 100570 466760 100576 466812
rect 100628 466800 100634 466812
rect 101490 466800 101496 466812
rect 100628 466772 101496 466800
rect 100628 466760 100634 466772
rect 101490 466760 101496 466772
rect 101548 466760 101554 466812
rect 62758 466352 62764 466404
rect 62816 466392 62822 466404
rect 63494 466392 63500 466404
rect 62816 466364 63500 466392
rect 62816 466352 62822 466364
rect 63494 466352 63500 466364
rect 63552 466392 63558 466404
rect 67634 466392 67640 466404
rect 63552 466364 67640 466392
rect 63552 466352 63558 466364
rect 67634 466352 67640 466364
rect 67692 466352 67698 466404
rect 100018 465740 100024 465792
rect 100076 465780 100082 465792
rect 114738 465780 114744 465792
rect 100076 465752 114744 465780
rect 100076 465740 100082 465752
rect 114738 465740 114744 465752
rect 114796 465740 114802 465792
rect 54938 465672 54944 465724
rect 54996 465712 55002 465724
rect 66898 465712 66904 465724
rect 54996 465684 66904 465712
rect 54996 465672 55002 465684
rect 66898 465672 66904 465684
rect 66956 465712 66962 465724
rect 67726 465712 67732 465724
rect 66956 465684 67732 465712
rect 66956 465672 66962 465684
rect 67726 465672 67732 465684
rect 67784 465672 67790 465724
rect 102318 465672 102324 465724
rect 102376 465712 102382 465724
rect 141050 465712 141056 465724
rect 102376 465684 141056 465712
rect 102376 465672 102382 465684
rect 141050 465672 141056 465684
rect 141108 465712 141114 465724
rect 151906 465712 151912 465724
rect 141108 465684 151912 465712
rect 141108 465672 141114 465684
rect 151906 465672 151912 465684
rect 151964 465672 151970 465724
rect 102226 465060 102232 465112
rect 102284 465100 102290 465112
rect 102284 465072 120028 465100
rect 102284 465060 102290 465072
rect 120000 465044 120028 465072
rect 102134 464992 102140 465044
rect 102192 465032 102198 465044
rect 107562 465032 107568 465044
rect 102192 465004 107568 465032
rect 102192 464992 102198 465004
rect 107562 464992 107568 465004
rect 107620 464992 107626 465044
rect 119982 464992 119988 465044
rect 120040 465032 120046 465044
rect 121638 465032 121644 465044
rect 120040 465004 121644 465032
rect 120040 464992 120046 465004
rect 121638 464992 121644 465004
rect 121696 464992 121702 465044
rect 60550 464380 60556 464432
rect 60608 464420 60614 464432
rect 67726 464420 67732 464432
rect 60608 464392 67732 464420
rect 60608 464380 60614 464392
rect 67726 464380 67732 464392
rect 67784 464380 67790 464432
rect 49510 464312 49516 464364
rect 49568 464352 49574 464364
rect 67634 464352 67640 464364
rect 49568 464324 67640 464352
rect 49568 464312 49574 464324
rect 67634 464312 67640 464324
rect 67692 464312 67698 464364
rect 107562 464312 107568 464364
rect 107620 464352 107626 464364
rect 143810 464352 143816 464364
rect 107620 464324 143816 464352
rect 107620 464312 107626 464324
rect 143810 464312 143816 464324
rect 143868 464312 143874 464364
rect 121454 463740 121460 463752
rect 117056 463712 121460 463740
rect 102134 463632 102140 463684
rect 102192 463672 102198 463684
rect 116578 463672 116584 463684
rect 102192 463644 116584 463672
rect 102192 463632 102198 463644
rect 116578 463632 116584 463644
rect 116636 463672 116642 463684
rect 117056 463672 117084 463712
rect 121454 463700 121460 463712
rect 121512 463700 121518 463752
rect 116636 463644 117084 463672
rect 116636 463632 116642 463644
rect 117222 463632 117228 463684
rect 117280 463672 117286 463684
rect 117498 463672 117504 463684
rect 117280 463644 117504 463672
rect 117280 463632 117286 463644
rect 117498 463632 117504 463644
rect 117556 463632 117562 463684
rect 106550 463360 106556 463412
rect 106608 463400 106614 463412
rect 108298 463400 108304 463412
rect 106608 463372 108304 463400
rect 106608 463360 106614 463372
rect 108298 463360 108304 463372
rect 108356 463360 108362 463412
rect 54478 462952 54484 463004
rect 54536 462992 54542 463004
rect 59078 462992 59084 463004
rect 54536 462964 59084 462992
rect 54536 462952 54542 462964
rect 59078 462952 59084 462964
rect 59136 462952 59142 463004
rect 106182 462952 106188 463004
rect 106240 462992 106246 463004
rect 136726 462992 136732 463004
rect 106240 462964 136732 462992
rect 106240 462952 106246 462964
rect 136726 462952 136732 462964
rect 136784 462992 136790 463004
rect 146386 462992 146392 463004
rect 136784 462964 146392 462992
rect 136784 462952 136790 462964
rect 146386 462952 146392 462964
rect 146444 462952 146450 463004
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 59078 462340 59084 462392
rect 59136 462380 59142 462392
rect 67634 462380 67640 462392
rect 59136 462352 67640 462380
rect 59136 462340 59142 462352
rect 67634 462340 67640 462352
rect 67692 462340 67698 462392
rect 102226 462272 102232 462324
rect 102284 462312 102290 462324
rect 133966 462312 133972 462324
rect 102284 462284 133972 462312
rect 102284 462272 102290 462284
rect 133966 462272 133972 462284
rect 134024 462312 134030 462324
rect 141050 462312 141056 462324
rect 134024 462284 141056 462312
rect 134024 462272 134030 462284
rect 141050 462272 141056 462284
rect 141108 462272 141114 462324
rect 102134 462204 102140 462256
rect 102192 462244 102198 462256
rect 106182 462244 106188 462256
rect 102192 462216 106188 462244
rect 102192 462204 102198 462216
rect 106182 462204 106188 462216
rect 106240 462204 106246 462256
rect 106550 460952 106556 460964
rect 106246 460924 106556 460952
rect 102134 460844 102140 460896
rect 102192 460884 102198 460896
rect 106246 460884 106274 460924
rect 106550 460912 106556 460924
rect 106608 460952 106614 460964
rect 147674 460952 147680 460964
rect 106608 460924 147680 460952
rect 106608 460912 106614 460924
rect 147674 460912 147680 460924
rect 147732 460912 147738 460964
rect 102192 460856 106274 460884
rect 102192 460844 102198 460856
rect 48130 460164 48136 460216
rect 48188 460204 48194 460216
rect 67634 460204 67640 460216
rect 48188 460176 67640 460204
rect 48188 460164 48194 460176
rect 67634 460164 67640 460176
rect 67692 460164 67698 460216
rect 102134 460164 102140 460216
rect 102192 460204 102198 460216
rect 106090 460204 106096 460216
rect 102192 460176 106096 460204
rect 102192 460164 102198 460176
rect 106090 460164 106096 460176
rect 106148 460204 106154 460216
rect 130010 460204 130016 460216
rect 106148 460176 130016 460204
rect 106148 460164 106154 460176
rect 130010 460164 130016 460176
rect 130068 460164 130074 460216
rect 111058 459620 111064 459672
rect 111116 459660 111122 459672
rect 119430 459660 119436 459672
rect 111116 459632 119436 459660
rect 111116 459620 111122 459632
rect 119430 459620 119436 459632
rect 119488 459620 119494 459672
rect 47670 459552 47676 459604
rect 47728 459592 47734 459604
rect 48130 459592 48136 459604
rect 47728 459564 48136 459592
rect 47728 459552 47734 459564
rect 48130 459552 48136 459564
rect 48188 459552 48194 459604
rect 102226 459552 102232 459604
rect 102284 459592 102290 459604
rect 103238 459592 103244 459604
rect 102284 459564 103244 459592
rect 102284 459552 102290 459564
rect 103238 459552 103244 459564
rect 103296 459592 103302 459604
rect 145006 459592 145012 459604
rect 103296 459564 145012 459592
rect 103296 459552 103302 459564
rect 145006 459552 145012 459564
rect 145064 459552 145070 459604
rect 63494 459484 63500 459536
rect 63552 459524 63558 459536
rect 64138 459524 64144 459536
rect 63552 459496 64144 459524
rect 63552 459484 63558 459496
rect 64138 459484 64144 459496
rect 64196 459524 64202 459536
rect 67634 459524 67640 459536
rect 64196 459496 67640 459524
rect 64196 459484 64202 459496
rect 67634 459484 67640 459496
rect 67692 459484 67698 459536
rect 102134 459484 102140 459536
rect 102192 459524 102198 459536
rect 111058 459524 111064 459536
rect 102192 459496 111064 459524
rect 102192 459484 102198 459496
rect 111058 459484 111064 459496
rect 111116 459484 111122 459536
rect 108298 458872 108304 458924
rect 108356 458912 108362 458924
rect 135254 458912 135260 458924
rect 108356 458884 135260 458912
rect 108356 458872 108362 458884
rect 135254 458872 135260 458884
rect 135312 458872 135318 458924
rect 32950 458804 32956 458856
rect 33008 458844 33014 458856
rect 63494 458844 63500 458856
rect 33008 458816 63500 458844
rect 33008 458804 33014 458816
rect 63494 458804 63500 458816
rect 63552 458804 63558 458856
rect 101306 458804 101312 458856
rect 101364 458844 101370 458856
rect 138658 458844 138664 458856
rect 101364 458816 138664 458844
rect 101364 458804 101370 458816
rect 138658 458804 138664 458816
rect 138716 458844 138722 458856
rect 142522 458844 142528 458856
rect 138716 458816 142528 458844
rect 138716 458804 138722 458816
rect 142522 458804 142528 458816
rect 142580 458804 142586 458856
rect 55858 458232 55864 458244
rect 55186 458204 55864 458232
rect 50338 458124 50344 458176
rect 50396 458164 50402 458176
rect 55186 458164 55214 458204
rect 55858 458192 55864 458204
rect 55916 458232 55922 458244
rect 67726 458232 67732 458244
rect 55916 458204 67732 458232
rect 55916 458192 55922 458204
rect 67726 458192 67732 458204
rect 67784 458192 67790 458244
rect 135254 458192 135260 458244
rect 135312 458232 135318 458244
rect 136910 458232 136916 458244
rect 135312 458204 136916 458232
rect 135312 458192 135318 458204
rect 136910 458192 136916 458204
rect 136968 458192 136974 458244
rect 50396 458136 55214 458164
rect 50396 458124 50402 458136
rect 39850 457512 39856 457564
rect 39908 457552 39914 457564
rect 50522 457552 50528 457564
rect 39908 457524 50528 457552
rect 39908 457512 39914 457524
rect 50522 457512 50528 457524
rect 50580 457512 50586 457564
rect 102226 457512 102232 457564
rect 102284 457552 102290 457564
rect 108298 457552 108304 457564
rect 102284 457524 108304 457552
rect 102284 457512 102290 457524
rect 108298 457512 108304 457524
rect 108356 457512 108362 457564
rect 34238 457444 34244 457496
rect 34296 457484 34302 457496
rect 36538 457484 36544 457496
rect 34296 457456 36544 457484
rect 34296 457444 34302 457456
rect 36538 457444 36544 457456
rect 36596 457484 36602 457496
rect 67634 457484 67640 457496
rect 36596 457456 67640 457484
rect 36596 457444 36602 457456
rect 67634 457444 67640 457456
rect 67692 457444 67698 457496
rect 103606 457444 103612 457496
rect 103664 457484 103670 457496
rect 142338 457484 142344 457496
rect 103664 457456 142344 457484
rect 103664 457444 103670 457456
rect 142338 457444 142344 457456
rect 142396 457484 142402 457496
rect 150526 457484 150532 457496
rect 142396 457456 150532 457484
rect 142396 457444 142402 457456
rect 150526 457444 150532 457456
rect 150584 457444 150590 457496
rect 50522 456764 50528 456816
rect 50580 456804 50586 456816
rect 50890 456804 50896 456816
rect 50580 456776 50896 456804
rect 50580 456764 50586 456776
rect 50890 456764 50896 456776
rect 50948 456804 50954 456816
rect 67634 456804 67640 456816
rect 50948 456776 67640 456804
rect 50948 456764 50954 456776
rect 67634 456764 67640 456776
rect 67692 456764 67698 456816
rect 108482 456764 108488 456816
rect 108540 456804 108546 456816
rect 108942 456804 108948 456816
rect 108540 456776 108948 456804
rect 108540 456764 108546 456776
rect 108942 456764 108948 456776
rect 109000 456804 109006 456816
rect 150434 456804 150440 456816
rect 109000 456776 150440 456804
rect 109000 456764 109006 456776
rect 150434 456764 150440 456776
rect 150492 456764 150498 456816
rect 446398 456764 446404 456816
rect 446456 456804 446462 456816
rect 580166 456804 580172 456816
rect 446456 456776 580172 456804
rect 446456 456764 446462 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 62114 456696 62120 456748
rect 62172 456736 62178 456748
rect 67726 456736 67732 456748
rect 62172 456708 67732 456736
rect 62172 456696 62178 456708
rect 67726 456696 67732 456708
rect 67784 456696 67790 456748
rect 35710 456016 35716 456068
rect 35768 456056 35774 456068
rect 62114 456056 62120 456068
rect 35768 456028 62120 456056
rect 35768 456016 35774 456028
rect 62114 456016 62120 456028
rect 62172 456016 62178 456068
rect 102870 456016 102876 456068
rect 102928 456056 102934 456068
rect 121546 456056 121552 456068
rect 102928 456028 121552 456056
rect 102928 456016 102934 456028
rect 121546 456016 121552 456028
rect 121604 456016 121610 456068
rect 56502 455336 56508 455388
rect 56560 455376 56566 455388
rect 57698 455376 57704 455388
rect 56560 455348 57704 455376
rect 56560 455336 56566 455348
rect 57698 455336 57704 455348
rect 57756 455336 57762 455388
rect 102134 455336 102140 455388
rect 102192 455376 102198 455388
rect 108482 455376 108488 455388
rect 102192 455348 108488 455376
rect 102192 455336 102198 455348
rect 108482 455336 108488 455348
rect 108540 455336 108546 455388
rect 108942 454928 108948 454980
rect 109000 454968 109006 454980
rect 111794 454968 111800 454980
rect 109000 454940 111800 454968
rect 109000 454928 109006 454940
rect 111794 454928 111800 454940
rect 111852 454928 111858 454980
rect 56502 454384 56508 454436
rect 56560 454424 56566 454436
rect 57238 454424 57244 454436
rect 56560 454396 57244 454424
rect 56560 454384 56566 454396
rect 57238 454384 57244 454396
rect 57296 454384 57302 454436
rect 57698 454044 57704 454096
rect 57756 454084 57762 454096
rect 67634 454084 67640 454096
rect 57756 454056 67640 454084
rect 57756 454044 57762 454056
rect 67634 454044 67640 454056
rect 67692 454044 67698 454096
rect 139578 454084 139584 454096
rect 108316 454056 139584 454084
rect 57606 453976 57612 454028
rect 57664 454016 57670 454028
rect 68002 454016 68008 454028
rect 57664 453988 68008 454016
rect 57664 453976 57670 453988
rect 68002 453976 68008 453988
rect 68060 453976 68066 454028
rect 102134 453976 102140 454028
rect 102192 454016 102198 454028
rect 108316 454016 108344 454056
rect 139578 454044 139584 454056
rect 139636 454044 139642 454096
rect 102192 453988 108344 454016
rect 102192 453976 102198 453988
rect 56502 453296 56508 453348
rect 56560 453336 56566 453348
rect 67634 453336 67640 453348
rect 56560 453308 67640 453336
rect 56560 453296 56566 453308
rect 67634 453296 67640 453308
rect 67692 453296 67698 453348
rect 102870 453296 102876 453348
rect 102928 453336 102934 453348
rect 118786 453336 118792 453348
rect 102928 453308 118792 453336
rect 102928 453296 102934 453308
rect 118786 453296 118792 453308
rect 118844 453296 118850 453348
rect 65610 452548 65616 452600
rect 65668 452588 65674 452600
rect 67634 452588 67640 452600
rect 65668 452560 67640 452588
rect 65668 452548 65674 452560
rect 67634 452548 67640 452560
rect 67692 452548 67698 452600
rect 45462 451868 45468 451920
rect 45520 451908 45526 451920
rect 46750 451908 46756 451920
rect 45520 451880 46756 451908
rect 45520 451868 45526 451880
rect 46750 451868 46756 451880
rect 46808 451908 46814 451920
rect 67358 451908 67364 451920
rect 46808 451880 67364 451908
rect 46808 451868 46814 451880
rect 67358 451868 67364 451880
rect 67416 451868 67422 451920
rect 102318 451868 102324 451920
rect 102376 451908 102382 451920
rect 116026 451908 116032 451920
rect 102376 451880 116032 451908
rect 102376 451868 102382 451880
rect 116026 451868 116032 451880
rect 116084 451868 116090 451920
rect 116026 451528 116032 451580
rect 116084 451568 116090 451580
rect 116578 451568 116584 451580
rect 116084 451540 116584 451568
rect 116084 451528 116090 451540
rect 116578 451528 116584 451540
rect 116636 451528 116642 451580
rect 30282 451256 30288 451308
rect 30340 451296 30346 451308
rect 33778 451296 33784 451308
rect 30340 451268 33784 451296
rect 30340 451256 30346 451268
rect 33778 451256 33784 451268
rect 33836 451256 33842 451308
rect 58986 451256 58992 451308
rect 59044 451296 59050 451308
rect 65610 451296 65616 451308
rect 59044 451268 65616 451296
rect 59044 451256 59050 451268
rect 65610 451256 65616 451268
rect 65668 451256 65674 451308
rect 102134 451256 102140 451308
rect 102192 451296 102198 451308
rect 139394 451296 139400 451308
rect 102192 451268 139400 451296
rect 102192 451256 102198 451268
rect 139394 451256 139400 451268
rect 139452 451256 139458 451308
rect 33796 451228 33824 451256
rect 67634 451228 67640 451240
rect 33796 451200 67640 451228
rect 67634 451188 67640 451200
rect 67692 451188 67698 451240
rect 107378 449896 107384 449948
rect 107436 449936 107442 449948
rect 138658 449936 138664 449948
rect 107436 449908 138664 449936
rect 107436 449896 107442 449908
rect 138658 449896 138664 449908
rect 138716 449896 138722 449948
rect 102134 449828 102140 449880
rect 102192 449868 102198 449880
rect 107396 449868 107424 449896
rect 102192 449840 107424 449868
rect 102192 449828 102198 449840
rect 102870 449216 102876 449268
rect 102928 449256 102934 449268
rect 106182 449256 106188 449268
rect 102928 449228 106188 449256
rect 102928 449216 102934 449228
rect 106182 449216 106188 449228
rect 106240 449256 106246 449268
rect 107654 449256 107660 449268
rect 106240 449228 107660 449256
rect 106240 449216 106246 449228
rect 107654 449216 107660 449228
rect 107712 449216 107718 449268
rect 105998 448672 106004 448724
rect 106056 448712 106062 448724
rect 123570 448712 123576 448724
rect 106056 448684 123576 448712
rect 106056 448672 106062 448684
rect 123570 448672 123576 448684
rect 123628 448672 123634 448724
rect 101582 448604 101588 448656
rect 101640 448644 101646 448656
rect 107470 448644 107476 448656
rect 101640 448616 107476 448644
rect 101640 448604 101646 448616
rect 107470 448604 107476 448616
rect 107528 448644 107534 448656
rect 113266 448644 113272 448656
rect 107528 448616 113272 448644
rect 107528 448604 107534 448616
rect 113266 448604 113272 448616
rect 113324 448604 113330 448656
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 58618 448576 58624 448588
rect 3200 448548 58624 448576
rect 3200 448536 3206 448548
rect 58618 448536 58624 448548
rect 58676 448536 58682 448588
rect 59262 448536 59268 448588
rect 59320 448576 59326 448588
rect 64138 448576 64144 448588
rect 59320 448548 64144 448576
rect 59320 448536 59326 448548
rect 64138 448536 64144 448548
rect 64196 448576 64202 448588
rect 67726 448576 67732 448588
rect 64196 448548 67732 448576
rect 64196 448536 64202 448548
rect 67726 448536 67732 448548
rect 67784 448536 67790 448588
rect 61930 448468 61936 448520
rect 61988 448508 61994 448520
rect 63402 448508 63408 448520
rect 61988 448480 63408 448508
rect 61988 448468 61994 448480
rect 63402 448468 63408 448480
rect 63460 448508 63466 448520
rect 67634 448508 67640 448520
rect 63460 448480 67640 448508
rect 63460 448468 63466 448480
rect 67634 448468 67640 448480
rect 67692 448468 67698 448520
rect 102134 448468 102140 448520
rect 102192 448508 102198 448520
rect 105630 448508 105636 448520
rect 102192 448480 105636 448508
rect 102192 448468 102198 448480
rect 105630 448468 105636 448480
rect 105688 448508 105694 448520
rect 105998 448508 106004 448520
rect 105688 448480 106004 448508
rect 105688 448468 105694 448480
rect 105998 448468 106004 448480
rect 106056 448468 106062 448520
rect 64782 447108 64788 447160
rect 64840 447148 64846 447160
rect 65610 447148 65616 447160
rect 64840 447120 65616 447148
rect 64840 447108 64846 447120
rect 65610 447108 65616 447120
rect 65668 447148 65674 447160
rect 67634 447148 67640 447160
rect 65668 447120 67640 447148
rect 65668 447108 65674 447120
rect 67634 447108 67640 447120
rect 67692 447108 67698 447160
rect 102226 447108 102232 447160
rect 102284 447148 102290 447160
rect 125870 447148 125876 447160
rect 102284 447120 125876 447148
rect 102284 447108 102290 447120
rect 125870 447108 125876 447120
rect 125928 447148 125934 447160
rect 131298 447148 131304 447160
rect 125928 447120 131304 447148
rect 125928 447108 125934 447120
rect 131298 447108 131304 447120
rect 131356 447108 131362 447160
rect 124214 446428 124220 446480
rect 124272 446468 124278 446480
rect 124398 446468 124404 446480
rect 124272 446440 124404 446468
rect 124272 446428 124278 446440
rect 124398 446428 124404 446440
rect 124456 446428 124462 446480
rect 104802 445816 104808 445868
rect 104860 445856 104866 445868
rect 112622 445856 112628 445868
rect 104860 445828 112628 445856
rect 104860 445816 104866 445828
rect 112622 445816 112628 445828
rect 112680 445816 112686 445868
rect 63126 445748 63132 445800
rect 63184 445788 63190 445800
rect 67634 445788 67640 445800
rect 63184 445760 67640 445788
rect 63184 445748 63190 445760
rect 67634 445748 67640 445760
rect 67692 445748 67698 445800
rect 102594 445748 102600 445800
rect 102652 445788 102658 445800
rect 135346 445788 135352 445800
rect 102652 445760 135352 445788
rect 102652 445748 102658 445760
rect 135346 445748 135352 445760
rect 135404 445748 135410 445800
rect 103238 445680 103244 445732
rect 103296 445720 103302 445732
rect 104802 445720 104808 445732
rect 103296 445692 104808 445720
rect 103296 445680 103302 445692
rect 104802 445680 104808 445692
rect 104860 445680 104866 445732
rect 102502 445612 102508 445664
rect 102560 445652 102566 445664
rect 104158 445652 104164 445664
rect 102560 445624 104164 445652
rect 102560 445612 102566 445624
rect 104158 445612 104164 445624
rect 104216 445612 104222 445664
rect 102226 445000 102232 445052
rect 102284 445040 102290 445052
rect 136634 445040 136640 445052
rect 102284 445012 136640 445040
rect 102284 445000 102290 445012
rect 136634 445000 136640 445012
rect 136692 445040 136698 445052
rect 142154 445040 142160 445052
rect 136692 445012 142160 445040
rect 136692 445000 136698 445012
rect 142154 445000 142160 445012
rect 142212 445000 142218 445052
rect 123478 444428 123484 444440
rect 122806 444400 123484 444428
rect 55674 444320 55680 444372
rect 55732 444360 55738 444372
rect 56410 444360 56416 444372
rect 55732 444332 56416 444360
rect 55732 444320 55738 444332
rect 56410 444320 56416 444332
rect 56468 444360 56474 444372
rect 67634 444360 67640 444372
rect 56468 444332 67640 444360
rect 56468 444320 56474 444332
rect 67634 444320 67640 444332
rect 67692 444320 67698 444372
rect 99650 444320 99656 444372
rect 99708 444360 99714 444372
rect 122806 444360 122834 444400
rect 123478 444388 123484 444400
rect 123536 444428 123542 444440
rect 129734 444428 129740 444440
rect 123536 444400 129740 444428
rect 123536 444388 123542 444400
rect 129734 444388 129740 444400
rect 129792 444388 129798 444440
rect 99708 444332 122834 444360
rect 99708 444320 99714 444332
rect 41322 443640 41328 443692
rect 41380 443680 41386 443692
rect 55674 443680 55680 443692
rect 41380 443652 55680 443680
rect 41380 443640 41386 443652
rect 55674 443640 55680 443652
rect 55732 443640 55738 443692
rect 60642 442892 60648 442944
rect 60700 442932 60706 442944
rect 64598 442932 64604 442944
rect 60700 442904 64604 442932
rect 60700 442892 60706 442904
rect 64598 442892 64604 442904
rect 64656 442892 64662 442944
rect 36998 442688 37004 442740
rect 37056 442728 37062 442740
rect 37182 442728 37188 442740
rect 37056 442700 37188 442728
rect 37056 442688 37062 442700
rect 37182 442688 37188 442700
rect 37240 442688 37246 442740
rect 36998 442212 37004 442264
rect 37056 442252 37062 442264
rect 67634 442252 67640 442264
rect 37056 442224 67640 442252
rect 37056 442212 37062 442224
rect 67634 442212 67640 442224
rect 67692 442212 67698 442264
rect 102870 442212 102876 442264
rect 102928 442252 102934 442264
rect 108758 442252 108764 442264
rect 102928 442224 108764 442252
rect 102928 442212 102934 442224
rect 108758 442212 108764 442224
rect 108816 442252 108822 442264
rect 130378 442252 130384 442264
rect 108816 442224 130384 442252
rect 108816 442212 108822 442224
rect 130378 442212 130384 442224
rect 130436 442212 130442 442264
rect 64598 441600 64604 441652
rect 64656 441640 64662 441652
rect 67726 441640 67732 441652
rect 64656 441612 67732 441640
rect 64656 441600 64662 441612
rect 67726 441600 67732 441612
rect 67784 441600 67790 441652
rect 63402 441532 63408 441584
rect 63460 441572 63466 441584
rect 63460 441544 64874 441572
rect 63460 441532 63466 441544
rect 64846 441504 64874 441544
rect 99282 441532 99288 441584
rect 99340 441572 99346 441584
rect 99374 441572 99380 441584
rect 99340 441544 99380 441572
rect 99340 441532 99346 441544
rect 99374 441532 99380 441544
rect 99432 441532 99438 441584
rect 65518 441504 65524 441516
rect 64846 441476 65524 441504
rect 65518 441464 65524 441476
rect 65576 441504 65582 441516
rect 67634 441504 67640 441516
rect 65576 441476 67640 441504
rect 65576 441464 65582 441476
rect 67634 441464 67640 441476
rect 67692 441464 67698 441516
rect 62022 440852 62028 440904
rect 62080 440892 62086 440904
rect 67634 440892 67640 440904
rect 62080 440864 67640 440892
rect 62080 440852 62086 440864
rect 67634 440852 67640 440864
rect 67692 440852 67698 440904
rect 117590 440892 117596 440904
rect 97920 440864 117596 440892
rect 97920 440700 97948 440864
rect 117590 440852 117596 440864
rect 117648 440852 117654 440904
rect 97902 440648 97908 440700
rect 97960 440648 97966 440700
rect 102594 440308 102600 440360
rect 102652 440348 102658 440360
rect 102652 440320 109034 440348
rect 102652 440308 102658 440320
rect 48038 440240 48044 440292
rect 48096 440280 48102 440292
rect 50982 440280 50988 440292
rect 48096 440252 50988 440280
rect 48096 440240 48102 440252
rect 50982 440240 50988 440252
rect 51040 440240 51046 440292
rect 61838 440240 61844 440292
rect 61896 440280 61902 440292
rect 62022 440280 62028 440292
rect 61896 440252 62028 440280
rect 61896 440240 61902 440252
rect 62022 440240 62028 440252
rect 62080 440240 62086 440292
rect 101490 440240 101496 440292
rect 101548 440280 101554 440292
rect 102042 440280 102048 440292
rect 101548 440252 102048 440280
rect 101548 440240 101554 440252
rect 102042 440240 102048 440252
rect 102100 440280 102106 440292
rect 105538 440280 105544 440292
rect 102100 440252 105544 440280
rect 102100 440240 102106 440252
rect 105538 440240 105544 440252
rect 105596 440240 105602 440292
rect 109006 440280 109034 440320
rect 133966 440280 133972 440292
rect 109006 440252 133972 440280
rect 133966 440240 133972 440252
rect 134024 440240 134030 440292
rect 64690 439560 64696 439612
rect 64748 439600 64754 439612
rect 75178 439600 75184 439612
rect 64748 439572 75184 439600
rect 64748 439560 64754 439572
rect 75178 439560 75184 439572
rect 75236 439560 75242 439612
rect 53742 439492 53748 439544
rect 53800 439532 53806 439544
rect 82814 439532 82820 439544
rect 53800 439504 82820 439532
rect 53800 439492 53806 439504
rect 82814 439492 82820 439504
rect 82872 439492 82878 439544
rect 69106 439220 69112 439272
rect 69164 439260 69170 439272
rect 71774 439260 71780 439272
rect 69164 439232 71780 439260
rect 69164 439220 69170 439232
rect 71774 439220 71780 439232
rect 71832 439220 71838 439272
rect 11698 439152 11704 439204
rect 11756 439192 11762 439204
rect 96430 439192 96436 439204
rect 11756 439164 96436 439192
rect 11756 439152 11762 439164
rect 96430 439152 96436 439164
rect 96488 439152 96494 439204
rect 88702 439084 88708 439136
rect 88760 439124 88766 439136
rect 121546 439124 121552 439136
rect 88760 439096 121552 439124
rect 88760 439084 88766 439096
rect 121546 439084 121552 439096
rect 121604 439084 121610 439136
rect 125502 439084 125508 439136
rect 125560 439124 125566 439136
rect 132678 439124 132684 439136
rect 125560 439096 132684 439124
rect 125560 439084 125566 439096
rect 132678 439084 132684 439096
rect 132736 439084 132742 439136
rect 94498 439016 94504 439068
rect 94556 439056 94562 439068
rect 128446 439056 128452 439068
rect 94556 439028 128452 439056
rect 94556 439016 94562 439028
rect 128446 439016 128452 439028
rect 128504 439056 128510 439068
rect 131482 439056 131488 439068
rect 128504 439028 131488 439056
rect 128504 439016 128510 439028
rect 131482 439016 131488 439028
rect 131540 439016 131546 439068
rect 39758 438948 39764 439000
rect 39816 438988 39822 439000
rect 39816 438960 64874 438988
rect 39816 438948 39822 438960
rect 64846 438920 64874 438960
rect 92474 438948 92480 439000
rect 92532 438988 92538 439000
rect 93210 438988 93216 439000
rect 92532 438960 93216 438988
rect 92532 438948 92538 438960
rect 93210 438948 93216 438960
rect 93268 438988 93274 439000
rect 131114 438988 131120 439000
rect 93268 438960 131120 438988
rect 93268 438948 93274 438960
rect 131114 438948 131120 438960
rect 131172 438948 131178 439000
rect 72602 438920 72608 438932
rect 64846 438892 72608 438920
rect 72602 438880 72608 438892
rect 72660 438920 72666 438932
rect 73338 438920 73344 438932
rect 72660 438892 73344 438920
rect 72660 438880 72666 438892
rect 73338 438880 73344 438892
rect 73396 438880 73402 438932
rect 119338 438880 119344 438932
rect 119396 438920 119402 438932
rect 136818 438920 136824 438932
rect 119396 438892 136824 438920
rect 119396 438880 119402 438892
rect 136818 438880 136824 438892
rect 136876 438880 136882 438932
rect 4798 438812 4804 438864
rect 4856 438852 4862 438864
rect 49602 438852 49608 438864
rect 4856 438824 49608 438852
rect 4856 438812 4862 438824
rect 49602 438812 49608 438824
rect 49660 438812 49666 438864
rect 99650 438812 99656 438864
rect 99708 438852 99714 438864
rect 124858 438852 124864 438864
rect 99708 438824 124864 438852
rect 99708 438812 99714 438824
rect 124858 438812 124864 438824
rect 124916 438852 124922 438864
rect 125502 438852 125508 438864
rect 124916 438824 125508 438852
rect 124916 438812 124922 438824
rect 125502 438812 125508 438824
rect 125560 438812 125566 438864
rect 46658 438744 46664 438796
rect 46716 438784 46722 438796
rect 78766 438784 78772 438796
rect 46716 438756 78772 438784
rect 46716 438744 46722 438756
rect 78766 438744 78772 438756
rect 78824 438744 78830 438796
rect 82814 438744 82820 438796
rect 82872 438784 82878 438796
rect 83458 438784 83464 438796
rect 82872 438756 83464 438784
rect 82872 438744 82878 438756
rect 83458 438744 83464 438756
rect 83516 438784 83522 438796
rect 87414 438784 87420 438796
rect 83516 438756 87420 438784
rect 83516 438744 83522 438756
rect 87414 438744 87420 438756
rect 87472 438744 87478 438796
rect 91278 438744 91284 438796
rect 91336 438784 91342 438796
rect 124214 438784 124220 438796
rect 91336 438756 124220 438784
rect 91336 438744 91342 438756
rect 124214 438744 124220 438756
rect 124272 438784 124278 438796
rect 124398 438784 124404 438796
rect 124272 438756 124404 438784
rect 124272 438744 124278 438756
rect 124398 438744 124404 438756
rect 124456 438744 124462 438796
rect 57882 438676 57888 438728
rect 57940 438716 57946 438728
rect 82262 438716 82268 438728
rect 57940 438688 82268 438716
rect 57940 438676 57946 438688
rect 82262 438676 82268 438688
rect 82320 438676 82326 438728
rect 96430 438676 96436 438728
rect 96488 438716 96494 438728
rect 125778 438716 125784 438728
rect 96488 438688 125784 438716
rect 96488 438676 96494 438688
rect 125778 438676 125784 438688
rect 125836 438676 125842 438728
rect 51718 438608 51724 438660
rect 51776 438648 51782 438660
rect 73890 438648 73896 438660
rect 51776 438620 73896 438648
rect 51776 438608 51782 438620
rect 73890 438608 73896 438620
rect 73948 438608 73954 438660
rect 99006 438608 99012 438660
rect 99064 438648 99070 438660
rect 119338 438648 119344 438660
rect 99064 438620 119344 438648
rect 99064 438608 99070 438620
rect 119338 438608 119344 438620
rect 119396 438608 119402 438660
rect 91002 438540 91008 438592
rect 91060 438580 91066 438592
rect 100018 438580 100024 438592
rect 91060 438552 100024 438580
rect 91060 438540 91066 438552
rect 100018 438540 100024 438552
rect 100076 438540 100082 438592
rect 93854 438472 93860 438524
rect 93912 438512 93918 438524
rect 95142 438512 95148 438524
rect 93912 438484 95148 438512
rect 93912 438472 93918 438484
rect 95142 438472 95148 438484
rect 95200 438512 95206 438524
rect 103514 438512 103520 438524
rect 95200 438484 103520 438512
rect 95200 438472 95206 438484
rect 103514 438472 103520 438484
rect 103572 438472 103578 438524
rect 58618 438404 58624 438456
rect 58676 438444 58682 438456
rect 99742 438444 99748 438456
rect 58676 438416 99748 438444
rect 58676 438404 58682 438416
rect 99742 438404 99748 438416
rect 99800 438404 99806 438456
rect 45186 438268 45192 438320
rect 45244 438308 45250 438320
rect 51718 438308 51724 438320
rect 45244 438280 51724 438308
rect 45244 438268 45250 438280
rect 51718 438268 51724 438280
rect 51776 438268 51782 438320
rect 45554 438200 45560 438252
rect 45612 438240 45618 438252
rect 46198 438240 46204 438252
rect 45612 438212 46204 438240
rect 45612 438200 45618 438212
rect 46198 438200 46204 438212
rect 46256 438240 46262 438252
rect 73246 438240 73252 438252
rect 46256 438212 73252 438240
rect 46256 438200 46262 438212
rect 73246 438200 73252 438212
rect 73304 438200 73310 438252
rect 49602 438132 49608 438184
rect 49660 438172 49666 438184
rect 50706 438172 50712 438184
rect 49660 438144 50712 438172
rect 49660 438132 49666 438144
rect 50706 438132 50712 438144
rect 50764 438172 50770 438184
rect 83550 438172 83556 438184
rect 50764 438144 83556 438172
rect 50764 438132 50770 438144
rect 83550 438132 83556 438144
rect 83608 438132 83614 438184
rect 89990 438132 89996 438184
rect 90048 438172 90054 438184
rect 91002 438172 91008 438184
rect 90048 438144 91008 438172
rect 90048 438132 90054 438144
rect 91002 438132 91008 438144
rect 91060 438132 91066 438184
rect 97718 437996 97724 438048
rect 97776 438036 97782 438048
rect 98638 438036 98644 438048
rect 97776 438008 98644 438036
rect 97776 437996 97782 438008
rect 98638 437996 98644 438008
rect 98696 437996 98702 438048
rect 86770 437452 86776 437504
rect 86828 437492 86834 437504
rect 87598 437492 87604 437504
rect 86828 437464 87604 437492
rect 86828 437452 86834 437464
rect 87598 437452 87604 437464
rect 87656 437452 87662 437504
rect 97442 437384 97448 437436
rect 97500 437424 97506 437436
rect 127158 437424 127164 437436
rect 97500 437396 127164 437424
rect 97500 437384 97506 437396
rect 127158 437384 127164 437396
rect 127216 437384 127222 437436
rect 46474 437316 46480 437368
rect 46532 437356 46538 437368
rect 80974 437356 80980 437368
rect 46532 437328 80980 437356
rect 46532 437316 46538 437328
rect 80974 437316 80980 437328
rect 81032 437316 81038 437368
rect 88242 437316 88248 437368
rect 88300 437356 88306 437368
rect 108390 437356 108396 437368
rect 88300 437328 108396 437356
rect 88300 437316 88306 437328
rect 108390 437316 108396 437328
rect 108448 437316 108454 437368
rect 50614 437248 50620 437300
rect 50672 437288 50678 437300
rect 82906 437288 82912 437300
rect 50672 437260 82912 437288
rect 50672 437248 50678 437260
rect 82906 437248 82912 437260
rect 82964 437248 82970 437300
rect 88978 437248 88984 437300
rect 89036 437288 89042 437300
rect 104894 437288 104900 437300
rect 89036 437260 104900 437288
rect 89036 437248 89042 437260
rect 104894 437248 104900 437260
rect 104952 437248 104958 437300
rect 43990 437180 43996 437232
rect 44048 437220 44054 437232
rect 77938 437220 77944 437232
rect 44048 437192 77944 437220
rect 44048 437180 44054 437192
rect 77938 437180 77944 437192
rect 77996 437220 78002 437232
rect 78398 437220 78404 437232
rect 77996 437192 78404 437220
rect 77996 437180 78002 437192
rect 78398 437180 78404 437192
rect 78456 437180 78462 437232
rect 80146 436432 80152 436484
rect 80204 436472 80210 436484
rect 80974 436472 80980 436484
rect 80204 436444 80980 436472
rect 80204 436432 80210 436444
rect 80974 436432 80980 436444
rect 81032 436432 81038 436484
rect 120258 436092 120264 436144
rect 120316 436132 120322 436144
rect 120718 436132 120724 436144
rect 120316 436104 120724 436132
rect 120316 436092 120322 436104
rect 120718 436092 120724 436104
rect 120776 436132 120782 436144
rect 128446 436132 128452 436144
rect 120776 436104 128452 436132
rect 120776 436092 120782 436104
rect 128446 436092 128452 436104
rect 128504 436092 128510 436144
rect 45278 436024 45284 436076
rect 45336 436064 45342 436076
rect 45462 436064 45468 436076
rect 45336 436036 45468 436064
rect 45336 436024 45342 436036
rect 45462 436024 45468 436036
rect 45520 436064 45526 436076
rect 76466 436064 76472 436076
rect 45520 436036 76472 436064
rect 45520 436024 45526 436036
rect 76466 436024 76472 436036
rect 76524 436024 76530 436076
rect 95050 436024 95056 436076
rect 95108 436064 95114 436076
rect 125686 436064 125692 436076
rect 95108 436036 125692 436064
rect 95108 436024 95114 436036
rect 125686 436024 125692 436036
rect 125744 436024 125750 436076
rect 56318 435956 56324 436008
rect 56376 435996 56382 436008
rect 81434 435996 81440 436008
rect 56376 435968 81440 435996
rect 56376 435956 56382 435968
rect 81434 435956 81440 435968
rect 81492 435956 81498 436008
rect 91922 435956 91928 436008
rect 91980 435996 91986 436008
rect 120258 435996 120264 436008
rect 91980 435968 120264 435996
rect 91980 435956 91986 435968
rect 120258 435956 120264 435968
rect 120316 435956 120322 436008
rect 57330 435888 57336 435940
rect 57388 435928 57394 435940
rect 76006 435928 76012 435940
rect 57388 435900 76012 435928
rect 57388 435888 57394 435900
rect 76006 435888 76012 435900
rect 76064 435928 76070 435940
rect 77110 435928 77116 435940
rect 76064 435900 77116 435928
rect 76064 435888 76070 435900
rect 77110 435888 77116 435900
rect 77168 435888 77174 435940
rect 48130 435344 48136 435396
rect 48188 435384 48194 435396
rect 71314 435384 71320 435396
rect 48188 435356 71320 435384
rect 48188 435344 48194 435356
rect 71314 435344 71320 435356
rect 71372 435344 71378 435396
rect 42702 434664 42708 434716
rect 42760 434704 42766 434716
rect 74718 434704 74724 434716
rect 42760 434676 74724 434704
rect 42760 434664 42766 434676
rect 74718 434664 74724 434676
rect 74776 434704 74782 434716
rect 75822 434704 75828 434716
rect 74776 434676 75828 434704
rect 74776 434664 74782 434676
rect 75822 434664 75828 434676
rect 75880 434664 75886 434716
rect 37090 434596 37096 434648
rect 37148 434636 37154 434648
rect 47578 434636 47584 434648
rect 37148 434608 47584 434636
rect 37148 434596 37154 434608
rect 47578 434596 47584 434608
rect 47636 434636 47642 434648
rect 48130 434636 48136 434648
rect 47636 434608 48136 434636
rect 47636 434596 47642 434608
rect 48130 434596 48136 434608
rect 48188 434596 48194 434648
rect 43806 433236 43812 433288
rect 43864 433276 43870 433288
rect 44082 433276 44088 433288
rect 43864 433248 44088 433276
rect 43864 433236 43870 433248
rect 44082 433236 44088 433248
rect 44140 433276 44146 433288
rect 74534 433276 74540 433288
rect 44140 433248 74540 433276
rect 44140 433236 44146 433248
rect 74534 433236 74540 433248
rect 74592 433236 74598 433288
rect 42702 432556 42708 432608
rect 42760 432596 42766 432608
rect 70670 432596 70676 432608
rect 42760 432568 70676 432596
rect 42760 432556 42766 432568
rect 70670 432556 70676 432568
rect 70728 432556 70734 432608
rect 38470 431876 38476 431928
rect 38528 431916 38534 431928
rect 42702 431916 42708 431928
rect 38528 431888 42708 431916
rect 38528 431876 38534 431888
rect 42702 431876 42708 431888
rect 42760 431876 42766 431928
rect 77938 431196 77944 431248
rect 77996 431236 78002 431248
rect 580166 431236 580172 431248
rect 77996 431208 580172 431236
rect 77996 431196 78002 431208
rect 580166 431196 580172 431208
rect 580224 431196 580230 431248
rect 42058 430584 42064 430636
rect 42116 430624 42122 430636
rect 42702 430624 42708 430636
rect 42116 430596 42708 430624
rect 42116 430584 42122 430596
rect 42702 430584 42708 430596
rect 42760 430584 42766 430636
rect 3418 429836 3424 429888
rect 3476 429876 3482 429888
rect 101582 429876 101588 429888
rect 3476 429848 101588 429876
rect 3476 429836 3482 429848
rect 101582 429836 101588 429848
rect 101640 429836 101646 429888
rect 3510 422288 3516 422340
rect 3568 422328 3574 422340
rect 3568 422300 111840 422328
rect 3568 422288 3574 422300
rect 111812 422260 111840 422300
rect 120166 422260 120172 422272
rect 111812 422232 120172 422260
rect 120166 422220 120172 422232
rect 120224 422220 120230 422272
rect 323578 418140 323584 418192
rect 323636 418180 323642 418192
rect 580166 418180 580172 418192
rect 323636 418152 580172 418180
rect 323636 418140 323642 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 59170 410524 59176 410576
rect 59228 410564 59234 410576
rect 89714 410564 89720 410576
rect 59228 410536 89720 410564
rect 59228 410524 59234 410536
rect 89714 410524 89720 410536
rect 89772 410524 89778 410576
rect 89714 409844 89720 409896
rect 89772 409884 89778 409896
rect 353294 409884 353300 409896
rect 89772 409856 353300 409884
rect 89772 409844 89778 409856
rect 353294 409844 353300 409856
rect 353352 409844 353358 409896
rect 40954 406376 40960 406428
rect 41012 406416 41018 406428
rect 71682 406416 71688 406428
rect 41012 406388 71688 406416
rect 41012 406376 41018 406388
rect 71682 406376 71688 406388
rect 71740 406376 71746 406428
rect 89806 406376 89812 406428
rect 89864 406416 89870 406428
rect 114646 406416 114652 406428
rect 89864 406388 114652 406416
rect 89864 406376 89870 406388
rect 114646 406376 114652 406388
rect 114704 406416 114710 406428
rect 115842 406416 115848 406428
rect 114704 406388 115848 406416
rect 114704 406376 114710 406388
rect 115842 406376 115848 406388
rect 115900 406376 115906 406428
rect 92474 405016 92480 405068
rect 92532 405056 92538 405068
rect 131298 405056 131304 405068
rect 92532 405028 131304 405056
rect 92532 405016 92538 405028
rect 131298 405016 131304 405028
rect 131356 405016 131362 405068
rect 106090 404948 106096 405000
rect 106148 404988 106154 405000
rect 145190 404988 145196 405000
rect 106148 404960 145196 404988
rect 106148 404948 106154 404960
rect 145190 404948 145196 404960
rect 145248 404948 145254 405000
rect 544378 404336 544384 404388
rect 544436 404376 544442 404388
rect 580166 404376 580172 404388
rect 544436 404348 580172 404376
rect 544436 404336 544442 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 36630 403588 36636 403640
rect 36688 403628 36694 403640
rect 75914 403628 75920 403640
rect 36688 403600 75920 403628
rect 36688 403588 36694 403600
rect 75914 403588 75920 403600
rect 75972 403588 75978 403640
rect 75914 403044 75920 403096
rect 75972 403084 75978 403096
rect 164878 403084 164884 403096
rect 75972 403056 164884 403084
rect 75972 403044 75978 403056
rect 164878 403044 164884 403056
rect 164936 403044 164942 403096
rect 67450 402976 67456 403028
rect 67508 403016 67514 403028
rect 367094 403016 367100 403028
rect 67508 402988 367100 403016
rect 67508 402976 67514 402988
rect 367094 402976 367100 402988
rect 367152 402976 367158 403028
rect 64782 401616 64788 401668
rect 64840 401656 64846 401668
rect 162118 401656 162124 401668
rect 64840 401628 162124 401656
rect 64840 401616 64846 401628
rect 162118 401616 162124 401628
rect 162176 401616 162182 401668
rect 35526 400936 35532 400988
rect 35584 400976 35590 400988
rect 70394 400976 70400 400988
rect 35584 400948 70400 400976
rect 35584 400936 35590 400948
rect 70394 400936 70400 400948
rect 70452 400936 70458 400988
rect 34422 400868 34428 400920
rect 34480 400908 34486 400920
rect 42794 400908 42800 400920
rect 34480 400880 42800 400908
rect 34480 400868 34486 400880
rect 42794 400868 42800 400880
rect 42852 400908 42858 400920
rect 80054 400908 80060 400920
rect 42852 400880 80060 400908
rect 42852 400868 42858 400880
rect 80054 400868 80060 400880
rect 80112 400868 80118 400920
rect 70394 400256 70400 400308
rect 70452 400296 70458 400308
rect 74534 400296 74540 400308
rect 70452 400268 74540 400296
rect 70452 400256 70458 400268
rect 74534 400256 74540 400268
rect 74592 400296 74598 400308
rect 153838 400296 153844 400308
rect 74592 400268 153844 400296
rect 74592 400256 74598 400268
rect 153838 400256 153844 400268
rect 153896 400256 153902 400308
rect 80054 400188 80060 400240
rect 80112 400228 80118 400240
rect 80238 400228 80244 400240
rect 80112 400200 80244 400228
rect 80112 400188 80118 400200
rect 80238 400188 80244 400200
rect 80296 400228 80302 400240
rect 320266 400228 320272 400240
rect 80296 400200 320272 400228
rect 80296 400188 80302 400200
rect 320266 400188 320272 400200
rect 320324 400188 320330 400240
rect 49418 399576 49424 399628
rect 49476 399616 49482 399628
rect 81434 399616 81440 399628
rect 49476 399588 81440 399616
rect 49476 399576 49482 399588
rect 81434 399576 81440 399588
rect 81492 399576 81498 399628
rect 52270 399508 52276 399560
rect 52328 399548 52334 399560
rect 88058 399548 88064 399560
rect 52328 399520 88064 399548
rect 52328 399508 52334 399520
rect 88058 399508 88064 399520
rect 88116 399508 88122 399560
rect 41046 399440 41052 399492
rect 41104 399480 41110 399492
rect 84930 399480 84936 399492
rect 41104 399452 84936 399480
rect 41104 399440 41110 399452
rect 84930 399440 84936 399452
rect 84988 399440 84994 399492
rect 95878 399440 95884 399492
rect 95936 399480 95942 399492
rect 108850 399480 108856 399492
rect 95936 399452 108856 399480
rect 95936 399440 95942 399452
rect 108850 399440 108856 399452
rect 108908 399480 108914 399492
rect 160738 399480 160744 399492
rect 108908 399452 160744 399480
rect 108908 399440 108914 399452
rect 160738 399440 160744 399452
rect 160796 399440 160802 399492
rect 87690 398964 87696 399016
rect 87748 399004 87754 399016
rect 88058 399004 88064 399016
rect 87748 398976 88064 399004
rect 87748 398964 87754 398976
rect 88058 398964 88064 398976
rect 88116 399004 88122 399016
rect 159358 399004 159364 399016
rect 88116 398976 159364 399004
rect 88116 398964 88122 398976
rect 159358 398964 159364 398976
rect 159416 398964 159422 399016
rect 68646 398896 68652 398948
rect 68704 398936 68710 398948
rect 228358 398936 228364 398948
rect 68704 398908 228364 398936
rect 68704 398896 68710 398908
rect 228358 398896 228364 398908
rect 228416 398896 228422 398948
rect 106274 398828 106280 398880
rect 106332 398868 106338 398880
rect 106918 398868 106924 398880
rect 106332 398840 106924 398868
rect 106332 398828 106338 398840
rect 106918 398828 106924 398840
rect 106976 398868 106982 398880
rect 358814 398868 358820 398880
rect 106976 398840 358820 398868
rect 106976 398828 106982 398840
rect 358814 398828 358820 398840
rect 358872 398828 358878 398880
rect 109862 398760 109868 398812
rect 109920 398800 109926 398812
rect 114094 398800 114100 398812
rect 109920 398772 114100 398800
rect 109920 398760 109926 398772
rect 114094 398760 114100 398772
rect 114152 398760 114158 398812
rect 53466 398148 53472 398200
rect 53524 398188 53530 398200
rect 85758 398188 85764 398200
rect 53524 398160 85764 398188
rect 53524 398148 53530 398160
rect 85758 398148 85764 398160
rect 85816 398148 85822 398200
rect 95050 398148 95056 398200
rect 95108 398188 95114 398200
rect 119614 398188 119620 398200
rect 95108 398160 119620 398188
rect 95108 398148 95114 398160
rect 119614 398148 119620 398160
rect 119672 398148 119678 398200
rect 51994 398080 52000 398132
rect 52052 398120 52058 398132
rect 87598 398120 87604 398132
rect 52052 398092 87604 398120
rect 52052 398080 52058 398092
rect 87598 398080 87604 398092
rect 87656 398080 87662 398132
rect 88334 398080 88340 398132
rect 88392 398120 88398 398132
rect 122834 398120 122840 398132
rect 88392 398092 122840 398120
rect 88392 398080 88398 398092
rect 122834 398080 122840 398092
rect 122892 398120 122898 398132
rect 157978 398120 157984 398132
rect 122892 398092 157984 398120
rect 122892 398080 122898 398092
rect 157978 398080 157984 398092
rect 158036 398080 158042 398132
rect 268378 397508 268384 397520
rect 69492 397480 268384 397508
rect 42610 397400 42616 397452
rect 42668 397440 42674 397452
rect 69198 397440 69204 397452
rect 42668 397412 69204 397440
rect 42668 397400 42674 397412
rect 69198 397400 69204 397412
rect 69256 397440 69262 397452
rect 69492 397440 69520 397480
rect 268378 397468 268384 397480
rect 268436 397468 268442 397520
rect 69256 397412 69520 397440
rect 69256 397400 69262 397412
rect 107470 396856 107476 396908
rect 107528 396896 107534 396908
rect 129826 396896 129832 396908
rect 107528 396868 129832 396896
rect 107528 396856 107534 396868
rect 129826 396856 129832 396868
rect 129884 396856 129890 396908
rect 57790 396788 57796 396840
rect 57848 396828 57854 396840
rect 83458 396828 83464 396840
rect 57848 396800 83464 396828
rect 57848 396788 57854 396800
rect 83458 396788 83464 396800
rect 83516 396788 83522 396840
rect 97810 396788 97816 396840
rect 97868 396828 97874 396840
rect 127250 396828 127256 396840
rect 97868 396800 127256 396828
rect 97868 396788 97874 396800
rect 127250 396788 127256 396800
rect 127308 396788 127314 396840
rect 46842 396720 46848 396772
rect 46900 396760 46906 396772
rect 78766 396760 78772 396772
rect 46900 396732 78772 396760
rect 46900 396720 46906 396732
rect 78766 396720 78772 396732
rect 78824 396720 78830 396772
rect 93946 396720 93952 396772
rect 94004 396760 94010 396772
rect 128538 396760 128544 396772
rect 94004 396732 128544 396760
rect 94004 396720 94010 396732
rect 128538 396720 128544 396732
rect 128596 396760 128602 396772
rect 154666 396760 154672 396772
rect 128596 396732 154672 396760
rect 128596 396720 128602 396732
rect 154666 396720 154672 396732
rect 154724 396720 154730 396772
rect 108298 396652 108304 396704
rect 108356 396692 108362 396704
rect 114554 396692 114560 396704
rect 108356 396664 114560 396692
rect 108356 396652 108362 396664
rect 114554 396652 114560 396664
rect 114612 396652 114618 396704
rect 129826 396108 129832 396160
rect 129884 396148 129890 396160
rect 130010 396148 130016 396160
rect 129884 396120 130016 396148
rect 129884 396108 129890 396120
rect 130010 396108 130016 396120
rect 130068 396148 130074 396160
rect 289078 396148 289084 396160
rect 130068 396120 289084 396148
rect 130068 396108 130074 396120
rect 289078 396108 289084 396120
rect 289136 396108 289142 396160
rect 55950 396080 55956 396092
rect 55186 396052 55956 396080
rect 46750 395972 46756 396024
rect 46808 396012 46814 396024
rect 55186 396012 55214 396052
rect 55950 396040 55956 396052
rect 56008 396080 56014 396092
rect 286318 396080 286324 396092
rect 56008 396052 286324 396080
rect 56008 396040 56014 396052
rect 286318 396040 286324 396052
rect 286376 396040 286382 396092
rect 46808 395984 55214 396012
rect 46808 395972 46814 395984
rect 96706 395292 96712 395344
rect 96764 395332 96770 395344
rect 130194 395332 130200 395344
rect 96764 395304 130200 395332
rect 96764 395292 96770 395304
rect 130194 395292 130200 395304
rect 130252 395332 130258 395344
rect 149146 395332 149152 395344
rect 130252 395304 149152 395332
rect 130252 395292 130258 395304
rect 149146 395292 149152 395304
rect 149204 395292 149210 395344
rect 39298 394748 39304 394800
rect 39356 394788 39362 394800
rect 115842 394788 115848 394800
rect 39356 394760 115848 394788
rect 39356 394748 39362 394760
rect 115842 394748 115848 394760
rect 115900 394748 115906 394800
rect 118786 394748 118792 394800
rect 118844 394788 118850 394800
rect 119982 394788 119988 394800
rect 118844 394760 119988 394788
rect 118844 394748 118850 394760
rect 119982 394748 119988 394760
rect 120040 394788 120046 394800
rect 122834 394788 122840 394800
rect 120040 394760 122840 394788
rect 120040 394748 120046 394760
rect 122834 394748 122840 394760
rect 122892 394748 122898 394800
rect 291838 394748 291844 394800
rect 291896 394788 291902 394800
rect 385678 394788 385684 394800
rect 291896 394760 385684 394788
rect 291896 394748 291902 394760
rect 385678 394748 385684 394760
rect 385736 394748 385742 394800
rect 55858 394680 55864 394732
rect 55916 394720 55922 394732
rect 64690 394720 64696 394732
rect 55916 394692 64696 394720
rect 55916 394680 55922 394692
rect 64690 394680 64696 394692
rect 64748 394720 64754 394732
rect 151814 394720 151820 394732
rect 64748 394692 151820 394720
rect 64748 394680 64754 394692
rect 151814 394680 151820 394692
rect 151872 394720 151878 394732
rect 304258 394720 304264 394732
rect 151872 394692 304264 394720
rect 151872 394680 151878 394692
rect 304258 394680 304264 394692
rect 304316 394680 304322 394732
rect 68738 394612 68744 394664
rect 68796 394652 68802 394664
rect 68922 394652 68928 394664
rect 68796 394624 68928 394652
rect 68796 394612 68802 394624
rect 68922 394612 68928 394624
rect 68980 394612 68986 394664
rect 115842 394612 115848 394664
rect 115900 394652 115906 394664
rect 118786 394652 118792 394664
rect 115900 394624 118792 394652
rect 115900 394612 115906 394624
rect 118786 394612 118792 394624
rect 118844 394612 118850 394664
rect 52086 394068 52092 394120
rect 52144 394108 52150 394120
rect 74718 394108 74724 394120
rect 52144 394080 74724 394108
rect 52144 394068 52150 394080
rect 74718 394068 74724 394080
rect 74776 394068 74782 394120
rect 110506 394068 110512 394120
rect 110564 394108 110570 394120
rect 130102 394108 130108 394120
rect 110564 394080 130108 394108
rect 110564 394068 110570 394080
rect 130102 394068 130108 394080
rect 130160 394108 130166 394120
rect 138106 394108 138112 394120
rect 130160 394080 138112 394108
rect 130160 394068 130166 394080
rect 138106 394068 138112 394080
rect 138164 394068 138170 394120
rect 54754 394000 54760 394052
rect 54812 394040 54818 394052
rect 82814 394040 82820 394052
rect 54812 394012 82820 394040
rect 54812 394000 54818 394012
rect 82814 394000 82820 394012
rect 82872 394000 82878 394052
rect 100662 394000 100668 394052
rect 100720 394040 100726 394052
rect 107654 394040 107660 394052
rect 100720 394012 107660 394040
rect 100720 394000 100726 394012
rect 107654 394000 107660 394012
rect 107712 394000 107718 394052
rect 108758 394000 108764 394052
rect 108816 394040 108822 394052
rect 131390 394040 131396 394052
rect 108816 394012 131396 394040
rect 108816 394000 108822 394012
rect 131390 394000 131396 394012
rect 131448 394000 131454 394052
rect 47854 393932 47860 393984
rect 47912 393972 47918 393984
rect 81434 393972 81440 393984
rect 47912 393944 81440 393972
rect 47912 393932 47918 393944
rect 81434 393932 81440 393944
rect 81492 393932 81498 393984
rect 95786 393932 95792 393984
rect 95844 393972 95850 393984
rect 127342 393972 127348 393984
rect 95844 393944 127348 393972
rect 95844 393932 95850 393944
rect 127342 393932 127348 393944
rect 127400 393972 127406 393984
rect 151998 393972 152004 393984
rect 127400 393944 152004 393972
rect 127400 393932 127406 393944
rect 151998 393932 152004 393944
rect 152056 393932 152062 393984
rect 82998 393456 83004 393508
rect 83056 393496 83062 393508
rect 146938 393496 146944 393508
rect 83056 393468 146944 393496
rect 83056 393456 83062 393468
rect 146938 393456 146944 393468
rect 146996 393456 147002 393508
rect 131390 393388 131396 393440
rect 131448 393428 131454 393440
rect 316678 393428 316684 393440
rect 131448 393400 316684 393428
rect 131448 393388 131454 393400
rect 316678 393388 316684 393400
rect 316736 393388 316742 393440
rect 68922 393320 68928 393372
rect 68980 393360 68986 393372
rect 278038 393360 278044 393372
rect 68980 393332 278044 393360
rect 68980 393320 68986 393332
rect 278038 393320 278044 393332
rect 278096 393320 278102 393372
rect 46750 392640 46756 392692
rect 46808 392680 46814 392692
rect 77294 392680 77300 392692
rect 46808 392652 77300 392680
rect 46808 392640 46814 392652
rect 77294 392640 77300 392652
rect 77352 392640 77358 392692
rect 106182 392640 106188 392692
rect 106240 392680 106246 392692
rect 131206 392680 131212 392692
rect 106240 392652 131212 392680
rect 106240 392640 106246 392652
rect 131206 392640 131212 392652
rect 131264 392680 131270 392692
rect 131264 392652 132494 392680
rect 131264 392640 131270 392652
rect 3418 392572 3424 392624
rect 3476 392612 3482 392624
rect 52454 392612 52460 392624
rect 3476 392584 52460 392612
rect 3476 392572 3482 392584
rect 52454 392572 52460 392584
rect 52512 392572 52518 392624
rect 56410 392572 56416 392624
rect 56468 392612 56474 392624
rect 86218 392612 86224 392624
rect 56468 392584 86224 392612
rect 56468 392572 56474 392584
rect 86218 392572 86224 392584
rect 86276 392572 86282 392624
rect 91002 392572 91008 392624
rect 91060 392612 91066 392624
rect 120258 392612 120264 392624
rect 91060 392584 120264 392612
rect 91060 392572 91066 392584
rect 120258 392572 120264 392584
rect 120316 392572 120322 392624
rect 132466 392612 132494 392652
rect 146294 392612 146300 392624
rect 132466 392584 146300 392612
rect 146294 392572 146300 392584
rect 146352 392572 146358 392624
rect 116670 392436 116676 392488
rect 116728 392476 116734 392488
rect 118694 392476 118700 392488
rect 116728 392448 118700 392476
rect 116728 392436 116734 392448
rect 118694 392436 118700 392448
rect 118752 392436 118758 392488
rect 43990 392164 43996 392216
rect 44048 392204 44054 392216
rect 88978 392204 88984 392216
rect 44048 392176 88984 392204
rect 44048 392164 44054 392176
rect 88978 392164 88984 392176
rect 89036 392164 89042 392216
rect 101030 392164 101036 392216
rect 101088 392204 101094 392216
rect 101398 392204 101404 392216
rect 101088 392176 101404 392204
rect 101088 392164 101094 392176
rect 101398 392164 101404 392176
rect 101456 392204 101462 392216
rect 135254 392204 135260 392216
rect 101456 392176 135260 392204
rect 101456 392164 101462 392176
rect 135254 392164 135260 392176
rect 135312 392164 135318 392216
rect 82906 392096 82912 392148
rect 82964 392136 82970 392148
rect 83642 392136 83648 392148
rect 82964 392108 83648 392136
rect 82964 392096 82970 392108
rect 83642 392096 83648 392108
rect 83700 392136 83706 392148
rect 140038 392136 140044 392148
rect 83700 392108 140044 392136
rect 83700 392096 83706 392108
rect 140038 392096 140044 392108
rect 140096 392096 140102 392148
rect 67358 392028 67364 392080
rect 67416 392068 67422 392080
rect 143626 392068 143632 392080
rect 67416 392040 143632 392068
rect 67416 392028 67422 392040
rect 143626 392028 143632 392040
rect 143684 392028 143690 392080
rect 52454 391960 52460 392012
rect 52512 392000 52518 392012
rect 53650 392000 53656 392012
rect 52512 391972 53656 392000
rect 52512 391960 52518 391972
rect 53650 391960 53656 391972
rect 53708 392000 53714 392012
rect 116670 392000 116676 392012
rect 53708 391972 116676 392000
rect 53708 391960 53714 391972
rect 116670 391960 116676 391972
rect 116728 391960 116734 392012
rect 120258 391960 120264 392012
rect 120316 392000 120322 392012
rect 120810 392000 120816 392012
rect 120316 391972 120816 392000
rect 120316 391960 120322 391972
rect 120810 391960 120816 391972
rect 120868 392000 120874 392012
rect 220078 392000 220084 392012
rect 120868 391972 220084 392000
rect 120868 391960 120874 391972
rect 220078 391960 220084 391972
rect 220136 391960 220142 392012
rect 41230 391892 41236 391944
rect 41288 391932 41294 391944
rect 82906 391932 82912 391944
rect 41288 391904 82912 391932
rect 41288 391892 41294 391904
rect 82906 391892 82912 391904
rect 82964 391892 82970 391944
rect 59078 391824 59084 391876
rect 59136 391864 59142 391876
rect 67358 391864 67364 391876
rect 59136 391836 67364 391864
rect 59136 391824 59142 391836
rect 67358 391824 67364 391836
rect 67416 391824 67422 391876
rect 53558 391212 53564 391264
rect 53616 391252 53622 391264
rect 75454 391252 75460 391264
rect 53616 391224 75460 391252
rect 53616 391212 53622 391224
rect 75454 391212 75460 391224
rect 75512 391212 75518 391264
rect 88978 391212 88984 391264
rect 89036 391252 89042 391264
rect 103606 391252 103612 391264
rect 89036 391224 103612 391252
rect 89036 391212 89042 391224
rect 103606 391212 103612 391224
rect 103664 391212 103670 391264
rect 110322 391212 110328 391264
rect 110380 391252 110386 391264
rect 134058 391252 134064 391264
rect 110380 391224 134064 391252
rect 110380 391212 110386 391224
rect 134058 391212 134064 391224
rect 134116 391252 134122 391264
rect 140774 391252 140780 391264
rect 134116 391224 140780 391252
rect 134116 391212 134122 391224
rect 140774 391212 140780 391224
rect 140832 391212 140838 391264
rect 50982 390668 50988 390720
rect 51040 390708 51046 390720
rect 79318 390708 79324 390720
rect 51040 390680 79324 390708
rect 51040 390668 51046 390680
rect 79318 390668 79324 390680
rect 79376 390668 79382 390720
rect 114094 390668 114100 390720
rect 114152 390708 114158 390720
rect 133138 390708 133144 390720
rect 114152 390680 133144 390708
rect 114152 390668 114158 390680
rect 133138 390668 133144 390680
rect 133196 390668 133202 390720
rect 75454 390600 75460 390652
rect 75512 390640 75518 390652
rect 134058 390640 134064 390652
rect 75512 390612 134064 390640
rect 75512 390600 75518 390612
rect 134058 390600 134064 390612
rect 134116 390600 134122 390652
rect 324406 390572 324412 390584
rect 67560 390544 324412 390572
rect 57698 390464 57704 390516
rect 57756 390504 57762 390516
rect 67560 390504 67588 390544
rect 324406 390532 324412 390544
rect 324464 390532 324470 390584
rect 57756 390476 67588 390504
rect 57756 390464 57762 390476
rect 109770 390124 109776 390176
rect 109828 390164 109834 390176
rect 114922 390164 114928 390176
rect 109828 390136 114928 390164
rect 109828 390124 109834 390136
rect 114922 390124 114928 390136
rect 114980 390124 114986 390176
rect 103330 390056 103336 390108
rect 103388 390096 103394 390108
rect 115198 390096 115204 390108
rect 103388 390068 115204 390096
rect 103388 390056 103394 390068
rect 115198 390056 115204 390068
rect 115256 390056 115262 390108
rect 114462 389920 114468 389972
rect 114520 389960 114526 389972
rect 124306 389960 124312 389972
rect 114520 389932 124312 389960
rect 114520 389920 114526 389932
rect 124306 389920 124312 389932
rect 124364 389960 124370 389972
rect 128538 389960 128544 389972
rect 124364 389932 128544 389960
rect 124364 389920 124370 389932
rect 128538 389920 128544 389932
rect 128596 389920 128602 389972
rect 115842 389852 115848 389904
rect 115900 389892 115906 389904
rect 120166 389892 120172 389904
rect 115900 389864 120172 389892
rect 115900 389852 115906 389864
rect 120166 389852 120172 389864
rect 120224 389892 120230 389904
rect 147858 389892 147864 389904
rect 120224 389864 147864 389892
rect 120224 389852 120230 389864
rect 147858 389852 147864 389864
rect 147916 389852 147922 389904
rect 41230 389784 41236 389836
rect 41288 389824 41294 389836
rect 73338 389824 73344 389836
rect 41288 389796 73344 389824
rect 41288 389784 41294 389796
rect 73338 389784 73344 389796
rect 73396 389784 73402 389836
rect 99282 389784 99288 389836
rect 99340 389824 99346 389836
rect 128354 389824 128360 389836
rect 99340 389796 128360 389824
rect 99340 389784 99346 389796
rect 128354 389784 128360 389796
rect 128412 389784 128418 389836
rect 119430 389580 119436 389632
rect 119488 389620 119494 389632
rect 120902 389620 120908 389632
rect 119488 389592 120908 389620
rect 119488 389580 119494 389592
rect 120902 389580 120908 389592
rect 120960 389580 120966 389632
rect 71682 389308 71688 389360
rect 71740 389348 71746 389360
rect 73338 389348 73344 389360
rect 71740 389320 73344 389348
rect 71740 389308 71746 389320
rect 73338 389308 73344 389320
rect 73396 389308 73402 389360
rect 49602 389172 49608 389224
rect 49660 389212 49666 389224
rect 53834 389212 53840 389224
rect 49660 389184 53840 389212
rect 49660 389172 49666 389184
rect 53834 389172 53840 389184
rect 53892 389172 53898 389224
rect 55030 389172 55036 389224
rect 55088 389212 55094 389224
rect 95510 389212 95516 389224
rect 55088 389184 95516 389212
rect 55088 389172 55094 389184
rect 95510 389172 95516 389184
rect 95568 389172 95574 389224
rect 128354 389172 128360 389224
rect 128412 389212 128418 389224
rect 130378 389212 130384 389224
rect 128412 389184 130384 389212
rect 128412 389172 128418 389184
rect 130378 389172 130384 389184
rect 130436 389172 130442 389224
rect 103606 389104 103612 389156
rect 103664 389144 103670 389156
rect 110414 389144 110420 389156
rect 103664 389116 110420 389144
rect 103664 389104 103670 389116
rect 110414 389104 110420 389116
rect 110472 389104 110478 389156
rect 112530 388628 112536 388680
rect 112588 388668 112594 388680
rect 121546 388668 121552 388680
rect 112588 388640 121552 388668
rect 112588 388628 112594 388640
rect 121546 388628 121552 388640
rect 121604 388628 121610 388680
rect 53834 388560 53840 388612
rect 53892 388600 53898 388612
rect 77478 388600 77484 388612
rect 53892 388572 77484 388600
rect 53892 388560 53898 388572
rect 77478 388560 77484 388572
rect 77536 388560 77542 388612
rect 94866 388560 94872 388612
rect 94924 388600 94930 388612
rect 102226 388600 102232 388612
rect 94924 388572 102232 388600
rect 94924 388560 94930 388572
rect 102226 388560 102232 388572
rect 102284 388560 102290 388612
rect 104618 388560 104624 388612
rect 104676 388600 104682 388612
rect 114462 388600 114468 388612
rect 104676 388572 114468 388600
rect 104676 388560 104682 388572
rect 114462 388560 114468 388572
rect 114520 388560 114526 388612
rect 69658 388492 69664 388544
rect 69716 388532 69722 388544
rect 88886 388532 88892 388544
rect 69716 388504 88892 388532
rect 69716 388492 69722 388504
rect 88886 388492 88892 388504
rect 88944 388492 88950 388544
rect 102594 388492 102600 388544
rect 102652 388532 102658 388544
rect 115934 388532 115940 388544
rect 102652 388504 115940 388532
rect 102652 388492 102658 388504
rect 115934 388492 115940 388504
rect 115992 388532 115998 388544
rect 159450 388532 159456 388544
rect 115992 388504 159456 388532
rect 115992 388492 115998 388504
rect 159450 388492 159456 388504
rect 159508 388492 159514 388544
rect 52362 388424 52368 388476
rect 52420 388464 52426 388476
rect 77294 388464 77300 388476
rect 52420 388436 77300 388464
rect 52420 388424 52426 388436
rect 77294 388424 77300 388436
rect 77352 388424 77358 388476
rect 110414 388424 110420 388476
rect 110472 388464 110478 388476
rect 309134 388464 309140 388476
rect 110472 388436 309140 388464
rect 110472 388424 110478 388436
rect 309134 388424 309140 388436
rect 309192 388424 309198 388476
rect 95418 388124 95424 388136
rect 80026 388096 95424 388124
rect 77294 388016 77300 388068
rect 77352 388056 77358 388068
rect 78490 388056 78496 388068
rect 77352 388028 78496 388056
rect 77352 388016 77358 388028
rect 78490 388016 78496 388028
rect 78548 388056 78554 388068
rect 80026 388056 80054 388096
rect 95418 388084 95424 388096
rect 95476 388084 95482 388136
rect 78548 388028 80054 388056
rect 78548 388016 78554 388028
rect 92842 388016 92848 388068
rect 92900 388056 92906 388068
rect 95878 388056 95884 388068
rect 92900 388028 95884 388056
rect 92900 388016 92906 388028
rect 95878 388016 95884 388028
rect 95936 388016 95942 388068
rect 52270 387948 52276 388000
rect 52328 387988 52334 388000
rect 69750 387988 69756 388000
rect 52328 387960 69756 387988
rect 52328 387948 52334 387960
rect 69750 387948 69756 387960
rect 69808 387948 69814 388000
rect 81434 387948 81440 388000
rect 81492 387988 81498 388000
rect 82538 387988 82544 388000
rect 81492 387960 82544 387988
rect 81492 387948 81498 387960
rect 82538 387948 82544 387960
rect 82596 387988 82602 388000
rect 86954 387988 86960 388000
rect 82596 387960 86960 387988
rect 82596 387948 82602 387960
rect 86954 387948 86960 387960
rect 87012 387948 87018 388000
rect 93302 387948 93308 388000
rect 93360 387988 93366 388000
rect 119338 387988 119344 388000
rect 93360 387960 119344 387988
rect 93360 387948 93366 387960
rect 119338 387948 119344 387960
rect 119396 387948 119402 388000
rect 53742 387880 53748 387932
rect 53800 387920 53806 387932
rect 87046 387920 87052 387932
rect 53800 387892 87052 387920
rect 53800 387880 53806 387892
rect 87046 387880 87052 387892
rect 87104 387880 87110 387932
rect 91554 387880 91560 387932
rect 91612 387920 91618 387932
rect 108298 387920 108304 387932
rect 91612 387892 108304 387920
rect 91612 387880 91618 387892
rect 108298 387880 108304 387892
rect 108356 387880 108362 387932
rect 114922 387880 114928 387932
rect 114980 387920 114986 387932
rect 184198 387920 184204 387932
rect 114980 387892 184204 387920
rect 114980 387880 114986 387892
rect 184198 387880 184204 387892
rect 184256 387880 184262 387932
rect 4798 387812 4804 387864
rect 4856 387852 4862 387864
rect 71774 387852 71780 387864
rect 4856 387824 71780 387852
rect 4856 387812 4862 387824
rect 71774 387812 71780 387824
rect 71832 387852 71838 387864
rect 72694 387852 72700 387864
rect 71832 387824 72700 387852
rect 71832 387812 71838 387824
rect 72694 387812 72700 387824
rect 72752 387852 72758 387864
rect 119430 387852 119436 387864
rect 72752 387824 119436 387852
rect 72752 387812 72758 387824
rect 119430 387812 119436 387824
rect 119488 387812 119494 387864
rect 121546 387812 121552 387864
rect 121604 387852 121610 387864
rect 244918 387852 244924 387864
rect 121604 387824 244924 387852
rect 121604 387812 121610 387824
rect 244918 387812 244924 387824
rect 244976 387812 244982 387864
rect 57790 387744 57796 387796
rect 57848 387784 57854 387796
rect 58618 387784 58624 387796
rect 57848 387756 58624 387784
rect 57848 387744 57854 387756
rect 58618 387744 58624 387756
rect 58676 387744 58682 387796
rect 107654 387744 107660 387796
rect 107712 387784 107718 387796
rect 108482 387784 108488 387796
rect 107712 387756 108488 387784
rect 107712 387744 107718 387756
rect 108482 387744 108488 387756
rect 108540 387744 108546 387796
rect 39942 387200 39948 387252
rect 40000 387240 40006 387252
rect 57238 387240 57244 387252
rect 40000 387212 57244 387240
rect 40000 387200 40006 387212
rect 57238 387200 57244 387212
rect 57296 387200 57302 387252
rect 57790 387200 57796 387252
rect 57848 387240 57854 387252
rect 77938 387240 77944 387252
rect 57848 387212 77944 387240
rect 57848 387200 57854 387212
rect 77938 387200 77944 387212
rect 77996 387200 78002 387252
rect 52178 387132 52184 387184
rect 52236 387172 52242 387184
rect 80146 387172 80152 387184
rect 52236 387144 80152 387172
rect 52236 387132 52242 387144
rect 80146 387132 80152 387144
rect 80204 387132 80210 387184
rect 86954 387132 86960 387184
rect 87012 387172 87018 387184
rect 154574 387172 154580 387184
rect 87012 387144 154580 387172
rect 87012 387132 87018 387144
rect 154574 387132 154580 387144
rect 154632 387132 154638 387184
rect 38470 387064 38476 387116
rect 38528 387104 38534 387116
rect 110598 387104 110604 387116
rect 38528 387076 110604 387104
rect 38528 387064 38534 387076
rect 110598 387064 110604 387076
rect 110656 387104 110662 387116
rect 115934 387104 115940 387116
rect 110656 387076 115940 387104
rect 110656 387064 110662 387076
rect 115934 387064 115940 387076
rect 115992 387064 115998 387116
rect 108482 386588 108488 386640
rect 108540 386628 108546 386640
rect 123662 386628 123668 386640
rect 108540 386600 123668 386628
rect 108540 386588 108546 386600
rect 123662 386588 123668 386600
rect 123720 386588 123726 386640
rect 57238 386520 57244 386572
rect 57296 386560 57302 386572
rect 84470 386560 84476 386572
rect 57296 386532 84476 386560
rect 57296 386520 57302 386532
rect 84470 386520 84476 386532
rect 84528 386520 84534 386572
rect 112162 386520 112168 386572
rect 112220 386560 112226 386572
rect 112438 386560 112444 386572
rect 112220 386532 112444 386560
rect 112220 386520 112226 386532
rect 112438 386520 112444 386532
rect 112496 386560 112502 386572
rect 167638 386560 167644 386572
rect 112496 386532 167644 386560
rect 112496 386520 112502 386532
rect 167638 386520 167644 386532
rect 167696 386520 167702 386572
rect 48222 386452 48228 386504
rect 48280 386492 48286 386504
rect 80606 386492 80612 386504
rect 48280 386464 80612 386492
rect 48280 386452 48286 386464
rect 80606 386452 80612 386464
rect 80664 386452 80670 386504
rect 107194 386452 107200 386504
rect 107252 386492 107258 386504
rect 127066 386492 127072 386504
rect 107252 386464 127072 386492
rect 107252 386452 107258 386464
rect 127066 386452 127072 386464
rect 127124 386452 127130 386504
rect 154574 386452 154580 386504
rect 154632 386492 154638 386504
rect 321554 386492 321560 386504
rect 154632 386464 321560 386492
rect 154632 386452 154638 386464
rect 321554 386452 321560 386464
rect 321612 386452 321618 386504
rect 323578 386424 323584 386436
rect 60016 386396 323584 386424
rect 60016 386368 60044 386396
rect 323578 386384 323584 386396
rect 323636 386384 323642 386436
rect 58986 386316 58992 386368
rect 59044 386356 59050 386368
rect 59998 386356 60004 386368
rect 59044 386328 60004 386356
rect 59044 386316 59050 386328
rect 59998 386316 60004 386328
rect 60056 386316 60062 386368
rect 76006 386152 76012 386164
rect 64846 386124 76012 386152
rect 54846 385704 54852 385756
rect 54904 385744 54910 385756
rect 64846 385744 64874 386124
rect 76006 386112 76012 386124
rect 76064 386112 76070 386164
rect 106090 386044 106096 386096
rect 106148 386084 106154 386096
rect 106148 386056 106228 386084
rect 106148 386044 106154 386056
rect 84286 386016 84292 386028
rect 54904 385716 64874 385744
rect 70366 385988 84292 386016
rect 54904 385704 54910 385716
rect 53558 385636 53564 385688
rect 53616 385676 53622 385688
rect 70366 385676 70394 385988
rect 84286 385976 84292 385988
rect 84344 385976 84350 386028
rect 106200 385744 106228 386056
rect 108298 385976 108304 386028
rect 108356 386016 108362 386028
rect 121546 386016 121552 386028
rect 108356 385988 121552 386016
rect 108356 385976 108362 385988
rect 121546 385976 121552 385988
rect 121604 385976 121610 386028
rect 134150 385744 134156 385756
rect 106200 385716 134156 385744
rect 134150 385704 134156 385716
rect 134208 385704 134214 385756
rect 53616 385648 70394 385676
rect 53616 385636 53622 385648
rect 95418 385636 95424 385688
rect 95476 385676 95482 385688
rect 128354 385676 128360 385688
rect 95476 385648 128360 385676
rect 95476 385636 95482 385648
rect 128354 385636 128360 385648
rect 128412 385636 128418 385688
rect 71774 385336 71780 385348
rect 64846 385308 71780 385336
rect 39666 385092 39672 385144
rect 39724 385132 39730 385144
rect 64846 385132 64874 385308
rect 71774 385296 71780 385308
rect 71832 385296 71838 385348
rect 92934 385336 92940 385348
rect 80026 385308 92940 385336
rect 39724 385104 64874 385132
rect 39724 385092 39730 385104
rect 48130 385024 48136 385076
rect 48188 385064 48194 385076
rect 53742 385064 53748 385076
rect 48188 385036 53748 385064
rect 48188 385024 48194 385036
rect 53742 385024 53748 385036
rect 53800 385064 53806 385076
rect 80026 385064 80054 385308
rect 92934 385296 92940 385308
rect 92992 385296 92998 385348
rect 104434 385296 104440 385348
rect 104492 385336 104498 385348
rect 104492 385308 113174 385336
rect 104492 385296 104498 385308
rect 53800 385036 80054 385064
rect 113146 385064 113174 385308
rect 121546 385092 121552 385144
rect 121604 385132 121610 385144
rect 263594 385132 263600 385144
rect 121604 385104 263600 385132
rect 121604 385092 121610 385104
rect 263594 385092 263600 385104
rect 263652 385092 263658 385144
rect 122650 385064 122656 385076
rect 113146 385036 122656 385064
rect 53800 385024 53806 385036
rect 122650 385024 122656 385036
rect 122708 385064 122714 385076
rect 122708 385036 122834 385064
rect 122708 385024 122714 385036
rect 61746 384956 61752 385008
rect 61804 384996 61810 385008
rect 67634 384996 67640 385008
rect 61804 384968 67640 384996
rect 61804 384956 61810 384968
rect 67634 384956 67640 384968
rect 67692 384956 67698 385008
rect 122806 384996 122834 385036
rect 128354 385024 128360 385076
rect 128412 385064 128418 385076
rect 301498 385064 301504 385076
rect 128412 385036 301504 385064
rect 128412 385024 128418 385036
rect 301498 385024 301504 385036
rect 301556 385024 301562 385076
rect 132494 384996 132500 385008
rect 122806 384968 132500 384996
rect 132494 384956 132500 384968
rect 132552 384956 132558 385008
rect 118510 384752 118516 384804
rect 118568 384792 118574 384804
rect 124306 384792 124312 384804
rect 118568 384764 124312 384792
rect 118568 384752 118574 384764
rect 124306 384752 124312 384764
rect 124364 384752 124370 384804
rect 60642 384480 60648 384532
rect 60700 384520 60706 384532
rect 61746 384520 61752 384532
rect 60700 384492 61752 384520
rect 60700 384480 60706 384492
rect 61746 384480 61752 384492
rect 61804 384480 61810 384532
rect 118602 384344 118608 384396
rect 118660 384384 118666 384396
rect 124122 384384 124128 384396
rect 118660 384356 124128 384384
rect 118660 384344 118666 384356
rect 124122 384344 124128 384356
rect 124180 384384 124186 384396
rect 127158 384384 127164 384396
rect 124180 384356 127164 384384
rect 124180 384344 124186 384356
rect 127158 384344 127164 384356
rect 127216 384344 127222 384396
rect 39942 383664 39948 383716
rect 40000 383704 40006 383716
rect 68738 383704 68744 383716
rect 40000 383676 68744 383704
rect 40000 383664 40006 383676
rect 68738 383664 68744 383676
rect 68796 383664 68802 383716
rect 126882 383120 126888 383172
rect 126940 383160 126946 383172
rect 147766 383160 147772 383172
rect 126940 383132 147772 383160
rect 126940 383120 126946 383132
rect 147766 383120 147772 383132
rect 147824 383120 147830 383172
rect 118602 383052 118608 383104
rect 118660 383092 118666 383104
rect 125502 383092 125508 383104
rect 118660 383064 125508 383092
rect 118660 383052 118666 383064
rect 125502 383052 125508 383064
rect 125560 383052 125566 383104
rect 119430 382984 119436 383036
rect 119488 383024 119494 383036
rect 147766 383024 147772 383036
rect 119488 382996 147772 383024
rect 119488 382984 119494 382996
rect 147766 382984 147772 382996
rect 147824 382984 147830 383036
rect 124306 382916 124312 382968
rect 124364 382956 124370 382968
rect 349798 382956 349804 382968
rect 124364 382928 349804 382956
rect 124364 382916 124370 382928
rect 349798 382916 349804 382928
rect 349856 382916 349862 382968
rect 125502 382644 125508 382696
rect 125560 382684 125566 382696
rect 126974 382684 126980 382696
rect 125560 382656 126980 382684
rect 125560 382644 125566 382656
rect 126974 382644 126980 382656
rect 127032 382644 127038 382696
rect 42702 382236 42708 382288
rect 42760 382276 42766 382288
rect 67634 382276 67640 382288
rect 42760 382248 67640 382276
rect 42760 382236 42766 382248
rect 67634 382236 67640 382248
rect 67692 382236 67698 382288
rect 147766 382236 147772 382288
rect 147824 382276 147830 382288
rect 209774 382276 209780 382288
rect 147824 382248 209780 382276
rect 147824 382236 147830 382248
rect 209774 382236 209780 382248
rect 209832 382236 209838 382288
rect 118602 382168 118608 382220
rect 118660 382208 118666 382220
rect 152090 382208 152096 382220
rect 118660 382180 152096 382208
rect 118660 382168 118666 382180
rect 152090 382168 152096 382180
rect 152148 382208 152154 382220
rect 153102 382208 153108 382220
rect 152148 382180 153108 382208
rect 152148 382168 152154 382180
rect 153102 382168 153108 382180
rect 153160 382168 153166 382220
rect 118602 381556 118608 381608
rect 118660 381596 118666 381608
rect 126238 381596 126244 381608
rect 118660 381568 126244 381596
rect 118660 381556 118666 381568
rect 126238 381556 126244 381568
rect 126296 381596 126302 381608
rect 126882 381596 126888 381608
rect 126296 381568 126888 381596
rect 126296 381556 126302 381568
rect 126882 381556 126888 381568
rect 126940 381556 126946 381608
rect 116394 381488 116400 381540
rect 116452 381528 116458 381540
rect 125594 381528 125600 381540
rect 116452 381500 125600 381528
rect 116452 381488 116458 381500
rect 125594 381488 125600 381500
rect 125652 381528 125658 381540
rect 137278 381528 137284 381540
rect 125652 381500 137284 381528
rect 125652 381488 125658 381500
rect 137278 381488 137284 381500
rect 137336 381488 137342 381540
rect 153102 381488 153108 381540
rect 153160 381528 153166 381540
rect 181438 381528 181444 381540
rect 153160 381500 181444 381528
rect 153160 381488 153166 381500
rect 181438 381488 181444 381500
rect 181496 381488 181502 381540
rect 42794 380128 42800 380180
rect 42852 380168 42858 380180
rect 43898 380168 43904 380180
rect 42852 380140 43904 380168
rect 42852 380128 42858 380140
rect 43898 380128 43904 380140
rect 43956 380168 43962 380180
rect 67910 380168 67916 380180
rect 43956 380140 67916 380168
rect 43956 380128 43962 380140
rect 67910 380128 67916 380140
rect 67968 380128 67974 380180
rect 118326 380128 118332 380180
rect 118384 380168 118390 380180
rect 189718 380168 189724 380180
rect 118384 380140 189724 380168
rect 118384 380128 118390 380140
rect 189718 380128 189724 380140
rect 189776 380128 189782 380180
rect 3418 378768 3424 378820
rect 3476 378808 3482 378820
rect 42794 378808 42800 378820
rect 3476 378780 42800 378808
rect 3476 378768 3482 378780
rect 42794 378768 42800 378780
rect 42852 378768 42858 378820
rect 130378 378768 130384 378820
rect 130436 378808 130442 378820
rect 163498 378808 163504 378820
rect 130436 378780 163504 378808
rect 130436 378768 130442 378780
rect 163498 378768 163504 378780
rect 163556 378768 163562 378820
rect 118602 378700 118608 378752
rect 118660 378740 118666 378752
rect 124122 378740 124128 378752
rect 118660 378712 124128 378740
rect 118660 378700 118666 378712
rect 124122 378700 124128 378712
rect 124180 378700 124186 378752
rect 118050 378156 118056 378208
rect 118108 378196 118114 378208
rect 129826 378196 129832 378208
rect 118108 378168 129832 378196
rect 118108 378156 118114 378168
rect 129826 378156 129832 378168
rect 129884 378156 129890 378208
rect 213178 378156 213184 378208
rect 213236 378196 213242 378208
rect 346394 378196 346400 378208
rect 213236 378168 346400 378196
rect 213236 378156 213242 378168
rect 346394 378156 346400 378168
rect 346452 378156 346458 378208
rect 353938 378156 353944 378208
rect 353996 378196 354002 378208
rect 580166 378196 580172 378208
rect 353996 378168 580172 378196
rect 353996 378156 354002 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 118234 378088 118240 378140
rect 118292 378128 118298 378140
rect 140958 378128 140964 378140
rect 118292 378100 140964 378128
rect 118292 378088 118298 378100
rect 140958 378088 140964 378100
rect 141016 378128 141022 378140
rect 141234 378128 141240 378140
rect 141016 378100 141240 378128
rect 141016 378088 141022 378100
rect 141234 378088 141240 378100
rect 141292 378088 141298 378140
rect 141234 377408 141240 377460
rect 141292 377448 141298 377460
rect 155954 377448 155960 377460
rect 141292 377420 155960 377448
rect 141292 377408 141298 377420
rect 155954 377408 155960 377420
rect 156012 377408 156018 377460
rect 171778 376864 171784 376916
rect 171836 376904 171842 376916
rect 305638 376904 305644 376916
rect 171836 376876 305644 376904
rect 171836 376864 171842 376876
rect 305638 376864 305644 376876
rect 305696 376864 305702 376916
rect 155954 376796 155960 376848
rect 156012 376836 156018 376848
rect 313274 376836 313280 376848
rect 156012 376808 313280 376836
rect 156012 376796 156018 376808
rect 313274 376796 313280 376808
rect 313332 376796 313338 376848
rect 65518 376768 65524 376780
rect 64846 376740 65524 376768
rect 34330 376660 34336 376712
rect 34388 376700 34394 376712
rect 64846 376700 64874 376740
rect 65518 376728 65524 376740
rect 65576 376768 65582 376780
rect 67634 376768 67640 376780
rect 65576 376740 67640 376768
rect 65576 376728 65582 376740
rect 67634 376728 67640 376740
rect 67692 376728 67698 376780
rect 263594 376728 263600 376780
rect 263652 376768 263658 376780
rect 520918 376768 520924 376780
rect 263652 376740 520924 376768
rect 263652 376728 263658 376740
rect 520918 376728 520924 376740
rect 520976 376728 520982 376780
rect 34388 376672 64874 376700
rect 34388 376660 34394 376672
rect 66162 376660 66168 376712
rect 66220 376700 66226 376712
rect 67726 376700 67732 376712
rect 66220 376672 67732 376700
rect 66220 376660 66226 376672
rect 67726 376660 67732 376672
rect 67784 376660 67790 376712
rect 118142 376660 118148 376712
rect 118200 376700 118206 376712
rect 143534 376700 143540 376712
rect 118200 376672 143540 376700
rect 118200 376660 118206 376672
rect 143534 376660 143540 376672
rect 143592 376700 143598 376712
rect 149054 376700 149060 376712
rect 143592 376672 149060 376700
rect 143592 376660 143598 376672
rect 149054 376660 149060 376672
rect 149112 376660 149118 376712
rect 119338 376048 119344 376100
rect 119396 376088 119402 376100
rect 297358 376088 297364 376100
rect 119396 376060 297364 376088
rect 119396 376048 119402 376060
rect 297358 376048 297364 376060
rect 297416 376048 297422 376100
rect 313274 376048 313280 376100
rect 313332 376088 313338 376100
rect 318794 376088 318800 376100
rect 313332 376060 318800 376088
rect 313332 376048 313338 376060
rect 318794 376048 318800 376060
rect 318852 376048 318858 376100
rect 133782 375980 133788 376032
rect 133840 376020 133846 376032
rect 143718 376020 143724 376032
rect 133840 375992 143724 376020
rect 133840 375980 133846 375992
rect 143718 375980 143724 375992
rect 143776 376020 143782 376032
rect 331214 376020 331220 376032
rect 143776 375992 331220 376020
rect 143776 375980 143782 375992
rect 331214 375980 331220 375992
rect 331272 375980 331278 376032
rect 233878 375436 233884 375488
rect 233936 375476 233942 375488
rect 347774 375476 347780 375488
rect 233936 375448 347780 375476
rect 233936 375436 233942 375448
rect 347774 375436 347780 375448
rect 347832 375436 347838 375488
rect 62022 375368 62028 375420
rect 62080 375408 62086 375420
rect 67082 375408 67088 375420
rect 62080 375380 67088 375408
rect 62080 375368 62086 375380
rect 67082 375368 67088 375380
rect 67140 375408 67146 375420
rect 67634 375408 67640 375420
rect 67140 375380 67640 375408
rect 67140 375368 67146 375380
rect 67634 375368 67640 375380
rect 67692 375368 67698 375420
rect 118602 375368 118608 375420
rect 118660 375408 118666 375420
rect 132586 375408 132592 375420
rect 118660 375380 132592 375408
rect 118660 375368 118666 375380
rect 132586 375368 132592 375380
rect 132644 375408 132650 375420
rect 133782 375408 133788 375420
rect 132644 375380 133788 375408
rect 132644 375368 132650 375380
rect 133782 375368 133788 375380
rect 133840 375368 133846 375420
rect 217962 375368 217968 375420
rect 218020 375408 218026 375420
rect 339494 375408 339500 375420
rect 218020 375380 339500 375408
rect 218020 375368 218026 375380
rect 339494 375368 339500 375380
rect 339552 375368 339558 375420
rect 138658 375300 138664 375352
rect 138716 375340 138722 375352
rect 141142 375340 141148 375352
rect 138716 375312 141148 375340
rect 138716 375300 138722 375312
rect 141142 375300 141148 375312
rect 141200 375300 141206 375352
rect 63310 374620 63316 374672
rect 63368 374660 63374 374672
rect 67634 374660 67640 374672
rect 63368 374632 67640 374660
rect 63368 374620 63374 374632
rect 67634 374620 67640 374632
rect 67692 374620 67698 374672
rect 129826 374620 129832 374672
rect 129884 374660 129890 374672
rect 265618 374660 265624 374672
rect 129884 374632 265624 374660
rect 129884 374620 129890 374632
rect 265618 374620 265624 374632
rect 265676 374620 265682 374672
rect 253198 374144 253204 374196
rect 253256 374184 253262 374196
rect 357434 374184 357440 374196
rect 253256 374156 357440 374184
rect 253256 374144 253262 374156
rect 357434 374144 357440 374156
rect 357492 374144 357498 374196
rect 141142 374076 141148 374128
rect 141200 374116 141206 374128
rect 327258 374116 327264 374128
rect 141200 374088 327264 374116
rect 141200 374076 141206 374088
rect 327258 374076 327264 374088
rect 327316 374076 327322 374128
rect 209774 374008 209780 374060
rect 209832 374048 209838 374060
rect 471974 374048 471980 374060
rect 209832 374020 471980 374048
rect 209832 374008 209838 374020
rect 471974 374008 471980 374020
rect 472032 374008 472038 374060
rect 60458 373940 60464 373992
rect 60516 373980 60522 373992
rect 67726 373980 67732 373992
rect 60516 373952 67732 373980
rect 60516 373940 60522 373952
rect 67726 373940 67732 373952
rect 67784 373940 67790 373992
rect 118602 373940 118608 373992
rect 118660 373980 118666 373992
rect 140866 373980 140872 373992
rect 118660 373952 140872 373980
rect 118660 373940 118666 373952
rect 140866 373940 140872 373952
rect 140924 373940 140930 373992
rect 64782 373260 64788 373312
rect 64840 373300 64846 373312
rect 67634 373300 67640 373312
rect 64840 373272 67640 373300
rect 64840 373260 64846 373272
rect 67634 373260 67640 373272
rect 67692 373260 67698 373312
rect 140866 373260 140872 373312
rect 140924 373300 140930 373312
rect 185578 373300 185584 373312
rect 140924 373272 185584 373300
rect 140924 373260 140930 373272
rect 185578 373260 185584 373272
rect 185636 373260 185642 373312
rect 220078 372988 220084 373040
rect 220136 373028 220142 373040
rect 220722 373028 220728 373040
rect 220136 373000 220728 373028
rect 220136 372988 220142 373000
rect 220722 372988 220728 373000
rect 220780 372988 220786 373040
rect 170398 372784 170404 372836
rect 170456 372824 170462 372836
rect 327166 372824 327172 372836
rect 170456 372796 327172 372824
rect 170456 372784 170462 372796
rect 327166 372784 327172 372796
rect 327224 372784 327230 372836
rect 117866 372716 117872 372768
rect 117924 372756 117930 372768
rect 284294 372756 284300 372768
rect 117924 372728 284300 372756
rect 117924 372716 117930 372728
rect 284294 372716 284300 372728
rect 284352 372716 284358 372768
rect 220722 372648 220728 372700
rect 220780 372688 220786 372700
rect 403618 372688 403624 372700
rect 220780 372660 403624 372688
rect 220780 372648 220786 372660
rect 403618 372648 403624 372660
rect 403676 372648 403682 372700
rect 59262 372580 59268 372632
rect 59320 372620 59326 372632
rect 60458 372620 60464 372632
rect 59320 372592 60464 372620
rect 59320 372580 59326 372592
rect 60458 372580 60464 372592
rect 60516 372580 60522 372632
rect 197998 372580 198004 372632
rect 198056 372620 198062 372632
rect 411898 372620 411904 372632
rect 198056 372592 411904 372620
rect 198056 372580 198062 372592
rect 411898 372580 411904 372592
rect 411956 372580 411962 372632
rect 3510 372512 3516 372564
rect 3568 372552 3574 372564
rect 39298 372552 39304 372564
rect 3568 372524 39304 372552
rect 3568 372512 3574 372524
rect 39298 372512 39304 372524
rect 39356 372512 39362 372564
rect 123570 371968 123576 372020
rect 123628 372008 123634 372020
rect 138014 372008 138020 372020
rect 123628 371980 138020 372008
rect 123628 371968 123634 371980
rect 138014 371968 138020 371980
rect 138072 372008 138078 372020
rect 139026 372008 139032 372020
rect 138072 371980 139032 372008
rect 138072 371968 138078 371980
rect 139026 371968 139032 371980
rect 139084 371968 139090 372020
rect 115842 371900 115848 371952
rect 115900 371940 115906 371952
rect 141050 371940 141056 371952
rect 115900 371912 141056 371940
rect 115900 371900 115906 371912
rect 141050 371900 141056 371912
rect 141108 371900 141114 371952
rect 120074 371832 120080 371884
rect 120132 371872 120138 371884
rect 135438 371872 135444 371884
rect 120132 371844 135444 371872
rect 120132 371832 120138 371844
rect 135438 371832 135444 371844
rect 135496 371832 135502 371884
rect 139486 371832 139492 371884
rect 139544 371872 139550 371884
rect 339586 371872 339592 371884
rect 139544 371844 339592 371872
rect 139544 371832 139550 371844
rect 339586 371832 339592 371844
rect 339644 371832 339650 371884
rect 139026 371356 139032 371408
rect 139084 371396 139090 371408
rect 139084 371368 142154 371396
rect 139084 371356 139090 371368
rect 135898 371288 135904 371340
rect 135956 371328 135962 371340
rect 139486 371328 139492 371340
rect 135956 371300 139492 371328
rect 135956 371288 135962 371300
rect 139486 371288 139492 371300
rect 139544 371288 139550 371340
rect 142126 371328 142154 371368
rect 342254 371328 342260 371340
rect 142126 371300 342260 371328
rect 342254 371288 342260 371300
rect 342312 371288 342318 371340
rect 117774 371220 117780 371272
rect 117832 371260 117838 371272
rect 338758 371260 338764 371272
rect 117832 371232 338764 371260
rect 117832 371220 117838 371232
rect 338758 371220 338764 371232
rect 338816 371220 338822 371272
rect 54938 370472 54944 370524
rect 54996 370512 55002 370524
rect 67634 370512 67640 370524
rect 54996 370484 67640 370512
rect 54996 370472 55002 370484
rect 67634 370472 67640 370484
rect 67692 370472 67698 370524
rect 118602 370472 118608 370524
rect 118660 370512 118666 370524
rect 120166 370512 120172 370524
rect 118660 370484 120172 370512
rect 118660 370472 118666 370484
rect 120166 370472 120172 370484
rect 120224 370512 120230 370524
rect 129826 370512 129832 370524
rect 120224 370484 129832 370512
rect 120224 370472 120230 370484
rect 129826 370472 129832 370484
rect 129884 370472 129890 370524
rect 284294 370472 284300 370524
rect 284352 370512 284358 370524
rect 337378 370512 337384 370524
rect 284352 370484 337384 370512
rect 284352 370472 284358 370484
rect 337378 370472 337384 370484
rect 337436 370472 337442 370524
rect 249702 370132 249708 370184
rect 249760 370172 249766 370184
rect 324958 370172 324964 370184
rect 249760 370144 324964 370172
rect 249760 370132 249766 370144
rect 324958 370132 324964 370144
rect 325016 370132 325022 370184
rect 169110 370064 169116 370116
rect 169168 370104 169174 370116
rect 282914 370104 282920 370116
rect 169168 370076 282920 370104
rect 169168 370064 169174 370076
rect 282914 370064 282920 370076
rect 282972 370064 282978 370116
rect 174630 369996 174636 370048
rect 174688 370036 174694 370048
rect 295334 370036 295340 370048
rect 174688 370008 295340 370036
rect 174688 369996 174694 370008
rect 295334 369996 295340 370008
rect 295392 369996 295398 370048
rect 212902 369928 212908 369980
rect 212960 369968 212966 369980
rect 417418 369968 417424 369980
rect 212960 369940 417424 369968
rect 212960 369928 212966 369940
rect 417418 369928 417424 369940
rect 417476 369928 417482 369980
rect 37182 369860 37188 369912
rect 37240 369900 37246 369912
rect 37240 369872 62160 369900
rect 37240 369860 37246 369872
rect 62132 369832 62160 369872
rect 223482 369860 223488 369912
rect 223540 369900 223546 369912
rect 464338 369900 464344 369912
rect 223540 369872 464344 369900
rect 223540 369860 223546 369872
rect 464338 369860 464344 369872
rect 464396 369860 464402 369912
rect 62758 369832 62764 369844
rect 62132 369804 62764 369832
rect 62758 369792 62764 369804
rect 62816 369832 62822 369844
rect 67634 369832 67640 369844
rect 62816 369804 67640 369832
rect 62816 369792 62822 369804
rect 67634 369792 67640 369804
rect 67692 369792 67698 369844
rect 118418 369792 118424 369844
rect 118476 369832 118482 369844
rect 132494 369832 132500 369844
rect 118476 369804 132500 369832
rect 118476 369792 118482 369804
rect 132494 369792 132500 369804
rect 132552 369832 132558 369844
rect 141418 369832 141424 369844
rect 132552 369804 141424 369832
rect 132552 369792 132558 369804
rect 141418 369792 141424 369804
rect 141476 369792 141482 369844
rect 120994 369180 121000 369232
rect 121052 369220 121058 369232
rect 125870 369220 125876 369232
rect 121052 369192 125876 369220
rect 121052 369180 121058 369192
rect 125870 369180 125876 369192
rect 125928 369180 125934 369232
rect 60366 369112 60372 369164
rect 60424 369152 60430 369164
rect 69658 369152 69664 369164
rect 60424 369124 69664 369152
rect 60424 369112 60430 369124
rect 69658 369112 69664 369124
rect 69716 369112 69722 369164
rect 118694 369112 118700 369164
rect 118752 369152 118758 369164
rect 255314 369152 255320 369164
rect 118752 369124 255320 369152
rect 118752 369112 118758 369124
rect 255314 369112 255320 369124
rect 255372 369112 255378 369164
rect 258718 368772 258724 368824
rect 258776 368812 258782 368824
rect 343634 368812 343640 368824
rect 258776 368784 343640 368812
rect 258776 368772 258782 368784
rect 343634 368772 343640 368784
rect 343692 368772 343698 368824
rect 194042 368704 194048 368756
rect 194100 368744 194106 368756
rect 333974 368744 333980 368756
rect 194100 368716 333980 368744
rect 194100 368704 194106 368716
rect 333974 368704 333980 368716
rect 334032 368704 334038 368756
rect 119338 368636 119344 368688
rect 119396 368676 119402 368688
rect 270218 368676 270224 368688
rect 119396 368648 270224 368676
rect 119396 368636 119402 368648
rect 270218 368636 270224 368648
rect 270276 368636 270282 368688
rect 282914 368636 282920 368688
rect 282972 368676 282978 368688
rect 335446 368676 335452 368688
rect 282972 368648 335452 368676
rect 282972 368636 282978 368648
rect 335446 368636 335452 368648
rect 335504 368636 335510 368688
rect 160830 368568 160836 368620
rect 160888 368608 160894 368620
rect 323118 368608 323124 368620
rect 160888 368580 323124 368608
rect 160888 368568 160894 368580
rect 323118 368568 323124 368580
rect 323176 368568 323182 368620
rect 49510 368500 49516 368552
rect 49568 368540 49574 368552
rect 53650 368540 53656 368552
rect 49568 368512 53656 368540
rect 49568 368500 49574 368512
rect 53650 368500 53656 368512
rect 53708 368540 53714 368552
rect 67634 368540 67640 368552
rect 53708 368512 67640 368540
rect 53708 368500 53714 368512
rect 67634 368500 67640 368512
rect 67692 368500 67698 368552
rect 255314 368500 255320 368552
rect 255372 368540 255378 368552
rect 457438 368540 457444 368552
rect 255372 368512 457444 368540
rect 255372 368500 255378 368512
rect 457438 368500 457444 368512
rect 457496 368500 457502 368552
rect 117774 367820 117780 367872
rect 117832 367860 117838 367872
rect 120074 367860 120080 367872
rect 117832 367832 120080 367860
rect 117832 367820 117838 367832
rect 120074 367820 120080 367832
rect 120132 367820 120138 367872
rect 118602 367752 118608 367804
rect 118660 367792 118666 367804
rect 122742 367792 122748 367804
rect 118660 367764 122748 367792
rect 118660 367752 118666 367764
rect 122742 367752 122748 367764
rect 122800 367792 122806 367804
rect 126422 367792 126428 367804
rect 122800 367764 126428 367792
rect 122800 367752 122806 367764
rect 126422 367752 126428 367764
rect 126480 367752 126486 367804
rect 269850 367412 269856 367464
rect 269908 367452 269914 367464
rect 270218 367452 270224 367464
rect 269908 367424 270224 367452
rect 269908 367412 269914 367424
rect 270218 367412 270224 367424
rect 270276 367452 270282 367464
rect 340874 367452 340880 367464
rect 270276 367424 340880 367452
rect 270276 367412 270282 367424
rect 340874 367412 340880 367424
rect 340932 367412 340938 367464
rect 286318 367344 286324 367396
rect 286376 367384 286382 367396
rect 286594 367384 286600 367396
rect 286376 367356 286600 367384
rect 286376 367344 286382 367356
rect 286594 367344 286600 367356
rect 286652 367384 286658 367396
rect 371878 367384 371884 367396
rect 286652 367356 371884 367384
rect 286652 367344 286658 367356
rect 371878 367344 371884 367356
rect 371936 367344 371942 367396
rect 166258 367276 166264 367328
rect 166316 367316 166322 367328
rect 300118 367316 300124 367328
rect 166316 367288 300124 367316
rect 166316 367276 166322 367288
rect 300118 367276 300124 367288
rect 300176 367276 300182 367328
rect 182910 367208 182916 367260
rect 182968 367248 182974 367260
rect 324498 367248 324504 367260
rect 182968 367220 324504 367248
rect 182968 367208 182974 367220
rect 324498 367208 324504 367220
rect 324556 367208 324562 367260
rect 126330 367140 126336 367192
rect 126388 367180 126394 367192
rect 293218 367180 293224 367192
rect 126388 367152 293224 367180
rect 126388 367140 126394 367152
rect 293218 367140 293224 367152
rect 293276 367140 293282 367192
rect 295334 367140 295340 367192
rect 295392 367180 295398 367192
rect 295610 367180 295616 367192
rect 295392 367152 295616 367180
rect 295392 367140 295398 367152
rect 295610 367140 295616 367152
rect 295668 367180 295674 367192
rect 350534 367180 350540 367192
rect 295668 367152 350540 367180
rect 295668 367140 295674 367152
rect 350534 367140 350540 367152
rect 350592 367140 350598 367192
rect 123478 367072 123484 367124
rect 123536 367112 123542 367124
rect 321830 367112 321836 367124
rect 123536 367084 321836 367112
rect 123536 367072 123542 367084
rect 321830 367072 321836 367084
rect 321888 367072 321894 367124
rect 59078 367004 59084 367056
rect 59136 367044 59142 367056
rect 67634 367044 67640 367056
rect 59136 367016 67640 367044
rect 59136 367004 59142 367016
rect 67634 367004 67640 367016
rect 67692 367004 67698 367056
rect 118142 367004 118148 367056
rect 118200 367044 118206 367056
rect 142246 367044 142252 367056
rect 118200 367016 142252 367044
rect 118200 367004 118206 367016
rect 142246 367004 142252 367016
rect 142304 367044 142310 367056
rect 144914 367044 144920 367056
rect 142304 367016 144920 367044
rect 142304 367004 142310 367016
rect 144914 367004 144920 367016
rect 144972 367004 144978 367056
rect 189810 366052 189816 366104
rect 189868 366092 189874 366104
rect 247034 366092 247040 366104
rect 189868 366064 247040 366092
rect 189868 366052 189874 366064
rect 247034 366052 247040 366064
rect 247092 366052 247098 366104
rect 275922 366052 275928 366104
rect 275980 366092 275986 366104
rect 320174 366092 320180 366104
rect 275980 366064 320180 366092
rect 275980 366052 275986 366064
rect 320174 366052 320180 366064
rect 320232 366052 320238 366104
rect 176102 365984 176108 366036
rect 176160 366024 176166 366036
rect 209038 366024 209044 366036
rect 176160 365996 209044 366024
rect 176160 365984 176166 365996
rect 209038 365984 209044 365996
rect 209096 365984 209102 366036
rect 244918 365984 244924 366036
rect 244976 366024 244982 366036
rect 358078 366024 358084 366036
rect 244976 365996 358084 366024
rect 244976 365984 244982 365996
rect 358078 365984 358084 365996
rect 358136 365984 358142 366036
rect 162210 365916 162216 365968
rect 162268 365956 162274 365968
rect 323026 365956 323032 365968
rect 162268 365928 323032 365956
rect 162268 365916 162274 365928
rect 323026 365916 323032 365928
rect 323084 365916 323090 365968
rect 169202 365848 169208 365900
rect 169260 365888 169266 365900
rect 238662 365888 238668 365900
rect 169260 365860 238668 365888
rect 169260 365848 169266 365860
rect 238662 365848 238668 365860
rect 238720 365848 238726 365900
rect 297358 365848 297364 365900
rect 297416 365888 297422 365900
rect 475378 365888 475384 365900
rect 297416 365860 475384 365888
rect 297416 365848 297422 365860
rect 475378 365848 475384 365860
rect 475436 365848 475442 365900
rect 146938 365780 146944 365832
rect 146996 365820 147002 365832
rect 327074 365820 327080 365832
rect 146996 365792 327080 365820
rect 146996 365780 147002 365792
rect 327074 365780 327080 365792
rect 327132 365780 327138 365832
rect 124950 365712 124956 365764
rect 125008 365752 125014 365764
rect 312722 365752 312728 365764
rect 125008 365724 312728 365752
rect 125008 365712 125014 365724
rect 312722 365712 312728 365724
rect 312780 365712 312786 365764
rect 118050 365644 118056 365696
rect 118108 365684 118114 365696
rect 133874 365684 133880 365696
rect 118108 365656 133880 365684
rect 118108 365644 118114 365656
rect 133874 365644 133880 365656
rect 133932 365644 133938 365696
rect 196802 364692 196808 364744
rect 196860 364732 196866 364744
rect 216582 364732 216588 364744
rect 196860 364704 216588 364732
rect 196860 364692 196866 364704
rect 216582 364692 216588 364704
rect 216640 364692 216646 364744
rect 181530 364624 181536 364676
rect 181588 364664 181594 364676
rect 242250 364664 242256 364676
rect 181588 364636 242256 364664
rect 181588 364624 181594 364636
rect 242250 364624 242256 364636
rect 242308 364624 242314 364676
rect 309962 364624 309968 364676
rect 310020 364664 310026 364676
rect 325786 364664 325792 364676
rect 310020 364636 325792 364664
rect 310020 364624 310026 364636
rect 325786 364624 325792 364636
rect 325844 364624 325850 364676
rect 195422 364556 195428 364608
rect 195480 364596 195486 364608
rect 227714 364596 227720 364608
rect 195480 364568 227720 364596
rect 195480 364556 195486 364568
rect 227714 364556 227720 364568
rect 227772 364556 227778 364608
rect 335354 364596 335360 364608
rect 238726 364568 335360 364596
rect 171870 364488 171876 364540
rect 171928 364528 171934 364540
rect 236086 364528 236092 364540
rect 171928 364500 236092 364528
rect 171928 364488 171934 364500
rect 236086 364488 236092 364500
rect 236144 364528 236150 364540
rect 238726 364528 238754 364568
rect 335354 364556 335360 364568
rect 335412 364556 335418 364608
rect 236144 364500 238754 364528
rect 236144 364488 236150 364500
rect 257338 364488 257344 364540
rect 257396 364528 257402 364540
rect 395338 364528 395344 364540
rect 257396 364500 395344 364528
rect 257396 364488 257402 364500
rect 395338 364488 395344 364500
rect 395396 364488 395402 364540
rect 119522 364420 119528 364472
rect 119580 364460 119586 364472
rect 258718 364460 258724 364472
rect 119580 364432 258724 364460
rect 119580 364420 119586 364432
rect 258718 364420 258724 364432
rect 258776 364420 258782 364472
rect 265618 364420 265624 364472
rect 265676 364460 265682 364472
rect 414658 364460 414664 364472
rect 265676 364432 414664 364460
rect 265676 364420 265682 364432
rect 414658 364420 414664 364432
rect 414716 364420 414722 364472
rect 43898 364352 43904 364404
rect 43956 364392 43962 364404
rect 47670 364392 47676 364404
rect 43956 364364 47676 364392
rect 43956 364352 43962 364364
rect 47670 364352 47676 364364
rect 47728 364392 47734 364404
rect 47728 364364 48314 364392
rect 47728 364352 47734 364364
rect 48286 364324 48314 364364
rect 117314 364352 117320 364404
rect 117372 364392 117378 364404
rect 117372 364364 118740 364392
rect 117372 364352 117378 364364
rect 67634 364324 67640 364336
rect 48286 364296 67640 364324
rect 67634 364284 67640 364296
rect 67692 364284 67698 364336
rect 118712 364324 118740 364364
rect 148962 364352 148968 364404
rect 149020 364392 149026 364404
rect 153194 364392 153200 364404
rect 149020 364364 153200 364392
rect 149020 364352 149026 364364
rect 153194 364352 153200 364364
rect 153252 364352 153258 364404
rect 198642 364352 198648 364404
rect 198700 364392 198706 364404
rect 579614 364392 579620 364404
rect 198700 364364 579620 364392
rect 198700 364352 198706 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 148980 364324 149008 364352
rect 118712 364296 149008 364324
rect 118142 364216 118148 364268
rect 118200 364256 118206 364268
rect 139302 364256 139308 364268
rect 118200 364228 139308 364256
rect 118200 364216 118206 364228
rect 139302 364216 139308 364228
rect 139360 364216 139366 364268
rect 187050 363196 187056 363248
rect 187108 363236 187114 363248
rect 206462 363236 206468 363248
rect 187108 363208 206468 363236
rect 187108 363196 187114 363208
rect 206462 363196 206468 363208
rect 206520 363196 206526 363248
rect 305638 363196 305644 363248
rect 305696 363236 305702 363248
rect 306282 363236 306288 363248
rect 305696 363208 306288 363236
rect 305696 363196 305702 363208
rect 306282 363196 306288 363208
rect 306340 363236 306346 363248
rect 320818 363236 320824 363248
rect 306340 363208 320824 363236
rect 306340 363196 306346 363208
rect 320818 363196 320824 363208
rect 320876 363196 320882 363248
rect 191098 363128 191104 363180
rect 191156 363168 191162 363180
rect 225782 363168 225788 363180
rect 191156 363140 225788 363168
rect 191156 363128 191162 363140
rect 225782 363128 225788 363140
rect 225840 363128 225846 363180
rect 242250 363128 242256 363180
rect 242308 363168 242314 363180
rect 351914 363168 351920 363180
rect 242308 363140 351920 363168
rect 242308 363128 242314 363140
rect 351914 363128 351920 363140
rect 351972 363128 351978 363180
rect 195330 363060 195336 363112
rect 195388 363100 195394 363112
rect 321646 363100 321652 363112
rect 195388 363072 321652 363100
rect 195388 363060 195394 363072
rect 321646 363060 321652 363072
rect 321704 363060 321710 363112
rect 192478 362992 192484 363044
rect 192536 363032 192542 363044
rect 233878 363032 233884 363044
rect 192536 363004 233884 363032
rect 192536 362992 192542 363004
rect 233878 362992 233884 363004
rect 233936 362992 233942 363044
rect 268378 362992 268384 363044
rect 268436 363032 268442 363044
rect 466454 363032 466460 363044
rect 268436 363004 466460 363032
rect 268436 362992 268442 363004
rect 466454 362992 466460 363004
rect 466512 362992 466518 363044
rect 35526 362924 35532 362976
rect 35584 362964 35590 362976
rect 69198 362964 69204 362976
rect 35584 362936 69204 362964
rect 35584 362924 35590 362936
rect 69198 362924 69204 362936
rect 69256 362924 69262 362976
rect 123570 362924 123576 362976
rect 123628 362964 123634 362976
rect 213178 362964 213184 362976
rect 123628 362936 213184 362964
rect 123628 362924 123634 362936
rect 213178 362924 213184 362936
rect 213236 362924 213242 362976
rect 216582 362924 216588 362976
rect 216640 362964 216646 362976
rect 510614 362964 510620 362976
rect 216640 362936 510620 362964
rect 216640 362924 216646 362936
rect 217428 362908 217456 362936
rect 510614 362924 510620 362936
rect 510672 362924 510678 362976
rect 64690 362856 64696 362908
rect 64748 362896 64754 362908
rect 67634 362896 67640 362908
rect 64748 362868 67640 362896
rect 64748 362856 64754 362868
rect 67634 362856 67640 362868
rect 67692 362856 67698 362908
rect 117958 362856 117964 362908
rect 118016 362896 118022 362908
rect 149238 362896 149244 362908
rect 118016 362868 149244 362896
rect 118016 362856 118022 362868
rect 149238 362856 149244 362868
rect 149296 362856 149302 362908
rect 217410 362856 217416 362908
rect 217468 362856 217474 362908
rect 228358 362856 228364 362908
rect 228416 362896 228422 362908
rect 229646 362896 229652 362908
rect 228416 362868 229652 362896
rect 228416 362856 228422 362868
rect 229646 362856 229652 362868
rect 229704 362856 229710 362908
rect 316678 362448 316684 362500
rect 316736 362488 316742 362500
rect 317322 362488 317328 362500
rect 316736 362460 317328 362488
rect 316736 362448 316742 362460
rect 317322 362448 317328 362460
rect 317380 362448 317386 362500
rect 199378 362312 199384 362364
rect 199436 362352 199442 362364
rect 249702 362352 249708 362364
rect 199436 362324 249708 362352
rect 199436 362312 199442 362324
rect 249702 362312 249708 362324
rect 249760 362352 249766 362364
rect 250898 362352 250904 362364
rect 249760 362324 250904 362352
rect 249760 362312 249766 362324
rect 250898 362312 250904 362324
rect 250956 362312 250962 362364
rect 149238 362244 149244 362296
rect 149296 362284 149302 362296
rect 175918 362284 175924 362296
rect 149296 362256 175924 362284
rect 149296 362244 149302 362256
rect 175918 362244 175924 362256
rect 175976 362244 175982 362296
rect 196618 362244 196624 362296
rect 196676 362284 196682 362296
rect 275922 362284 275928 362296
rect 196676 362256 275928 362284
rect 196676 362244 196682 362256
rect 275922 362244 275928 362256
rect 275980 362284 275986 362296
rect 276658 362284 276664 362296
rect 275980 362256 276664 362284
rect 275980 362244 275986 362256
rect 276658 362244 276664 362256
rect 276716 362244 276722 362296
rect 117682 362176 117688 362228
rect 117740 362216 117746 362228
rect 144270 362216 144276 362228
rect 117740 362188 144276 362216
rect 117740 362176 117746 362188
rect 144270 362176 144276 362188
rect 144328 362176 144334 362228
rect 166350 362176 166356 362228
rect 166408 362216 166414 362228
rect 309962 362216 309968 362228
rect 166408 362188 309968 362216
rect 166408 362176 166414 362188
rect 309962 362176 309968 362188
rect 310020 362176 310026 362228
rect 213178 362108 213184 362160
rect 213236 362148 213242 362160
rect 214834 362148 214840 362160
rect 213236 362120 214840 362148
rect 213236 362108 213242 362120
rect 214834 362108 214840 362120
rect 214892 362108 214898 362160
rect 217962 362040 217968 362092
rect 218020 362080 218026 362092
rect 219342 362080 219348 362092
rect 218020 362052 219348 362080
rect 218020 362040 218026 362052
rect 219342 362040 219348 362052
rect 219400 362040 219406 362092
rect 258718 361904 258724 361956
rect 258776 361944 258782 361956
rect 259914 361944 259920 361956
rect 258776 361916 259920 361944
rect 258776 361904 258782 361916
rect 259914 361904 259920 361916
rect 259972 361904 259978 361956
rect 289170 361904 289176 361956
rect 289228 361944 289234 361956
rect 319438 361944 319444 361956
rect 289228 361916 319444 361944
rect 289228 361904 289234 361916
rect 319438 361904 319444 361916
rect 319496 361904 319502 361956
rect 281166 361836 281172 361888
rect 281224 361876 281230 361888
rect 360838 361876 360844 361888
rect 281224 361848 360844 361876
rect 281224 361836 281230 361848
rect 360838 361836 360844 361848
rect 360896 361836 360902 361888
rect 310790 361768 310796 361820
rect 310848 361808 310854 361820
rect 399478 361808 399484 361820
rect 310848 361780 399484 361808
rect 310848 361768 310854 361780
rect 399478 361768 399484 361780
rect 399536 361768 399542 361820
rect 225782 361700 225788 361752
rect 225840 361740 225846 361752
rect 317046 361740 317052 361752
rect 225840 361712 317052 361740
rect 225840 361700 225846 361712
rect 317046 361700 317052 361712
rect 317104 361700 317110 361752
rect 184842 361632 184848 361684
rect 184900 361672 184906 361684
rect 202598 361672 202604 361684
rect 184900 361644 202604 361672
rect 184900 361632 184906 361644
rect 202598 361632 202604 361644
rect 202656 361632 202662 361684
rect 249702 361632 249708 361684
rect 249760 361672 249766 361684
rect 345658 361672 345664 361684
rect 249760 361644 345664 361672
rect 249760 361632 249766 361644
rect 345658 361632 345664 361644
rect 345716 361632 345722 361684
rect 143718 361564 143724 361616
rect 143776 361604 143782 361616
rect 144270 361604 144276 361616
rect 143776 361576 144276 361604
rect 143776 361564 143782 361576
rect 144270 361564 144276 361576
rect 144328 361604 144334 361616
rect 240594 361604 240600 361616
rect 144328 361576 240600 361604
rect 144328 361564 144334 361576
rect 240594 361564 240600 361576
rect 240652 361564 240658 361616
rect 281166 361604 281172 361616
rect 252480 361576 281172 361604
rect 145098 361496 145104 361548
rect 145156 361536 145162 361548
rect 252480 361536 252508 361576
rect 281166 361564 281172 361576
rect 281224 361564 281230 361616
rect 301498 361564 301504 361616
rect 301556 361604 301562 361616
rect 410518 361604 410524 361616
rect 301556 361576 410524 361604
rect 301556 361564 301562 361576
rect 410518 361564 410524 361576
rect 410576 361564 410582 361616
rect 145156 361508 252508 361536
rect 145156 361496 145162 361508
rect 32950 360816 32956 360868
rect 33008 360856 33014 360868
rect 42794 360856 42800 360868
rect 33008 360828 42800 360856
rect 33008 360816 33014 360828
rect 42794 360816 42800 360828
rect 42852 360816 42858 360868
rect 118602 360816 118608 360868
rect 118660 360856 118666 360868
rect 121638 360856 121644 360868
rect 118660 360828 121644 360856
rect 118660 360816 118666 360828
rect 121638 360816 121644 360828
rect 121696 360856 121702 360868
rect 145098 360856 145104 360868
rect 121696 360828 145104 360856
rect 121696 360816 121702 360828
rect 145098 360816 145104 360828
rect 145156 360816 145162 360868
rect 308490 360816 308496 360868
rect 308548 360856 308554 360868
rect 309134 360856 309140 360868
rect 308548 360828 309140 360856
rect 308548 360816 308554 360828
rect 309134 360816 309140 360828
rect 309192 360856 309198 360868
rect 356698 360856 356704 360868
rect 309192 360828 356704 360856
rect 309192 360816 309198 360828
rect 356698 360816 356704 360828
rect 356756 360816 356762 360868
rect 119430 360544 119436 360596
rect 119488 360584 119494 360596
rect 314654 360584 314660 360596
rect 119488 360556 314660 360584
rect 119488 360544 119494 360556
rect 314654 360544 314660 360556
rect 314712 360544 314718 360596
rect 278130 360476 278136 360528
rect 278188 360516 278194 360528
rect 278590 360516 278596 360528
rect 278188 360488 278596 360516
rect 278188 360476 278194 360488
rect 278590 360476 278596 360488
rect 278648 360516 278654 360528
rect 352558 360516 352564 360528
rect 278648 360488 352564 360516
rect 278648 360476 278654 360488
rect 352558 360476 352564 360488
rect 352616 360476 352622 360528
rect 199470 360408 199476 360460
rect 199528 360448 199534 360460
rect 310790 360448 310796 360460
rect 199528 360420 310796 360448
rect 199528 360408 199534 360420
rect 310790 360408 310796 360420
rect 310848 360408 310854 360460
rect 196710 360340 196716 360392
rect 196768 360380 196774 360392
rect 257338 360380 257344 360392
rect 196768 360352 257344 360380
rect 196768 360340 196774 360352
rect 257338 360340 257344 360352
rect 257396 360340 257402 360392
rect 272150 360340 272156 360392
rect 272208 360380 272214 360392
rect 406378 360380 406384 360392
rect 272208 360352 406384 360380
rect 272208 360340 272214 360352
rect 406378 360340 406384 360352
rect 406436 360340 406442 360392
rect 133138 360272 133144 360324
rect 133196 360312 133202 360324
rect 324314 360312 324320 360324
rect 133196 360284 324320 360312
rect 133196 360272 133202 360284
rect 324314 360272 324320 360284
rect 324372 360272 324378 360324
rect 42794 360204 42800 360256
rect 42852 360244 42858 360256
rect 44082 360244 44088 360256
rect 42852 360216 44088 360244
rect 42852 360204 42858 360216
rect 44082 360204 44088 360216
rect 44140 360244 44146 360256
rect 67634 360244 67640 360256
rect 44140 360216 67640 360244
rect 44140 360204 44146 360216
rect 67634 360204 67640 360216
rect 67692 360204 67698 360256
rect 198826 360204 198832 360256
rect 198884 360244 198890 360256
rect 204530 360244 204536 360256
rect 198884 360216 204536 360244
rect 198884 360204 198890 360216
rect 204530 360204 204536 360216
rect 204588 360204 204594 360256
rect 312722 360204 312728 360256
rect 312780 360244 312786 360256
rect 322934 360244 322940 360256
rect 312780 360216 322940 360244
rect 312780 360204 312786 360216
rect 322934 360204 322940 360216
rect 322992 360204 322998 360256
rect 118142 360136 118148 360188
rect 118200 360176 118206 360188
rect 146478 360176 146484 360188
rect 118200 360148 146484 360176
rect 118200 360136 118206 360148
rect 146478 360136 146484 360148
rect 146536 360136 146542 360188
rect 317506 359592 317512 359644
rect 317564 359632 317570 359644
rect 319530 359632 319536 359644
rect 317564 359604 319536 359632
rect 317564 359592 317570 359604
rect 319530 359592 319536 359604
rect 319588 359592 319594 359644
rect 50890 359524 50896 359576
rect 50948 359564 50954 359576
rect 67634 359564 67640 359576
rect 50948 359536 67640 359564
rect 50948 359524 50954 359536
rect 67634 359524 67640 359536
rect 67692 359524 67698 359576
rect 36538 359456 36544 359508
rect 36596 359496 36602 359508
rect 41046 359496 41052 359508
rect 36596 359468 41052 359496
rect 36596 359456 36602 359468
rect 41046 359456 41052 359468
rect 41104 359496 41110 359508
rect 67726 359496 67732 359508
rect 41104 359468 67732 359496
rect 41104 359456 41110 359468
rect 67726 359456 67732 359468
rect 67784 359456 67790 359508
rect 118602 359456 118608 359508
rect 118660 359496 118666 359508
rect 120718 359496 120724 359508
rect 118660 359468 120724 359496
rect 118660 359456 118666 359468
rect 120718 359456 120724 359468
rect 120776 359496 120782 359508
rect 137002 359496 137008 359508
rect 120776 359468 137008 359496
rect 120776 359456 120782 359468
rect 137002 359456 137008 359468
rect 137060 359456 137066 359508
rect 205606 359468 215294 359496
rect 205606 359292 205634 359468
rect 212534 359428 212540 359440
rect 201466 359264 205634 359292
rect 212460 359400 212540 359428
rect 201466 359088 201494 359264
rect 212460 359088 212488 359400
rect 212534 359388 212540 359400
rect 212592 359388 212598 359440
rect 195946 359060 201494 359088
rect 205606 359060 212488 359088
rect 193950 358912 193956 358964
rect 194008 358952 194014 358964
rect 195946 358952 195974 359060
rect 194008 358924 195974 358952
rect 194008 358912 194014 358924
rect 199838 358912 199844 358964
rect 199896 358952 199902 358964
rect 205606 358952 205634 359060
rect 215266 359020 215294 359468
rect 314838 359388 314844 359440
rect 314896 359428 314902 359440
rect 320358 359428 320364 359440
rect 314896 359400 320364 359428
rect 314896 359388 314902 359400
rect 320358 359388 320364 359400
rect 320416 359388 320422 359440
rect 215266 358992 216674 359020
rect 199896 358924 205634 358952
rect 216646 358952 216674 358992
rect 321646 358952 321652 358964
rect 216646 358924 321652 358952
rect 199896 358912 199902 358924
rect 321646 358912 321652 358924
rect 321704 358912 321710 358964
rect 167730 358844 167736 358896
rect 167788 358884 167794 358896
rect 329834 358884 329840 358896
rect 167788 358856 195974 358884
rect 167788 358844 167794 358856
rect 195946 358816 195974 358856
rect 215266 358856 329840 358884
rect 215266 358816 215294 358856
rect 329834 358844 329840 358856
rect 329892 358844 329898 358896
rect 195946 358788 215294 358816
rect 320358 358776 320364 358828
rect 320416 358816 320422 358828
rect 495434 358816 495440 358828
rect 320416 358788 495440 358816
rect 320416 358776 320422 358788
rect 495434 358776 495440 358788
rect 495492 358776 495498 358828
rect 118050 358708 118056 358760
rect 118108 358748 118114 358760
rect 120994 358748 121000 358760
rect 118108 358720 121000 358748
rect 118108 358708 118114 358720
rect 120994 358708 121000 358720
rect 121052 358708 121058 358760
rect 125502 358708 125508 358760
rect 125560 358748 125566 358760
rect 128630 358748 128636 358760
rect 125560 358720 128636 358748
rect 125560 358708 125566 358720
rect 128630 358708 128636 358720
rect 128688 358708 128694 358760
rect 57698 358028 57704 358080
rect 57756 358068 57762 358080
rect 67634 358068 67640 358080
rect 57756 358040 67640 358068
rect 57756 358028 57762 358040
rect 67634 358028 67640 358040
rect 67692 358028 67698 358080
rect 118602 358028 118608 358080
rect 118660 358068 118666 358080
rect 122834 358068 122840 358080
rect 118660 358040 122840 358068
rect 118660 358028 118666 358040
rect 122834 358028 122840 358040
rect 122892 358068 122898 358080
rect 146938 358068 146944 358080
rect 122892 358040 146944 358068
rect 122892 358028 122898 358040
rect 146938 358028 146944 358040
rect 146996 358068 147002 358080
rect 198826 358068 198832 358080
rect 146996 358040 198832 358068
rect 146996 358028 147002 358040
rect 198826 358028 198832 358040
rect 198884 358028 198890 358080
rect 319530 358028 319536 358080
rect 319588 358068 319594 358080
rect 469214 358068 469220 358080
rect 319588 358040 469220 358068
rect 319588 358028 319594 358040
rect 469214 358028 469220 358040
rect 469272 358028 469278 358080
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 15838 357456 15844 357468
rect 3200 357428 15844 357456
rect 3200 357416 3206 357428
rect 15838 357416 15844 357428
rect 15896 357416 15902 357468
rect 128630 357416 128636 357468
rect 128688 357456 128694 357468
rect 197998 357456 198004 357468
rect 128688 357428 198004 357456
rect 128688 357416 128694 357428
rect 197998 357416 198004 357428
rect 198056 357416 198062 357468
rect 35710 357348 35716 357400
rect 35768 357388 35774 357400
rect 66898 357388 66904 357400
rect 35768 357360 66904 357388
rect 35768 357348 35774 357360
rect 66898 357348 66904 357360
rect 66956 357388 66962 357400
rect 67542 357388 67548 357400
rect 66956 357360 67548 357388
rect 66956 357348 66962 357360
rect 67542 357348 67548 357360
rect 67600 357348 67606 357400
rect 150618 357348 150624 357400
rect 150676 357388 150682 357400
rect 151906 357388 151912 357400
rect 150676 357360 151912 357388
rect 150676 357348 150682 357360
rect 151906 357348 151912 357360
rect 151964 357388 151970 357400
rect 199838 357388 199844 357400
rect 151964 357360 199844 357388
rect 151964 357348 151970 357360
rect 199838 357348 199844 357360
rect 199896 357348 199902 357400
rect 118602 356736 118608 356788
rect 118660 356776 118666 356788
rect 186958 356776 186964 356788
rect 118660 356748 186964 356776
rect 118660 356736 118666 356748
rect 186958 356736 186964 356748
rect 187016 356736 187022 356788
rect 124858 356668 124864 356720
rect 124916 356708 124922 356720
rect 198274 356708 198280 356720
rect 124916 356680 198280 356708
rect 124916 356668 124922 356680
rect 198274 356668 198280 356680
rect 198332 356708 198338 356720
rect 198642 356708 198648 356720
rect 198332 356680 198648 356708
rect 198332 356668 198338 356680
rect 198642 356668 198648 356680
rect 198700 356668 198706 356720
rect 41138 356056 41144 356108
rect 41196 356096 41202 356108
rect 68002 356096 68008 356108
rect 41196 356068 68008 356096
rect 41196 356056 41202 356068
rect 68002 356056 68008 356068
rect 68060 356056 68066 356108
rect 118602 356056 118608 356108
rect 118660 356096 118666 356108
rect 150618 356096 150624 356108
rect 118660 356068 150624 356096
rect 118660 356056 118666 356068
rect 150618 356056 150624 356068
rect 150676 356056 150682 356108
rect 118510 355988 118516 356040
rect 118568 356028 118574 356040
rect 143810 356028 143816 356040
rect 118568 356000 143816 356028
rect 118568 355988 118574 356000
rect 143810 355988 143816 356000
rect 143868 356028 143874 356040
rect 144822 356028 144828 356040
rect 143868 356000 144828 356028
rect 143868 355988 143874 356000
rect 144822 355988 144828 356000
rect 144880 355988 144886 356040
rect 56502 355376 56508 355428
rect 56560 355416 56566 355428
rect 67634 355416 67640 355428
rect 56560 355388 67640 355416
rect 56560 355376 56566 355388
rect 67634 355376 67640 355388
rect 67692 355376 67698 355428
rect 55950 355308 55956 355360
rect 56008 355348 56014 355360
rect 67726 355348 67732 355360
rect 56008 355320 67732 355348
rect 56008 355308 56014 355320
rect 67726 355308 67732 355320
rect 67784 355308 67790 355360
rect 144822 355308 144828 355360
rect 144880 355348 144886 355360
rect 182818 355348 182824 355360
rect 144880 355320 182824 355348
rect 144880 355308 144886 355320
rect 182818 355308 182824 355320
rect 182876 355308 182882 355360
rect 319898 355308 319904 355360
rect 319956 355348 319962 355360
rect 458174 355348 458180 355360
rect 319956 355320 458180 355348
rect 319956 355308 319962 355320
rect 458174 355308 458180 355320
rect 458232 355308 458238 355360
rect 135162 354628 135168 354680
rect 135220 354668 135226 354680
rect 146386 354668 146392 354680
rect 135220 354640 146392 354668
rect 135220 354628 135226 354640
rect 146386 354628 146392 354640
rect 146444 354668 146450 354680
rect 198182 354668 198188 354680
rect 146444 354640 198188 354668
rect 146444 354628 146450 354640
rect 198182 354628 198188 354640
rect 198240 354628 198246 354680
rect 118602 354356 118608 354408
rect 118660 354396 118666 354408
rect 121454 354396 121460 354408
rect 118660 354368 121460 354396
rect 118660 354356 118666 354368
rect 121454 354356 121460 354368
rect 121512 354356 121518 354408
rect 322842 354356 322848 354408
rect 322900 354396 322906 354408
rect 324498 354396 324504 354408
rect 322900 354368 324504 354396
rect 322900 354356 322906 354368
rect 324498 354356 324504 354368
rect 324556 354356 324562 354408
rect 117774 354016 117780 354068
rect 117832 354056 117838 354068
rect 133874 354056 133880 354068
rect 117832 354028 133880 354056
rect 117832 354016 117838 354028
rect 133874 354016 133880 354028
rect 133932 354056 133938 354068
rect 135162 354056 135168 354068
rect 133932 354028 135168 354056
rect 133932 354016 133938 354028
rect 135162 354016 135168 354028
rect 135220 354016 135226 354068
rect 121454 353948 121460 354000
rect 121512 353988 121518 354000
rect 142246 353988 142252 354000
rect 121512 353960 142252 353988
rect 121512 353948 121518 353960
rect 142246 353948 142252 353960
rect 142304 353988 142310 354000
rect 196802 353988 196808 354000
rect 142304 353960 196808 353988
rect 142304 353948 142310 353960
rect 196802 353948 196808 353960
rect 196860 353948 196866 354000
rect 508498 353948 508504 354000
rect 508556 353988 508562 354000
rect 579614 353988 579620 354000
rect 508556 353960 579620 353988
rect 508556 353948 508562 353960
rect 579614 353948 579620 353960
rect 579672 353948 579678 354000
rect 59998 353200 60004 353252
rect 60056 353240 60062 353252
rect 66990 353240 66996 353252
rect 60056 353212 66996 353240
rect 60056 353200 60062 353212
rect 66990 353200 66996 353212
rect 67048 353240 67054 353252
rect 67542 353240 67548 353252
rect 67048 353212 67548 353240
rect 67048 353200 67054 353212
rect 67542 353200 67548 353212
rect 67600 353200 67606 353252
rect 41414 352520 41420 352572
rect 41472 352560 41478 352572
rect 42610 352560 42616 352572
rect 41472 352532 42616 352560
rect 41472 352520 41478 352532
rect 42610 352520 42616 352532
rect 42668 352560 42674 352572
rect 68922 352560 68928 352572
rect 42668 352532 68928 352560
rect 42668 352520 42674 352532
rect 68922 352520 68928 352532
rect 68980 352520 68986 352572
rect 126422 352520 126428 352572
rect 126480 352560 126486 352572
rect 140130 352560 140136 352572
rect 126480 352532 140136 352560
rect 126480 352520 126486 352532
rect 140130 352520 140136 352532
rect 140188 352520 140194 352572
rect 21358 351908 21364 351960
rect 21416 351948 21422 351960
rect 41414 351948 41420 351960
rect 21416 351920 41420 351948
rect 21416 351908 21422 351920
rect 41414 351908 41420 351920
rect 41472 351908 41478 351960
rect 61654 351840 61660 351892
rect 61712 351880 61718 351892
rect 64138 351880 64144 351892
rect 61712 351852 64144 351880
rect 61712 351840 61718 351852
rect 64138 351840 64144 351852
rect 64196 351880 64202 351892
rect 67634 351880 67640 351892
rect 64196 351852 67640 351880
rect 64196 351840 64202 351852
rect 67634 351840 67640 351852
rect 67692 351840 67698 351892
rect 117406 351840 117412 351892
rect 117464 351880 117470 351892
rect 147674 351880 147680 351892
rect 117464 351852 147680 351880
rect 117464 351840 117470 351852
rect 147674 351840 147680 351852
rect 147732 351840 147738 351892
rect 118602 351772 118608 351824
rect 118660 351812 118666 351824
rect 145190 351812 145196 351824
rect 118660 351784 145196 351812
rect 118660 351772 118666 351784
rect 145190 351772 145196 351784
rect 145248 351772 145254 351824
rect 147674 351160 147680 351212
rect 147732 351200 147738 351212
rect 178678 351200 178684 351212
rect 147732 351172 178684 351200
rect 147732 351160 147738 351172
rect 178678 351160 178684 351172
rect 178736 351160 178742 351212
rect 319438 351160 319444 351212
rect 319496 351200 319502 351212
rect 452654 351200 452660 351212
rect 319496 351172 452660 351200
rect 319496 351160 319502 351172
rect 452654 351160 452660 351172
rect 452712 351160 452718 351212
rect 120902 350588 120908 350600
rect 120092 350560 120908 350588
rect 118602 350480 118608 350532
rect 118660 350520 118666 350532
rect 120092 350520 120120 350560
rect 120902 350548 120908 350560
rect 120960 350588 120966 350600
rect 132770 350588 132776 350600
rect 120960 350560 132776 350588
rect 120960 350548 120966 350560
rect 132770 350548 132776 350560
rect 132828 350548 132834 350600
rect 141418 350548 141424 350600
rect 141476 350588 141482 350600
rect 142430 350588 142436 350600
rect 141476 350560 142436 350588
rect 141476 350548 141482 350560
rect 142430 350548 142436 350560
rect 142488 350588 142494 350600
rect 197354 350588 197360 350600
rect 142488 350560 197360 350588
rect 142488 350548 142494 350560
rect 197354 350548 197360 350560
rect 197412 350548 197418 350600
rect 118660 350492 120120 350520
rect 118660 350480 118666 350492
rect 322658 349800 322664 349852
rect 322716 349840 322722 349852
rect 323118 349840 323124 349852
rect 322716 349812 323124 349840
rect 322716 349800 322722 349812
rect 323118 349800 323124 349812
rect 323176 349840 323182 349852
rect 489178 349840 489184 349852
rect 323176 349812 489184 349840
rect 323176 349800 323182 349812
rect 489178 349800 489184 349812
rect 489236 349800 489242 349852
rect 61930 349120 61936 349172
rect 61988 349160 61994 349172
rect 64690 349160 64696 349172
rect 61988 349132 64696 349160
rect 61988 349120 61994 349132
rect 64690 349120 64696 349132
rect 64748 349160 64754 349172
rect 67634 349160 67640 349172
rect 64748 349132 67640 349160
rect 64748 349120 64754 349132
rect 67634 349120 67640 349132
rect 67692 349120 67698 349172
rect 35618 349052 35624 349104
rect 35676 349092 35682 349104
rect 69658 349092 69664 349104
rect 35676 349064 69664 349092
rect 35676 349052 35682 349064
rect 69658 349052 69664 349064
rect 69716 349052 69722 349104
rect 118602 349052 118608 349104
rect 118660 349092 118666 349104
rect 145006 349092 145012 349104
rect 118660 349064 145012 349092
rect 118660 349052 118666 349064
rect 145006 349052 145012 349064
rect 145064 349092 145070 349104
rect 146202 349092 146208 349104
rect 145064 349064 146208 349092
rect 145064 349052 145070 349064
rect 146202 349052 146208 349064
rect 146260 349052 146266 349104
rect 63126 348984 63132 349036
rect 63184 349024 63190 349036
rect 65610 349024 65616 349036
rect 63184 348996 65616 349024
rect 63184 348984 63190 348996
rect 65610 348984 65616 348996
rect 65668 349024 65674 349036
rect 67634 349024 67640 349036
rect 65668 348996 67640 349024
rect 65668 348984 65674 348996
rect 67634 348984 67640 348996
rect 67692 348984 67698 349036
rect 118510 348984 118516 349036
rect 118568 349024 118574 349036
rect 142338 349024 142344 349036
rect 118568 348996 142344 349024
rect 118568 348984 118574 348996
rect 142338 348984 142344 348996
rect 142396 349024 142402 349036
rect 143442 349024 143448 349036
rect 142396 348996 143448 349024
rect 142396 348984 142402 348996
rect 143442 348984 143448 348996
rect 143500 348984 143506 349036
rect 322198 348372 322204 348424
rect 322256 348412 322262 348424
rect 334618 348412 334624 348424
rect 322256 348384 334624 348412
rect 322256 348372 322262 348384
rect 334618 348372 334624 348384
rect 334676 348372 334682 348424
rect 63218 347692 63224 347744
rect 63276 347732 63282 347744
rect 66162 347732 66168 347744
rect 63276 347704 66168 347732
rect 63276 347692 63282 347704
rect 66162 347692 66168 347704
rect 66220 347732 66226 347744
rect 67634 347732 67640 347744
rect 66220 347704 67640 347732
rect 66220 347692 66226 347704
rect 67634 347692 67640 347704
rect 67692 347692 67698 347744
rect 118602 347012 118608 347064
rect 118660 347052 118666 347064
rect 132586 347052 132592 347064
rect 118660 347024 132592 347052
rect 118660 347012 118666 347024
rect 132586 347012 132592 347024
rect 132644 347052 132650 347064
rect 133782 347052 133788 347064
rect 132644 347024 133788 347052
rect 132644 347012 132650 347024
rect 133782 347012 133788 347024
rect 133840 347012 133846 347064
rect 322290 347012 322296 347064
rect 322348 347052 322354 347064
rect 356054 347052 356060 347064
rect 322348 347024 356060 347052
rect 322348 347012 322354 347024
rect 356054 347012 356060 347024
rect 356112 347012 356118 347064
rect 133782 346468 133788 346520
rect 133840 346508 133846 346520
rect 180058 346508 180064 346520
rect 133840 346480 180064 346508
rect 133840 346468 133846 346480
rect 180058 346468 180064 346480
rect 180116 346468 180122 346520
rect 179322 346400 179328 346452
rect 179380 346440 179386 346452
rect 197354 346440 197360 346452
rect 179380 346412 197360 346440
rect 179380 346400 179386 346412
rect 197354 346400 197360 346412
rect 197412 346400 197418 346452
rect 15838 346332 15844 346384
rect 15896 346372 15902 346384
rect 68830 346372 68836 346384
rect 15896 346344 68836 346372
rect 15896 346332 15902 346344
rect 68830 346332 68836 346344
rect 68888 346332 68894 346384
rect 116578 346332 116584 346384
rect 116636 346372 116642 346384
rect 117314 346372 117320 346384
rect 116636 346344 117320 346372
rect 116636 346332 116642 346344
rect 117314 346332 117320 346344
rect 117372 346332 117378 346384
rect 118602 346332 118608 346384
rect 118660 346372 118666 346384
rect 136910 346372 136916 346384
rect 118660 346344 136916 346372
rect 118660 346332 118666 346344
rect 136910 346332 136916 346344
rect 136968 346372 136974 346384
rect 137186 346372 137192 346384
rect 136968 346344 137192 346372
rect 136968 346332 136974 346344
rect 137186 346332 137192 346344
rect 137244 346332 137250 346384
rect 2774 346264 2780 346316
rect 2832 346304 2838 346316
rect 4798 346304 4804 346316
rect 2832 346276 4804 346304
rect 2832 346264 2838 346276
rect 4798 346264 4804 346276
rect 4856 346264 4862 346316
rect 137186 345652 137192 345704
rect 137244 345692 137250 345704
rect 180150 345692 180156 345704
rect 137244 345664 180156 345692
rect 137244 345652 137250 345664
rect 180150 345652 180156 345664
rect 180208 345652 180214 345704
rect 45278 345040 45284 345092
rect 45336 345080 45342 345092
rect 68646 345080 68652 345092
rect 45336 345052 68652 345080
rect 45336 345040 45342 345052
rect 68646 345040 68652 345052
rect 68704 345040 68710 345092
rect 118510 345040 118516 345092
rect 118568 345080 118574 345092
rect 140866 345080 140872 345092
rect 118568 345052 140872 345080
rect 118568 345040 118574 345052
rect 140866 345040 140872 345052
rect 140924 345040 140930 345092
rect 320266 345040 320272 345092
rect 320324 345080 320330 345092
rect 461578 345080 461584 345092
rect 320324 345052 461584 345080
rect 320324 345040 320330 345052
rect 461578 345040 461584 345052
rect 461636 345040 461642 345092
rect 118602 344972 118608 345024
rect 118660 345012 118666 345024
rect 150434 345012 150440 345024
rect 118660 344984 150440 345012
rect 118660 344972 118666 344984
rect 150434 344972 150440 344984
rect 150492 344972 150498 345024
rect 41322 344292 41328 344344
rect 41380 344332 41386 344344
rect 59078 344332 59084 344344
rect 41380 344304 59084 344332
rect 41380 344292 41386 344304
rect 59078 344292 59084 344304
rect 59136 344292 59142 344344
rect 150434 344292 150440 344344
rect 150492 344332 150498 344344
rect 188338 344332 188344 344344
rect 150492 344304 188344 344332
rect 150492 344292 150498 344304
rect 188338 344292 188344 344304
rect 188396 344292 188402 344344
rect 59078 343612 59084 343664
rect 59136 343652 59142 343664
rect 67634 343652 67640 343664
rect 59136 343624 67640 343652
rect 59136 343612 59142 343624
rect 67634 343612 67640 343624
rect 67692 343612 67698 343664
rect 117774 343544 117780 343596
rect 117832 343584 117838 343596
rect 139578 343584 139584 343596
rect 117832 343556 139584 343584
rect 117832 343544 117838 343556
rect 139578 343544 139584 343556
rect 139636 343544 139642 343596
rect 118602 342864 118608 342916
rect 118660 342904 118666 342916
rect 128722 342904 128728 342916
rect 118660 342876 128728 342904
rect 118660 342864 118666 342876
rect 128722 342864 128728 342876
rect 128780 342864 128786 342916
rect 139578 342864 139584 342916
rect 139636 342904 139642 342916
rect 193858 342904 193864 342916
rect 139636 342876 193864 342904
rect 139636 342864 139642 342876
rect 193858 342864 193864 342876
rect 193916 342864 193922 342916
rect 322474 342864 322480 342916
rect 322532 342904 322538 342916
rect 327258 342904 327264 342916
rect 322532 342876 327264 342904
rect 322532 342864 322538 342876
rect 327258 342864 327264 342876
rect 327316 342904 327322 342916
rect 352650 342904 352656 342916
rect 327316 342876 352656 342904
rect 327316 342864 327322 342876
rect 352650 342864 352656 342876
rect 352708 342864 352714 342916
rect 64598 342252 64604 342304
rect 64656 342292 64662 342304
rect 67634 342292 67640 342304
rect 64656 342264 67640 342292
rect 64656 342252 64662 342264
rect 67634 342252 67640 342264
rect 67692 342252 67698 342304
rect 323578 342292 323584 342304
rect 323491 342264 323584 342292
rect 323578 342252 323584 342264
rect 323636 342292 323642 342304
rect 493870 342292 493876 342304
rect 323636 342264 493876 342292
rect 323636 342252 323642 342264
rect 493870 342252 493876 342264
rect 493928 342252 493934 342304
rect 322842 342184 322848 342236
rect 322900 342224 322906 342236
rect 323596 342224 323624 342252
rect 322900 342196 323624 342224
rect 322900 342184 322906 342196
rect 118142 341572 118148 341624
rect 118200 341612 118206 341624
rect 131298 341612 131304 341624
rect 118200 341584 131304 341612
rect 118200 341572 118206 341584
rect 131298 341572 131304 341584
rect 131356 341572 131362 341624
rect 36998 341504 37004 341556
rect 37056 341544 37062 341556
rect 67910 341544 67916 341556
rect 37056 341516 67916 341544
rect 37056 341504 37062 341516
rect 67910 341504 67916 341516
rect 67968 341504 67974 341556
rect 118510 341504 118516 341556
rect 118568 341544 118574 341556
rect 138198 341544 138204 341556
rect 118568 341516 138204 341544
rect 118568 341504 118574 341516
rect 138198 341504 138204 341516
rect 138256 341504 138262 341556
rect 63402 340892 63408 340944
rect 63460 340932 63466 340944
rect 66162 340932 66168 340944
rect 63460 340904 66168 340932
rect 63460 340892 63466 340904
rect 66162 340892 66168 340904
rect 66220 340932 66226 340944
rect 67634 340932 67640 340944
rect 66220 340904 67640 340932
rect 66220 340892 66226 340904
rect 67634 340892 67640 340904
rect 67692 340892 67698 340944
rect 138198 340892 138204 340944
rect 138256 340932 138262 340944
rect 190454 340932 190460 340944
rect 138256 340904 190460 340932
rect 138256 340892 138262 340904
rect 190454 340892 190460 340904
rect 190512 340892 190518 340944
rect 117314 340824 117320 340876
rect 117372 340864 117378 340876
rect 135898 340864 135904 340876
rect 117372 340836 135904 340864
rect 117372 340824 117378 340836
rect 135898 340824 135904 340836
rect 135956 340824 135962 340876
rect 117406 340756 117412 340808
rect 117464 340796 117470 340808
rect 130010 340796 130016 340808
rect 117464 340768 130016 340796
rect 117464 340756 117470 340768
rect 130010 340756 130016 340768
rect 130068 340756 130074 340808
rect 69290 340688 69296 340740
rect 69348 340728 69354 340740
rect 69750 340728 69756 340740
rect 69348 340700 69756 340728
rect 69348 340688 69354 340700
rect 69750 340688 69756 340700
rect 69808 340688 69814 340740
rect 58618 340212 58624 340264
rect 58676 340252 58682 340264
rect 70394 340252 70400 340264
rect 58676 340224 70400 340252
rect 58676 340212 58682 340224
rect 70394 340212 70400 340224
rect 70452 340212 70458 340264
rect 43806 340144 43812 340196
rect 43864 340184 43870 340196
rect 43864 340156 64874 340184
rect 43864 340144 43870 340156
rect 64846 339912 64874 340156
rect 427814 340144 427820 340196
rect 427872 340184 427878 340196
rect 497458 340184 497464 340196
rect 427872 340156 497464 340184
rect 427872 340144 427878 340156
rect 497458 340144 497464 340156
rect 497516 340144 497522 340196
rect 75822 339912 75828 339924
rect 64846 339884 75828 339912
rect 75822 339872 75828 339884
rect 75880 339872 75886 339924
rect 61838 339532 61844 339584
rect 61896 339572 61902 339584
rect 64598 339572 64604 339584
rect 61896 339544 64604 339572
rect 61896 339532 61902 339544
rect 64598 339532 64604 339544
rect 64656 339572 64662 339584
rect 67634 339572 67640 339584
rect 64656 339544 67640 339572
rect 64656 339532 64662 339544
rect 67634 339532 67640 339544
rect 67692 339532 67698 339584
rect 111058 339532 111064 339584
rect 111116 339572 111122 339584
rect 115658 339572 115664 339584
rect 111116 339544 115664 339572
rect 111116 339532 111122 339544
rect 115658 339532 115664 339544
rect 115716 339532 115722 339584
rect 54846 339464 54852 339516
rect 54904 339504 54910 339516
rect 78398 339504 78404 339516
rect 54904 339476 78404 339504
rect 54904 339464 54910 339476
rect 78398 339464 78404 339476
rect 78456 339464 78462 339516
rect 107470 339464 107476 339516
rect 107528 339504 107534 339516
rect 117406 339504 117412 339516
rect 107528 339476 117412 339504
rect 107528 339464 107534 339476
rect 117406 339464 117412 339476
rect 117464 339464 117470 339516
rect 170490 339464 170496 339516
rect 170548 339504 170554 339516
rect 197354 339504 197360 339516
rect 170548 339476 197360 339504
rect 170548 339464 170554 339476
rect 197354 339464 197360 339476
rect 197412 339464 197418 339516
rect 46658 339396 46664 339448
rect 46716 339436 46722 339448
rect 52178 339436 52184 339448
rect 46716 339408 52184 339436
rect 46716 339396 46722 339408
rect 52178 339396 52184 339408
rect 52236 339436 52242 339448
rect 82262 339436 82268 339448
rect 52236 339408 82268 339436
rect 52236 339396 52242 339408
rect 82262 339396 82268 339408
rect 82320 339396 82326 339448
rect 87414 339396 87420 339448
rect 87472 339436 87478 339448
rect 87690 339436 87696 339448
rect 87472 339408 87696 339436
rect 87472 339396 87478 339408
rect 87690 339396 87696 339408
rect 87748 339436 87754 339448
rect 124858 339436 124864 339448
rect 87748 339408 124864 339436
rect 87748 339396 87754 339408
rect 124858 339396 124864 339408
rect 124916 339396 124922 339448
rect 194042 339436 194048 339448
rect 132466 339408 194048 339436
rect 60366 339328 60372 339380
rect 60424 339368 60430 339380
rect 92566 339368 92572 339380
rect 60424 339340 92572 339368
rect 60424 339328 60430 339340
rect 92566 339328 92572 339340
rect 92624 339368 92630 339380
rect 93118 339368 93124 339380
rect 92624 339340 93124 339368
rect 92624 339328 92630 339340
rect 93118 339328 93124 339340
rect 93176 339328 93182 339380
rect 94590 339328 94596 339380
rect 94648 339368 94654 339380
rect 95142 339368 95148 339380
rect 94648 339340 95148 339368
rect 94648 339328 94654 339340
rect 95142 339328 95148 339340
rect 95200 339368 95206 339380
rect 128446 339368 128452 339380
rect 95200 339340 128452 339368
rect 95200 339328 95206 339340
rect 128446 339328 128452 339340
rect 128504 339368 128510 339380
rect 132466 339368 132494 339408
rect 194042 339396 194048 339408
rect 194100 339396 194106 339448
rect 128504 339340 132494 339368
rect 128504 339328 128510 339340
rect 46198 339260 46204 339312
rect 46256 339300 46262 339312
rect 73890 339300 73896 339312
rect 46256 339272 73896 339300
rect 46256 339260 46262 339272
rect 73890 339260 73896 339272
rect 73948 339260 73954 339312
rect 113174 339260 113180 339312
rect 113232 339300 113238 339312
rect 113726 339300 113732 339312
rect 113232 339272 113732 339300
rect 113232 339260 113238 339272
rect 113726 339260 113732 339272
rect 113784 339300 113790 339312
rect 138014 339300 138020 339312
rect 113784 339272 138020 339300
rect 113784 339260 113790 339272
rect 138014 339260 138020 339272
rect 138072 339260 138078 339312
rect 52086 339192 52092 339244
rect 52144 339232 52150 339244
rect 76466 339232 76472 339244
rect 52144 339204 76472 339232
rect 52144 339192 52150 339204
rect 76466 339192 76472 339204
rect 76524 339192 76530 339244
rect 105446 339192 105452 339244
rect 105504 339232 105510 339244
rect 106182 339232 106188 339244
rect 105504 339204 106188 339232
rect 105504 339192 105510 339204
rect 106182 339192 106188 339204
rect 106240 339232 106246 339244
rect 117498 339232 117504 339244
rect 106240 339204 117504 339232
rect 106240 339192 106246 339204
rect 117498 339192 117504 339204
rect 117556 339192 117562 339244
rect 68830 338784 68836 338836
rect 68888 338824 68894 338836
rect 98638 338824 98644 338836
rect 68888 338796 98644 338824
rect 68888 338784 68894 338796
rect 98638 338784 98644 338796
rect 98696 338784 98702 338836
rect 66990 338716 66996 338768
rect 67048 338756 67054 338768
rect 77478 338756 77484 338768
rect 67048 338728 77484 338756
rect 67048 338716 67054 338728
rect 77478 338716 77484 338728
rect 77536 338716 77542 338768
rect 91738 338716 91744 338768
rect 91796 338756 91802 338768
rect 121638 338756 121644 338768
rect 91796 338728 121644 338756
rect 91796 338716 91802 338728
rect 121638 338716 121644 338728
rect 121696 338716 121702 338768
rect 323026 338376 323032 338428
rect 323084 338416 323090 338428
rect 323578 338416 323584 338428
rect 323084 338388 323584 338416
rect 323084 338376 323090 338388
rect 323578 338376 323584 338388
rect 323636 338376 323642 338428
rect 79686 338240 79692 338292
rect 79744 338280 79750 338292
rect 83642 338280 83648 338292
rect 79744 338252 83648 338280
rect 79744 338240 79750 338252
rect 83642 338240 83648 338252
rect 83700 338240 83706 338292
rect 76466 338172 76472 338224
rect 76524 338212 76530 338224
rect 83458 338212 83464 338224
rect 76524 338184 83464 338212
rect 76524 338172 76530 338184
rect 83458 338172 83464 338184
rect 83516 338172 83522 338224
rect 87598 338144 87604 338156
rect 84166 338116 87604 338144
rect 49418 337968 49424 338020
rect 49476 338008 49482 338020
rect 83550 338008 83556 338020
rect 49476 337980 83556 338008
rect 49476 337968 49482 337980
rect 83550 337968 83556 337980
rect 83608 338008 83614 338020
rect 84166 338008 84194 338116
rect 87598 338104 87604 338116
rect 87656 338104 87662 338156
rect 113818 338036 113824 338088
rect 113876 338076 113882 338088
rect 118050 338076 118056 338088
rect 113876 338048 118056 338076
rect 113876 338036 113882 338048
rect 118050 338036 118056 338048
rect 118108 338036 118114 338088
rect 199470 338076 199476 338088
rect 135732 338048 199476 338076
rect 83608 337980 84194 338008
rect 83608 337968 83614 337980
rect 112530 337968 112536 338020
rect 112588 338008 112594 338020
rect 135346 338008 135352 338020
rect 112588 337980 135352 338008
rect 112588 337968 112594 337980
rect 135346 337968 135352 337980
rect 135404 338008 135410 338020
rect 135622 338008 135628 338020
rect 135404 337980 135628 338008
rect 135404 337968 135410 337980
rect 135622 337968 135628 337980
rect 135680 337968 135686 338020
rect 45186 337900 45192 337952
rect 45244 337940 45250 337952
rect 74534 337940 74540 337952
rect 45244 337912 74540 337940
rect 45244 337900 45250 337912
rect 74534 337900 74540 337912
rect 74592 337940 74598 337952
rect 75270 337940 75276 337952
rect 74592 337912 75276 337940
rect 74592 337900 74598 337912
rect 75270 337900 75276 337912
rect 75328 337900 75334 337952
rect 119430 337940 119436 337952
rect 103486 337912 119436 337940
rect 42058 337832 42064 337884
rect 42116 337872 42122 337884
rect 70486 337872 70492 337884
rect 42116 337844 70492 337872
rect 42116 337832 42122 337844
rect 70486 337832 70492 337844
rect 70544 337832 70550 337884
rect 57882 337764 57888 337816
rect 57940 337804 57946 337816
rect 84194 337804 84200 337816
rect 57940 337776 84200 337804
rect 57940 337764 57946 337776
rect 84194 337764 84200 337776
rect 84252 337764 84258 337816
rect 99650 337764 99656 337816
rect 99708 337804 99714 337816
rect 100662 337804 100668 337816
rect 99708 337776 100668 337804
rect 99708 337764 99714 337776
rect 100662 337764 100668 337776
rect 100720 337804 100726 337816
rect 103486 337804 103514 337912
rect 119430 337900 119436 337912
rect 119488 337900 119494 337952
rect 104802 337832 104808 337884
rect 104860 337872 104866 337884
rect 132678 337872 132684 337884
rect 104860 337844 132684 337872
rect 104860 337832 104866 337844
rect 132678 337832 132684 337844
rect 132736 337872 132742 337884
rect 135732 337872 135760 338048
rect 199470 338036 199476 338048
rect 199528 338036 199534 338088
rect 136634 337968 136640 338020
rect 136692 338008 136698 338020
rect 136818 338008 136824 338020
rect 136692 337980 136824 338008
rect 136692 337968 136698 337980
rect 136818 337968 136824 337980
rect 136876 338008 136882 338020
rect 196710 338008 196716 338020
rect 136876 337980 196716 338008
rect 136876 337968 136882 337980
rect 196710 337968 196716 337980
rect 196768 337968 196774 338020
rect 132736 337844 135760 337872
rect 132736 337832 132742 337844
rect 100720 337776 103514 337804
rect 100720 337764 100726 337776
rect 50706 337696 50712 337748
rect 50764 337736 50770 337748
rect 86126 337736 86132 337748
rect 50764 337708 86132 337736
rect 50764 337696 50770 337708
rect 86126 337696 86132 337708
rect 86184 337736 86190 337748
rect 86862 337736 86868 337748
rect 86184 337708 86868 337736
rect 86184 337696 86190 337708
rect 86862 337696 86868 337708
rect 86920 337696 86926 337748
rect 91278 337696 91284 337748
rect 91336 337736 91342 337748
rect 103606 337736 103612 337748
rect 91336 337708 103612 337736
rect 91336 337696 91342 337708
rect 103606 337696 103612 337708
rect 103664 337696 103670 337748
rect 109954 337696 109960 337748
rect 110012 337736 110018 337748
rect 111794 337736 111800 337748
rect 110012 337708 111800 337736
rect 110012 337696 110018 337708
rect 111794 337696 111800 337708
rect 111852 337696 111858 337748
rect 75822 337492 75828 337544
rect 75880 337532 75886 337544
rect 104158 337532 104164 337544
rect 75880 337504 104164 337532
rect 75880 337492 75886 337504
rect 104158 337492 104164 337504
rect 104216 337492 104222 337544
rect 107378 337492 107384 337544
rect 107436 337532 107442 337544
rect 110230 337532 110236 337544
rect 107436 337504 110236 337532
rect 107436 337492 107442 337504
rect 110230 337492 110236 337504
rect 110288 337492 110294 337544
rect 78398 337424 78404 337476
rect 78456 337464 78462 337476
rect 98730 337464 98736 337476
rect 78456 337436 98736 337464
rect 78456 337424 78462 337436
rect 98730 337424 98736 337436
rect 98788 337424 98794 337476
rect 103514 337424 103520 337476
rect 103572 337464 103578 337476
rect 133874 337464 133880 337476
rect 103572 337436 133880 337464
rect 103572 337424 103578 337436
rect 133874 337424 133880 337436
rect 133932 337464 133938 337476
rect 136634 337464 136640 337476
rect 133932 337436 136640 337464
rect 133932 337424 133938 337436
rect 136634 337424 136640 337436
rect 136692 337424 136698 337476
rect 91002 337356 91008 337408
rect 91060 337396 91066 337408
rect 91922 337396 91928 337408
rect 91060 337368 91928 337396
rect 91060 337356 91066 337368
rect 91922 337356 91928 337368
rect 91980 337356 91986 337408
rect 131206 337396 131212 337408
rect 93826 337368 131212 337396
rect 82814 337288 82820 337340
rect 82872 337328 82878 337340
rect 84838 337328 84844 337340
rect 82872 337300 84844 337328
rect 82872 337288 82878 337300
rect 84838 337288 84844 337300
rect 84896 337288 84902 337340
rect 86862 337288 86868 337340
rect 86920 337328 86926 337340
rect 93826 337328 93854 337368
rect 131206 337356 131212 337368
rect 131264 337396 131270 337408
rect 134518 337396 134524 337408
rect 131264 337368 134524 337396
rect 131264 337356 131270 337368
rect 134518 337356 134524 337368
rect 134576 337356 134582 337408
rect 135622 337356 135628 337408
rect 135680 337396 135686 337408
rect 185670 337396 185676 337408
rect 135680 337368 185676 337396
rect 135680 337356 135686 337368
rect 185670 337356 185676 337368
rect 185728 337356 185734 337408
rect 86920 337300 93854 337328
rect 86920 337288 86926 337300
rect 103054 337220 103060 337272
rect 103112 337260 103118 337272
rect 104802 337260 104808 337272
rect 103112 337232 104808 337260
rect 103112 337220 103118 337232
rect 104802 337220 104808 337232
rect 104860 337220 104866 337272
rect 70026 337084 70032 337136
rect 70084 337124 70090 337136
rect 76558 337124 76564 337136
rect 70084 337096 76564 337124
rect 70084 337084 70090 337096
rect 76558 337084 76564 337096
rect 76616 337084 76622 337136
rect 111610 336744 111616 336796
rect 111668 336784 111674 336796
rect 113818 336784 113824 336796
rect 111668 336756 113824 336784
rect 111668 336744 111674 336756
rect 113818 336744 113824 336756
rect 113876 336744 113882 336796
rect 195054 336744 195060 336796
rect 195112 336784 195118 336796
rect 197354 336784 197360 336796
rect 195112 336756 197360 336784
rect 195112 336744 195118 336756
rect 197354 336744 197360 336756
rect 197412 336744 197418 336796
rect 46842 336676 46848 336728
rect 46900 336716 46906 336728
rect 80790 336716 80796 336728
rect 46900 336688 80796 336716
rect 46900 336676 46906 336688
rect 80790 336676 80796 336688
rect 80848 336676 80854 336728
rect 100938 336676 100944 336728
rect 100996 336716 101002 336728
rect 101950 336716 101956 336728
rect 100996 336688 101956 336716
rect 100996 336676 101002 336688
rect 101950 336676 101956 336688
rect 102008 336716 102014 336728
rect 102008 336688 103514 336716
rect 102008 336676 102014 336688
rect 56410 336608 56416 336660
rect 56468 336648 56474 336660
rect 88978 336648 88984 336660
rect 56468 336620 88984 336648
rect 56468 336608 56474 336620
rect 88978 336608 88984 336620
rect 89036 336608 89042 336660
rect 103486 336648 103514 336688
rect 110598 336676 110604 336728
rect 110656 336716 110662 336728
rect 111702 336716 111708 336728
rect 110656 336688 111708 336716
rect 110656 336676 110662 336688
rect 111702 336676 111708 336688
rect 111760 336676 111766 336728
rect 111794 336676 111800 336728
rect 111852 336716 111858 336728
rect 133966 336716 133972 336728
rect 111852 336688 133972 336716
rect 111852 336676 111858 336688
rect 133966 336676 133972 336688
rect 134024 336676 134030 336728
rect 322474 336676 322480 336728
rect 322532 336716 322538 336728
rect 327166 336716 327172 336728
rect 322532 336688 327172 336716
rect 322532 336676 322538 336688
rect 327166 336676 327172 336688
rect 327224 336716 327230 336728
rect 328362 336716 328368 336728
rect 327224 336688 328368 336716
rect 327224 336676 327230 336688
rect 328362 336676 328368 336688
rect 328420 336676 328426 336728
rect 127250 336648 127256 336660
rect 103486 336620 127256 336648
rect 127250 336608 127256 336620
rect 127308 336608 127314 336660
rect 52178 336540 52184 336592
rect 52236 336580 52242 336592
rect 54754 336580 54760 336592
rect 52236 336552 54760 336580
rect 52236 336540 52242 336552
rect 54754 336540 54760 336552
rect 54812 336580 54818 336592
rect 82814 336580 82820 336592
rect 54812 336552 82820 336580
rect 54812 336540 54818 336552
rect 82814 336540 82820 336552
rect 82872 336540 82878 336592
rect 100294 336540 100300 336592
rect 100352 336580 100358 336592
rect 125778 336580 125784 336592
rect 100352 336552 125784 336580
rect 100352 336540 100358 336552
rect 125778 336540 125784 336552
rect 125836 336580 125842 336592
rect 126882 336580 126888 336592
rect 125836 336552 126888 336580
rect 125836 336540 125842 336552
rect 126882 336540 126888 336552
rect 126940 336540 126946 336592
rect 70394 336472 70400 336524
rect 70452 336512 70458 336524
rect 90358 336512 90364 336524
rect 70452 336484 90364 336512
rect 70452 336472 70458 336484
rect 90358 336472 90364 336484
rect 90416 336472 90422 336524
rect 97902 336472 97908 336524
rect 97960 336512 97966 336524
rect 117958 336512 117964 336524
rect 97960 336484 117964 336512
rect 97960 336472 97966 336484
rect 117958 336472 117964 336484
rect 118016 336472 118022 336524
rect 50798 336404 50804 336456
rect 50856 336444 50862 336456
rect 71958 336444 71964 336456
rect 50856 336416 71964 336444
rect 50856 336404 50862 336416
rect 71958 336404 71964 336416
rect 72016 336444 72022 336456
rect 72418 336444 72424 336456
rect 72016 336416 72424 336444
rect 72016 336404 72022 336416
rect 72418 336404 72424 336416
rect 72476 336404 72482 336456
rect 111702 336404 111708 336456
rect 111760 336444 111766 336456
rect 124398 336444 124404 336456
rect 111760 336416 124404 336444
rect 111760 336404 111766 336416
rect 124398 336404 124404 336416
rect 124456 336404 124462 336456
rect 47578 336336 47584 336388
rect 47636 336376 47642 336388
rect 71314 336376 71320 336388
rect 47636 336348 71320 336376
rect 47636 336336 47642 336348
rect 71314 336336 71320 336348
rect 71372 336336 71378 336388
rect 106090 336336 106096 336388
rect 106148 336376 106154 336388
rect 111794 336376 111800 336388
rect 106148 336348 111800 336376
rect 106148 336336 106154 336348
rect 111794 336336 111800 336348
rect 111852 336336 111858 336388
rect 59078 335996 59084 336048
rect 59136 336036 59142 336048
rect 77386 336036 77392 336048
rect 59136 336008 77392 336036
rect 59136 335996 59142 336008
rect 77386 335996 77392 336008
rect 77444 335996 77450 336048
rect 86218 335996 86224 336048
rect 86276 336036 86282 336048
rect 121546 336036 121552 336048
rect 86276 336008 121552 336036
rect 86276 335996 86282 336008
rect 121546 335996 121552 336008
rect 121604 335996 121610 336048
rect 126882 335996 126888 336048
rect 126940 336036 126946 336048
rect 136726 336036 136732 336048
rect 126940 336008 136732 336036
rect 126940 335996 126946 336008
rect 136726 335996 136732 336008
rect 136784 335996 136790 336048
rect 328362 335996 328368 336048
rect 328420 336036 328426 336048
rect 388438 336036 388444 336048
rect 328420 336008 388444 336036
rect 328420 335996 328426 336008
rect 388438 335996 388444 336008
rect 388496 335996 388502 336048
rect 173158 335316 173164 335368
rect 173216 335356 173222 335368
rect 197354 335356 197360 335368
rect 173216 335328 197360 335356
rect 173216 335316 173222 335328
rect 197354 335316 197360 335328
rect 197412 335316 197418 335368
rect 53558 335248 53564 335300
rect 53616 335288 53622 335300
rect 87690 335288 87696 335300
rect 53616 335260 87696 335288
rect 53616 335248 53622 335260
rect 87690 335248 87696 335260
rect 87748 335248 87754 335300
rect 115106 335248 115112 335300
rect 115164 335288 115170 335300
rect 141142 335288 141148 335300
rect 115164 335260 141148 335288
rect 115164 335248 115170 335260
rect 141142 335248 141148 335260
rect 141200 335248 141206 335300
rect 53466 335180 53472 335232
rect 53524 335220 53530 335232
rect 86310 335220 86316 335232
rect 53524 335192 86316 335220
rect 53524 335180 53530 335192
rect 86310 335180 86316 335192
rect 86368 335180 86374 335232
rect 140682 335180 140688 335232
rect 140740 335220 140746 335232
rect 195054 335220 195060 335232
rect 140740 335192 195060 335220
rect 140740 335180 140746 335192
rect 195054 335180 195060 335192
rect 195112 335180 195118 335232
rect 41230 335112 41236 335164
rect 41288 335152 41294 335164
rect 71774 335152 71780 335164
rect 41288 335124 71780 335152
rect 41288 335112 41294 335124
rect 71774 335112 71780 335124
rect 71832 335152 71838 335164
rect 73062 335152 73068 335164
rect 71832 335124 73068 335152
rect 71832 335112 71838 335124
rect 73062 335112 73068 335124
rect 73120 335112 73126 335164
rect 86310 334772 86316 334824
rect 86368 334812 86374 334824
rect 86770 334812 86776 334824
rect 86368 334784 86776 334812
rect 86368 334772 86374 334784
rect 86770 334772 86776 334784
rect 86828 334772 86834 334824
rect 98362 334704 98368 334756
rect 98420 334744 98426 334756
rect 126422 334744 126428 334756
rect 98420 334716 126428 334744
rect 98420 334704 98426 334716
rect 126422 334704 126428 334716
rect 126480 334744 126486 334756
rect 131482 334744 131488 334756
rect 126480 334716 131488 334744
rect 126480 334704 126486 334716
rect 131482 334704 131488 334716
rect 131540 334704 131546 334756
rect 140130 334704 140136 334756
rect 140188 334744 140194 334756
rect 140682 334744 140688 334756
rect 140188 334716 140688 334744
rect 140188 334704 140194 334716
rect 140682 334704 140688 334716
rect 140740 334704 140746 334756
rect 69658 334636 69664 334688
rect 69716 334676 69722 334688
rect 109034 334676 109040 334688
rect 69716 334648 109040 334676
rect 69716 334636 69722 334648
rect 109034 334636 109040 334648
rect 109092 334636 109098 334688
rect 54846 334568 54852 334620
rect 54904 334608 54910 334620
rect 103054 334608 103060 334620
rect 54904 334580 103060 334608
rect 54904 334568 54910 334580
rect 103054 334568 103060 334580
rect 103112 334568 103118 334620
rect 129734 334568 129740 334620
rect 129792 334608 129798 334620
rect 140866 334608 140872 334620
rect 129792 334580 140872 334608
rect 129792 334568 129798 334580
rect 140866 334568 140872 334580
rect 140924 334568 140930 334620
rect 321738 334568 321744 334620
rect 321796 334608 321802 334620
rect 328454 334608 328460 334620
rect 321796 334580 328460 334608
rect 321796 334568 321802 334580
rect 328454 334568 328460 334580
rect 328512 334568 328518 334620
rect 48038 333956 48044 334008
rect 48096 333996 48102 334008
rect 53558 333996 53564 334008
rect 48096 333968 53564 333996
rect 48096 333956 48102 333968
rect 53558 333956 53564 333968
rect 53616 333956 53622 334008
rect 115106 333956 115112 334008
rect 115164 333996 115170 334008
rect 115382 333996 115388 334008
rect 115164 333968 115388 333996
rect 115164 333956 115170 333968
rect 115382 333956 115388 333968
rect 115440 333956 115446 334008
rect 51994 333888 52000 333940
rect 52052 333928 52058 333940
rect 89070 333928 89076 333940
rect 52052 333900 89076 333928
rect 52052 333888 52058 333900
rect 89070 333888 89076 333900
rect 89128 333888 89134 333940
rect 108022 333888 108028 333940
rect 108080 333928 108086 333940
rect 131390 333928 131396 333940
rect 108080 333900 131396 333928
rect 108080 333888 108086 333900
rect 131390 333888 131396 333900
rect 131448 333888 131454 333940
rect 45462 333820 45468 333872
rect 45520 333860 45526 333872
rect 76650 333860 76656 333872
rect 45520 333832 76656 333860
rect 45520 333820 45526 333832
rect 76650 333820 76656 333832
rect 76708 333820 76714 333872
rect 60458 333752 60464 333804
rect 60516 333792 60522 333804
rect 81618 333792 81624 333804
rect 60516 333764 81624 333792
rect 60516 333752 60522 333764
rect 81618 333752 81624 333764
rect 81676 333752 81682 333804
rect 76650 333412 76656 333464
rect 76708 333452 76714 333464
rect 77110 333452 77116 333464
rect 76708 333424 77116 333452
rect 76708 333412 76714 333424
rect 77110 333412 77116 333424
rect 77168 333412 77174 333464
rect 107562 333276 107568 333328
rect 107620 333316 107626 333328
rect 115934 333316 115940 333328
rect 107620 333288 115940 333316
rect 107620 333276 107626 333288
rect 115934 333276 115940 333288
rect 115992 333276 115998 333328
rect 109034 333208 109040 333260
rect 109092 333248 109098 333260
rect 136634 333248 136640 333260
rect 109092 333220 136640 333248
rect 109092 333208 109098 333220
rect 136634 333208 136640 333220
rect 136692 333248 136698 333260
rect 166258 333248 166264 333260
rect 136692 333220 166264 333248
rect 136692 333208 136698 333220
rect 166258 333208 166264 333220
rect 166316 333208 166322 333260
rect 352650 333208 352656 333260
rect 352708 333248 352714 333260
rect 465074 333248 465080 333260
rect 352708 333220 465080 333248
rect 352708 333208 352714 333220
rect 465074 333208 465080 333220
rect 465132 333208 465138 333260
rect 81618 332664 81624 332716
rect 81676 332704 81682 332716
rect 82078 332704 82084 332716
rect 81676 332676 82084 332704
rect 81676 332664 81682 332676
rect 82078 332664 82084 332676
rect 82136 332664 82142 332716
rect 73798 332596 73804 332648
rect 73856 332636 73862 332648
rect 198826 332636 198832 332648
rect 73856 332608 198832 332636
rect 73856 332596 73862 332608
rect 198826 332596 198832 332608
rect 198884 332636 198890 332648
rect 199010 332636 199016 332648
rect 198884 332608 199016 332636
rect 198884 332596 198890 332608
rect 199010 332596 199016 332608
rect 199068 332596 199074 332648
rect 46750 332528 46756 332580
rect 46808 332568 46814 332580
rect 79410 332568 79416 332580
rect 46808 332540 79416 332568
rect 46808 332528 46814 332540
rect 79410 332528 79416 332540
rect 79468 332528 79474 332580
rect 94498 332528 94504 332580
rect 94556 332568 94562 332580
rect 124214 332568 124220 332580
rect 94556 332540 124220 332568
rect 94556 332528 94562 332540
rect 124214 332528 124220 332540
rect 124272 332568 124278 332580
rect 126974 332568 126980 332580
rect 124272 332540 126980 332568
rect 124272 332528 124278 332540
rect 126974 332528 126980 332540
rect 127032 332528 127038 332580
rect 188522 332528 188528 332580
rect 188580 332568 188586 332580
rect 198090 332568 198096 332580
rect 188580 332540 198096 332568
rect 188580 332528 188586 332540
rect 198090 332528 198096 332540
rect 198148 332528 198154 332580
rect 97810 332460 97816 332512
rect 97868 332500 97874 332512
rect 118142 332500 118148 332512
rect 97868 332472 118148 332500
rect 97868 332460 97874 332472
rect 118142 332460 118148 332472
rect 118200 332460 118206 332512
rect 97074 331916 97080 331968
rect 97132 331956 97138 331968
rect 97810 331956 97816 331968
rect 97132 331928 97816 331956
rect 97132 331916 97138 331928
rect 97810 331916 97816 331928
rect 97868 331916 97874 331968
rect 37090 331848 37096 331900
rect 37148 331888 37154 331900
rect 108022 331888 108028 331900
rect 37148 331860 108028 331888
rect 37148 331848 37154 331860
rect 108022 331848 108028 331860
rect 108080 331848 108086 331900
rect 322198 331712 322204 331764
rect 322256 331752 322262 331764
rect 325694 331752 325700 331764
rect 322256 331724 325700 331752
rect 322256 331712 322262 331724
rect 325694 331712 325700 331724
rect 325752 331712 325758 331764
rect 7558 331236 7564 331288
rect 7616 331276 7622 331288
rect 37090 331276 37096 331288
rect 7616 331248 37096 331276
rect 7616 331236 7622 331248
rect 37090 331236 37096 331248
rect 37148 331236 37154 331288
rect 122190 331236 122196 331288
rect 122248 331276 122254 331288
rect 122650 331276 122656 331288
rect 122248 331248 122656 331276
rect 122248 331236 122254 331248
rect 122650 331236 122656 331248
rect 122708 331276 122714 331288
rect 165522 331276 165528 331288
rect 122708 331248 165528 331276
rect 122708 331236 122714 331248
rect 165522 331236 165528 331248
rect 165580 331276 165586 331288
rect 197354 331276 197360 331288
rect 165580 331248 197360 331276
rect 165580 331236 165586 331248
rect 197354 331236 197360 331248
rect 197412 331236 197418 331288
rect 93210 331168 93216 331220
rect 93268 331208 93274 331220
rect 120810 331208 120816 331220
rect 93268 331180 120816 331208
rect 93268 331168 93274 331180
rect 120810 331168 120816 331180
rect 120868 331208 120874 331220
rect 124214 331208 124220 331220
rect 120868 331180 124220 331208
rect 120868 331168 120874 331180
rect 124214 331168 124220 331180
rect 124272 331168 124278 331220
rect 104894 330760 104900 330812
rect 104952 330800 104958 330812
rect 128630 330800 128636 330812
rect 104952 330772 128636 330800
rect 104952 330760 104958 330772
rect 128630 330760 128636 330772
rect 128688 330760 128694 330812
rect 69106 330692 69112 330744
rect 69164 330732 69170 330744
rect 115198 330732 115204 330744
rect 69164 330704 115204 330732
rect 69164 330692 69170 330704
rect 115198 330692 115204 330704
rect 115256 330692 115262 330744
rect 129734 330692 129740 330744
rect 129792 330732 129798 330744
rect 169202 330732 169208 330744
rect 129792 330704 169208 330732
rect 129792 330692 129798 330704
rect 169202 330692 169208 330704
rect 169260 330692 169266 330744
rect 111794 330624 111800 330676
rect 111852 330664 111858 330676
rect 182910 330664 182916 330676
rect 111852 330636 182916 330664
rect 111852 330624 111858 330636
rect 182910 330624 182916 330636
rect 182968 330624 182974 330676
rect 66162 330556 66168 330608
rect 66220 330596 66226 330608
rect 151078 330596 151084 330608
rect 66220 330568 151084 330596
rect 66220 330556 66226 330568
rect 151078 330556 151084 330568
rect 151136 330556 151142 330608
rect 60550 330488 60556 330540
rect 60608 330528 60614 330540
rect 191098 330528 191104 330540
rect 60608 330500 191104 330528
rect 60608 330488 60614 330500
rect 191098 330488 191104 330500
rect 191156 330488 191162 330540
rect 322198 330488 322204 330540
rect 322256 330528 322262 330540
rect 325786 330528 325792 330540
rect 322256 330500 325792 330528
rect 322256 330488 322262 330500
rect 325786 330488 325792 330500
rect 325844 330528 325850 330540
rect 328546 330528 328552 330540
rect 325844 330500 328552 330528
rect 325844 330488 325850 330500
rect 328546 330488 328552 330500
rect 328604 330488 328610 330540
rect 129734 329848 129740 329860
rect 117976 329820 129740 329848
rect 56502 329740 56508 329792
rect 56560 329780 56566 329792
rect 117976 329780 118004 329820
rect 129734 329808 129740 329820
rect 129792 329808 129798 329860
rect 56560 329752 118004 329780
rect 56560 329740 56566 329752
rect 123662 329740 123668 329792
rect 123720 329780 123726 329792
rect 124306 329780 124312 329792
rect 123720 329752 124312 329780
rect 123720 329740 123726 329752
rect 124306 329740 124312 329752
rect 124364 329740 124370 329792
rect 55122 329128 55128 329180
rect 55180 329168 55186 329180
rect 94590 329168 94596 329180
rect 55180 329140 94596 329168
rect 55180 329128 55186 329140
rect 94590 329128 94596 329140
rect 94648 329128 94654 329180
rect 85574 329060 85580 329112
rect 85632 329100 85638 329112
rect 199378 329100 199384 329112
rect 85632 329072 199384 329100
rect 85632 329060 85638 329072
rect 199378 329060 199384 329072
rect 199436 329060 199442 329112
rect 124306 328448 124312 328500
rect 124364 328488 124370 328500
rect 169662 328488 169668 328500
rect 124364 328460 169668 328488
rect 124364 328448 124370 328460
rect 169662 328448 169668 328460
rect 169720 328488 169726 328500
rect 197354 328488 197360 328500
rect 169720 328460 197360 328488
rect 169720 328448 169726 328460
rect 197354 328448 197360 328460
rect 197412 328448 197418 328500
rect 107746 327904 107752 327956
rect 107804 327944 107810 327956
rect 162210 327944 162216 327956
rect 107804 327916 162216 327944
rect 107804 327904 107810 327916
rect 162210 327904 162216 327916
rect 162268 327904 162274 327956
rect 171962 327904 171968 327956
rect 172020 327944 172026 327956
rect 198274 327944 198280 327956
rect 172020 327916 198280 327944
rect 172020 327904 172026 327916
rect 198274 327904 198280 327916
rect 198332 327904 198338 327956
rect 66898 327836 66904 327888
rect 66956 327876 66962 327888
rect 122098 327876 122104 327888
rect 66956 327848 122104 327876
rect 66956 327836 66962 327848
rect 122098 327836 122104 327848
rect 122156 327836 122162 327888
rect 57790 327768 57796 327820
rect 57848 327808 57854 327820
rect 111058 327808 111064 327820
rect 57848 327780 111064 327808
rect 57848 327768 57854 327780
rect 111058 327768 111064 327780
rect 111116 327768 111122 327820
rect 112438 327768 112444 327820
rect 112496 327808 112502 327820
rect 171778 327808 171784 327820
rect 112496 327780 171784 327808
rect 112496 327768 112502 327780
rect 171778 327768 171784 327780
rect 171836 327768 171842 327820
rect 103606 327700 103612 327752
rect 103664 327740 103670 327752
rect 169110 327740 169116 327752
rect 103664 327712 169116 327740
rect 103664 327700 103670 327712
rect 169110 327700 169116 327712
rect 169168 327700 169174 327752
rect 322842 327700 322848 327752
rect 322900 327740 322906 327752
rect 324406 327740 324412 327752
rect 322900 327712 324412 327740
rect 322900 327700 322906 327712
rect 324406 327700 324412 327712
rect 324464 327740 324470 327752
rect 482278 327740 482284 327752
rect 324464 327712 482284 327740
rect 324464 327700 324470 327712
rect 482278 327700 482284 327712
rect 482336 327700 482342 327752
rect 195514 327088 195520 327140
rect 195572 327128 195578 327140
rect 197354 327128 197360 327140
rect 195572 327100 197360 327128
rect 195572 327088 195578 327100
rect 197354 327088 197360 327100
rect 197412 327088 197418 327140
rect 56502 326476 56508 326528
rect 56560 326516 56566 326528
rect 132494 326516 132500 326528
rect 56560 326488 132500 326516
rect 56560 326476 56566 326488
rect 132494 326476 132500 326488
rect 132552 326476 132558 326528
rect 88334 326408 88340 326460
rect 88392 326448 88398 326460
rect 171870 326448 171876 326460
rect 88392 326420 171876 326448
rect 88392 326408 88398 326420
rect 171870 326408 171876 326420
rect 171928 326408 171934 326460
rect 70394 326340 70400 326392
rect 70452 326380 70458 326392
rect 195422 326380 195428 326392
rect 70452 326352 195428 326380
rect 70452 326340 70458 326352
rect 195422 326340 195428 326352
rect 195480 326340 195486 326392
rect 110322 325660 110328 325712
rect 110380 325700 110386 325712
rect 115290 325700 115296 325712
rect 110380 325672 115296 325700
rect 110380 325660 110386 325672
rect 115290 325660 115296 325672
rect 115348 325660 115354 325712
rect 170582 325660 170588 325712
rect 170640 325700 170646 325712
rect 173158 325700 173164 325712
rect 170640 325672 173164 325700
rect 170640 325660 170646 325672
rect 173158 325660 173164 325672
rect 173216 325660 173222 325712
rect 104710 324980 104716 325032
rect 104768 325020 104774 325032
rect 128538 325020 128544 325032
rect 104768 324992 128544 325020
rect 104768 324980 104774 324992
rect 128538 324980 128544 324992
rect 128596 325020 128602 325032
rect 128596 324992 132494 325020
rect 128596 324980 128602 324992
rect 52086 324912 52092 324964
rect 52144 324952 52150 324964
rect 122190 324952 122196 324964
rect 52144 324924 122196 324952
rect 52144 324912 52150 324924
rect 122190 324912 122196 324924
rect 122248 324912 122254 324964
rect 132466 324952 132494 324992
rect 162210 324952 162216 324964
rect 132466 324924 162216 324952
rect 162210 324912 162216 324924
rect 162268 324912 162274 324964
rect 322750 324912 322756 324964
rect 322808 324952 322814 324964
rect 323210 324952 323216 324964
rect 322808 324924 323216 324952
rect 322808 324912 322814 324924
rect 323210 324912 323216 324924
rect 323268 324952 323274 324964
rect 329834 324952 329840 324964
rect 323268 324924 329840 324952
rect 323268 324912 323274 324924
rect 329834 324912 329840 324924
rect 329892 324912 329898 324964
rect 334618 324912 334624 324964
rect 334676 324952 334682 324964
rect 375926 324952 375932 324964
rect 334676 324924 375932 324952
rect 334676 324912 334682 324924
rect 375926 324912 375932 324924
rect 375984 324912 375990 324964
rect 375926 324300 375932 324352
rect 375984 324340 375990 324352
rect 376662 324340 376668 324352
rect 375984 324312 376668 324340
rect 375984 324300 375990 324312
rect 376662 324300 376668 324312
rect 376720 324340 376726 324352
rect 580166 324340 580172 324352
rect 376720 324312 580172 324340
rect 376720 324300 376726 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 79318 323688 79324 323740
rect 79376 323728 79382 323740
rect 104710 323728 104716 323740
rect 79376 323700 104716 323728
rect 79376 323688 79382 323700
rect 104710 323688 104716 323700
rect 104768 323688 104774 323740
rect 75270 323620 75276 323672
rect 75328 323660 75334 323672
rect 114554 323660 114560 323672
rect 75328 323632 114560 323660
rect 75328 323620 75334 323632
rect 114554 323620 114560 323632
rect 114612 323660 114618 323672
rect 160830 323660 160836 323672
rect 114612 323632 160836 323660
rect 114612 323620 114618 323632
rect 160830 323620 160836 323632
rect 160888 323620 160894 323672
rect 80698 323552 80704 323604
rect 80756 323592 80762 323604
rect 189810 323592 189816 323604
rect 80756 323564 189816 323592
rect 80756 323552 80762 323564
rect 189810 323552 189816 323564
rect 189868 323552 189874 323604
rect 322474 322940 322480 322992
rect 322532 322980 322538 322992
rect 329834 322980 329840 322992
rect 322532 322952 329840 322980
rect 322532 322940 322538 322952
rect 329834 322940 329840 322952
rect 329892 322940 329898 322992
rect 126882 322872 126888 322924
rect 126940 322912 126946 322924
rect 134058 322912 134064 322924
rect 126940 322884 134064 322912
rect 126940 322872 126946 322884
rect 134058 322872 134064 322884
rect 134116 322912 134122 322924
rect 197354 322912 197360 322924
rect 134116 322884 197360 322912
rect 134116 322872 134122 322884
rect 197354 322872 197360 322884
rect 197412 322872 197418 322924
rect 75270 322396 75276 322448
rect 75328 322436 75334 322448
rect 124306 322436 124312 322448
rect 75328 322408 124312 322436
rect 75328 322396 75334 322408
rect 124306 322396 124312 322408
rect 124364 322396 124370 322448
rect 50798 322328 50804 322380
rect 50856 322368 50862 322380
rect 107470 322368 107476 322380
rect 50856 322340 107476 322368
rect 50856 322328 50862 322340
rect 107470 322328 107476 322340
rect 107528 322328 107534 322380
rect 54938 322260 54944 322312
rect 54996 322300 55002 322312
rect 131114 322300 131120 322312
rect 54996 322272 131120 322300
rect 54996 322260 55002 322272
rect 131114 322260 131120 322272
rect 131172 322260 131178 322312
rect 95326 322192 95332 322244
rect 95384 322232 95390 322244
rect 174630 322232 174636 322244
rect 95384 322204 174636 322232
rect 95384 322192 95390 322204
rect 174630 322192 174636 322204
rect 174688 322192 174694 322244
rect 131114 321580 131120 321632
rect 131172 321620 131178 321632
rect 170490 321620 170496 321632
rect 131172 321592 170496 321620
rect 131172 321580 131178 321592
rect 170490 321580 170496 321592
rect 170548 321580 170554 321632
rect 80790 320832 80796 320884
rect 80848 320872 80854 320884
rect 191098 320872 191104 320884
rect 80848 320844 191104 320872
rect 80848 320832 80854 320844
rect 191098 320832 191104 320844
rect 191156 320832 191162 320884
rect 172422 320152 172428 320204
rect 172480 320192 172486 320204
rect 197354 320192 197360 320204
rect 172480 320164 197360 320192
rect 172480 320152 172486 320164
rect 197354 320152 197360 320164
rect 197412 320152 197418 320204
rect 71314 319472 71320 319524
rect 71372 319512 71378 319524
rect 135898 319512 135904 319524
rect 71372 319484 135904 319512
rect 71372 319472 71378 319484
rect 135898 319472 135904 319484
rect 135956 319472 135962 319524
rect 177942 319472 177948 319524
rect 178000 319512 178006 319524
rect 198182 319512 198188 319524
rect 178000 319484 198188 319512
rect 178000 319472 178006 319484
rect 198182 319472 198188 319484
rect 198240 319472 198246 319524
rect 101398 319404 101404 319456
rect 101456 319444 101462 319456
rect 181530 319444 181536 319456
rect 101456 319416 181536 319444
rect 101456 319404 101462 319416
rect 181530 319404 181536 319416
rect 181588 319404 181594 319456
rect 66162 318792 66168 318844
rect 66220 318832 66226 318844
rect 177942 318832 177948 318844
rect 66220 318804 177948 318832
rect 66220 318792 66226 318804
rect 177942 318792 177948 318804
rect 178000 318792 178006 318844
rect 322842 318792 322848 318844
rect 322900 318832 322906 318844
rect 323670 318832 323676 318844
rect 322900 318804 323676 318832
rect 322900 318792 322906 318804
rect 323670 318792 323676 318804
rect 323728 318792 323734 318844
rect 93210 318180 93216 318232
rect 93268 318220 93274 318232
rect 115382 318220 115388 318232
rect 93268 318192 115388 318220
rect 93268 318180 93274 318192
rect 115382 318180 115388 318192
rect 115440 318180 115446 318232
rect 84286 318112 84292 318164
rect 84344 318152 84350 318164
rect 113818 318152 113824 318164
rect 84344 318124 113824 318152
rect 84344 318112 84350 318124
rect 113818 318112 113824 318124
rect 113876 318112 113882 318164
rect 111242 318044 111248 318096
rect 111300 318084 111306 318096
rect 173158 318084 173164 318096
rect 111300 318056 173164 318084
rect 111300 318044 111306 318056
rect 173158 318044 173164 318056
rect 173216 318044 173222 318096
rect 115290 317432 115296 317484
rect 115348 317472 115354 317484
rect 197170 317472 197176 317484
rect 115348 317444 197176 317472
rect 115348 317432 115354 317444
rect 197170 317432 197176 317444
rect 197228 317472 197234 317484
rect 198642 317472 198648 317484
rect 197228 317444 198648 317472
rect 197228 317432 197234 317444
rect 198642 317432 198648 317444
rect 198700 317432 198706 317484
rect 102870 317364 102876 317416
rect 102928 317404 102934 317416
rect 129918 317404 129924 317416
rect 102928 317376 129924 317404
rect 102928 317364 102934 317376
rect 129918 317364 129924 317376
rect 129976 317364 129982 317416
rect 322474 317364 322480 317416
rect 322532 317404 322538 317416
rect 335538 317404 335544 317416
rect 322532 317376 335544 317404
rect 322532 317364 322538 317376
rect 335538 317364 335544 317376
rect 335596 317404 335602 317416
rect 336642 317404 336648 317416
rect 335596 317376 336648 317404
rect 335596 317364 335602 317376
rect 336642 317364 336648 317376
rect 336700 317364 336706 317416
rect 93946 316820 93952 316872
rect 94004 316860 94010 316872
rect 116670 316860 116676 316872
rect 94004 316832 116676 316860
rect 94004 316820 94010 316832
rect 116670 316820 116676 316832
rect 116728 316820 116734 316872
rect 75178 316752 75184 316804
rect 75236 316792 75242 316804
rect 142982 316792 142988 316804
rect 75236 316764 142988 316792
rect 75236 316752 75242 316764
rect 142982 316752 142988 316764
rect 143040 316752 143046 316804
rect 42610 316684 42616 316736
rect 42668 316724 42674 316736
rect 122834 316724 122840 316736
rect 42668 316696 122840 316724
rect 42668 316684 42674 316696
rect 122834 316684 122840 316696
rect 122892 316684 122898 316736
rect 130378 316684 130384 316736
rect 130436 316724 130442 316736
rect 167730 316724 167736 316736
rect 130436 316696 167736 316724
rect 130436 316684 130442 316696
rect 167730 316684 167736 316696
rect 167788 316684 167794 316736
rect 336642 316684 336648 316736
rect 336700 316724 336706 316736
rect 454678 316724 454684 316736
rect 336700 316696 454684 316724
rect 336700 316684 336706 316696
rect 454678 316684 454684 316696
rect 454736 316684 454742 316736
rect 130286 316004 130292 316056
rect 130344 316044 130350 316056
rect 181530 316044 181536 316056
rect 130344 316016 181536 316044
rect 130344 316004 130350 316016
rect 181530 316004 181536 316016
rect 181588 316004 181594 316056
rect 99282 315324 99288 315376
rect 99340 315364 99346 315376
rect 142430 315364 142436 315376
rect 99340 315336 142436 315364
rect 99340 315324 99346 315336
rect 142430 315324 142436 315336
rect 142488 315324 142494 315376
rect 75914 315256 75920 315308
rect 75972 315296 75978 315308
rect 133138 315296 133144 315308
rect 75972 315268 133144 315296
rect 75972 315256 75978 315268
rect 133138 315256 133144 315268
rect 133196 315256 133202 315308
rect 111058 314644 111064 314696
rect 111116 314684 111122 314696
rect 175182 314684 175188 314696
rect 111116 314656 175188 314684
rect 111116 314644 111122 314656
rect 175182 314644 175188 314656
rect 175240 314684 175246 314696
rect 197354 314684 197360 314696
rect 175240 314656 197360 314684
rect 175240 314644 175246 314656
rect 197354 314644 197360 314656
rect 197412 314644 197418 314696
rect 91002 314576 91008 314628
rect 91060 314616 91066 314628
rect 124306 314616 124312 314628
rect 91060 314588 124312 314616
rect 91060 314576 91066 314588
rect 124306 314576 124312 314588
rect 124364 314616 124370 314628
rect 125502 314616 125508 314628
rect 124364 314588 125508 314616
rect 124364 314576 124370 314588
rect 125502 314576 125508 314588
rect 125560 314576 125566 314628
rect 322474 314576 322480 314628
rect 322532 314616 322538 314628
rect 333974 314616 333980 314628
rect 322532 314588 333980 314616
rect 322532 314576 322538 314588
rect 333974 314576 333980 314588
rect 334032 314576 334038 314628
rect 76558 313964 76564 314016
rect 76616 314004 76622 314016
rect 176010 314004 176016 314016
rect 76616 313976 176016 314004
rect 76616 313964 76622 313976
rect 176010 313964 176016 313976
rect 176068 313964 176074 314016
rect 3418 313896 3424 313948
rect 3476 313936 3482 313948
rect 116670 313936 116676 313948
rect 3476 313908 116676 313936
rect 3476 313896 3482 313908
rect 116670 313896 116676 313908
rect 116728 313896 116734 313948
rect 333974 313896 333980 313948
rect 334032 313936 334038 313948
rect 500954 313936 500960 313948
rect 334032 313908 500960 313936
rect 334032 313896 334038 313908
rect 500954 313896 500960 313908
rect 501012 313896 501018 313948
rect 125502 313352 125508 313404
rect 125560 313392 125566 313404
rect 133966 313392 133972 313404
rect 125560 313364 133972 313392
rect 125560 313352 125566 313364
rect 133966 313352 133972 313364
rect 134024 313352 134030 313404
rect 83550 313284 83556 313336
rect 83608 313324 83614 313336
rect 108666 313324 108672 313336
rect 83608 313296 108672 313324
rect 83608 313284 83614 313296
rect 108666 313284 108672 313296
rect 108724 313284 108730 313336
rect 129182 313284 129188 313336
rect 129240 313324 129246 313336
rect 197354 313324 197360 313336
rect 129240 313296 197360 313324
rect 129240 313284 129246 313296
rect 197354 313284 197360 313296
rect 197412 313284 197418 313336
rect 108684 313256 108712 313284
rect 142154 313256 142160 313268
rect 108684 313228 142160 313256
rect 142154 313216 142160 313228
rect 142212 313256 142218 313268
rect 143442 313256 143448 313268
rect 142212 313228 143448 313256
rect 142212 313216 142218 313228
rect 143442 313216 143448 313228
rect 143500 313216 143506 313268
rect 86310 312604 86316 312656
rect 86368 312644 86374 312656
rect 116578 312644 116584 312656
rect 86368 312616 116584 312644
rect 86368 312604 86374 312616
rect 116578 312604 116584 312616
rect 116636 312604 116642 312656
rect 143442 312604 143448 312656
rect 143500 312644 143506 312656
rect 195422 312644 195428 312656
rect 143500 312616 195428 312644
rect 143500 312604 143506 312616
rect 195422 312604 195428 312616
rect 195480 312604 195486 312656
rect 72418 312536 72424 312588
rect 72476 312576 72482 312588
rect 149698 312576 149704 312588
rect 72476 312548 149704 312576
rect 72476 312536 72482 312548
rect 149698 312536 149704 312548
rect 149756 312536 149762 312588
rect 504358 312536 504364 312588
rect 504416 312576 504422 312588
rect 580258 312576 580264 312588
rect 504416 312548 580264 312576
rect 504416 312536 504422 312548
rect 580258 312536 580264 312548
rect 580316 312536 580322 312588
rect 322842 311992 322848 312044
rect 322900 312032 322906 312044
rect 324406 312032 324412 312044
rect 322900 312004 324412 312032
rect 322900 311992 322906 312004
rect 324406 311992 324412 312004
rect 324464 311992 324470 312044
rect 73890 311176 73896 311228
rect 73948 311216 73954 311228
rect 120074 311216 120080 311228
rect 73948 311188 120080 311216
rect 73948 311176 73954 311188
rect 120074 311176 120080 311188
rect 120132 311176 120138 311228
rect 45370 311108 45376 311160
rect 45428 311148 45434 311160
rect 176102 311148 176108 311160
rect 45428 311120 176108 311148
rect 45428 311108 45434 311120
rect 176102 311108 176108 311120
rect 176160 311108 176166 311160
rect 324406 311108 324412 311160
rect 324464 311148 324470 311160
rect 413278 311148 413284 311160
rect 324464 311120 413284 311148
rect 324464 311108 324470 311120
rect 413278 311108 413284 311120
rect 413336 311108 413342 311160
rect 89714 310496 89720 310548
rect 89772 310536 89778 310548
rect 190362 310536 190368 310548
rect 89772 310508 190368 310536
rect 89772 310496 89778 310508
rect 190362 310496 190368 310508
rect 190420 310536 190426 310548
rect 197354 310536 197360 310548
rect 190420 310508 197360 310536
rect 190420 310496 190426 310508
rect 197354 310496 197360 310508
rect 197412 310496 197418 310548
rect 100662 310428 100668 310480
rect 100720 310468 100726 310480
rect 103606 310468 103612 310480
rect 100720 310440 103612 310468
rect 100720 310428 100726 310440
rect 103606 310428 103612 310440
rect 103664 310428 103670 310480
rect 120074 310428 120080 310480
rect 120132 310468 120138 310480
rect 120810 310468 120816 310480
rect 120132 310440 120816 310468
rect 120132 310428 120138 310440
rect 120810 310428 120816 310440
rect 120868 310468 120874 310480
rect 195238 310468 195244 310480
rect 120868 310440 195244 310468
rect 120868 310428 120874 310440
rect 195238 310428 195244 310440
rect 195296 310428 195302 310480
rect 106090 309816 106096 309868
rect 106148 309856 106154 309868
rect 113818 309856 113824 309868
rect 106148 309828 113824 309856
rect 106148 309816 106154 309828
rect 113818 309816 113824 309828
rect 113876 309816 113882 309868
rect 89070 309748 89076 309800
rect 89128 309788 89134 309800
rect 142798 309788 142804 309800
rect 89128 309760 142804 309788
rect 89128 309748 89134 309760
rect 142798 309748 142804 309760
rect 142856 309748 142862 309800
rect 322474 309748 322480 309800
rect 322532 309788 322538 309800
rect 327074 309788 327080 309800
rect 322532 309760 327080 309788
rect 322532 309748 322538 309760
rect 327074 309748 327080 309760
rect 327132 309788 327138 309800
rect 377398 309788 377404 309800
rect 327132 309760 377404 309788
rect 327132 309748 327138 309760
rect 377398 309748 377404 309760
rect 377456 309748 377462 309800
rect 56318 309136 56324 309188
rect 56376 309176 56382 309188
rect 198090 309176 198096 309188
rect 56376 309148 198096 309176
rect 56376 309136 56382 309148
rect 198090 309136 198096 309148
rect 198148 309136 198154 309188
rect 195238 309068 195244 309120
rect 195296 309108 195302 309120
rect 195514 309108 195520 309120
rect 195296 309080 195520 309108
rect 195296 309068 195302 309080
rect 195514 309068 195520 309080
rect 195572 309068 195578 309120
rect 101950 308524 101956 308576
rect 102008 308564 102014 308576
rect 133138 308564 133144 308576
rect 102008 308536 133144 308564
rect 102008 308524 102014 308536
rect 133138 308524 133144 308536
rect 133196 308524 133202 308576
rect 106182 308456 106188 308508
rect 106240 308496 106246 308508
rect 138658 308496 138664 308508
rect 106240 308468 138664 308496
rect 106240 308456 106246 308468
rect 138658 308456 138664 308468
rect 138716 308456 138722 308508
rect 93118 308388 93124 308440
rect 93176 308428 93182 308440
rect 140130 308428 140136 308440
rect 93176 308400 140136 308428
rect 93176 308388 93182 308400
rect 140130 308388 140136 308400
rect 140188 308388 140194 308440
rect 68830 307776 68836 307828
rect 68888 307816 68894 307828
rect 195238 307816 195244 307828
rect 68888 307788 195244 307816
rect 68888 307776 68894 307788
rect 195238 307776 195244 307788
rect 195296 307776 195302 307828
rect 322474 307708 322480 307760
rect 322532 307748 322538 307760
rect 331214 307748 331220 307760
rect 322532 307720 331220 307748
rect 322532 307708 322538 307720
rect 331214 307708 331220 307720
rect 331272 307708 331278 307760
rect 104802 307096 104808 307148
rect 104860 307136 104866 307148
rect 145650 307136 145656 307148
rect 104860 307108 145656 307136
rect 104860 307096 104866 307108
rect 145650 307096 145656 307108
rect 145708 307096 145714 307148
rect 79410 307028 79416 307080
rect 79468 307068 79474 307080
rect 128998 307068 129004 307080
rect 79468 307040 129004 307068
rect 79468 307028 79474 307040
rect 128998 307028 129004 307040
rect 129056 307028 129062 307080
rect 331214 307028 331220 307080
rect 331272 307068 331278 307080
rect 447778 307068 447784 307080
rect 331272 307040 447784 307068
rect 331272 307028 331278 307040
rect 447778 307028 447784 307040
rect 447836 307028 447842 307080
rect 71038 306416 71044 306468
rect 71096 306456 71102 306468
rect 171778 306456 171784 306468
rect 71096 306428 171784 306456
rect 71096 306416 71102 306428
rect 171778 306416 171784 306428
rect 171836 306416 171842 306468
rect 182174 306388 182180 306400
rect 48286 306360 182180 306388
rect 48286 306332 48314 306360
rect 182174 306348 182180 306360
rect 182232 306348 182238 306400
rect 3418 306280 3424 306332
rect 3476 306320 3482 306332
rect 21358 306320 21364 306332
rect 3476 306292 21364 306320
rect 3476 306280 3482 306292
rect 21358 306280 21364 306292
rect 21416 306280 21422 306332
rect 41046 306280 41052 306332
rect 41104 306320 41110 306332
rect 48286 306320 48320 306332
rect 41104 306292 48320 306320
rect 41104 306280 41110 306292
rect 48314 306280 48320 306292
rect 48372 306280 48378 306332
rect 68738 305668 68744 305720
rect 68796 305708 68802 305720
rect 120074 305708 120080 305720
rect 68796 305680 120080 305708
rect 68796 305668 68802 305680
rect 120074 305668 120080 305680
rect 120132 305668 120138 305720
rect 83642 305600 83648 305652
rect 83700 305640 83706 305652
rect 148410 305640 148416 305652
rect 83700 305612 148416 305640
rect 83700 305600 83706 305612
rect 148410 305600 148416 305612
rect 148468 305600 148474 305652
rect 99374 304988 99380 305040
rect 99432 305028 99438 305040
rect 169110 305028 169116 305040
rect 99432 305000 169116 305028
rect 99432 304988 99438 305000
rect 169110 304988 169116 305000
rect 169168 304988 169174 305040
rect 322474 304988 322480 305040
rect 322532 305028 322538 305040
rect 327166 305028 327172 305040
rect 322532 305000 327172 305028
rect 322532 304988 322538 305000
rect 327166 304988 327172 305000
rect 327224 304988 327230 305040
rect 104158 304376 104164 304428
rect 104216 304416 104222 304428
rect 137370 304416 137376 304428
rect 104216 304388 137376 304416
rect 104216 304376 104222 304388
rect 137370 304376 137376 304388
rect 137428 304376 137434 304428
rect 90358 304308 90364 304360
rect 90416 304348 90422 304360
rect 129090 304348 129096 304360
rect 90416 304320 129096 304348
rect 90416 304308 90422 304320
rect 129090 304308 129096 304320
rect 129148 304308 129154 304360
rect 87598 304240 87604 304292
rect 87656 304280 87662 304292
rect 167730 304280 167736 304292
rect 87656 304252 167736 304280
rect 87656 304240 87662 304252
rect 167730 304240 167736 304252
rect 167788 304240 167794 304292
rect 56410 303696 56416 303748
rect 56468 303736 56474 303748
rect 117866 303736 117872 303748
rect 56468 303708 117872 303736
rect 56468 303696 56474 303708
rect 117866 303696 117872 303708
rect 117924 303696 117930 303748
rect 90266 303628 90272 303680
rect 90324 303668 90330 303680
rect 171962 303668 171968 303680
rect 90324 303640 171968 303668
rect 90324 303628 90330 303640
rect 171962 303628 171968 303640
rect 172020 303628 172026 303680
rect 187234 303628 187240 303680
rect 187292 303668 187298 303680
rect 197354 303668 197360 303680
rect 187292 303640 197360 303668
rect 187292 303628 187298 303640
rect 197354 303628 197360 303640
rect 197412 303628 197418 303680
rect 52362 302880 52368 302932
rect 52420 302920 52426 302932
rect 70486 302920 70492 302932
rect 52420 302892 70492 302920
rect 52420 302880 52426 302892
rect 70486 302880 70492 302892
rect 70544 302880 70550 302932
rect 97350 302880 97356 302932
rect 97408 302920 97414 302932
rect 196618 302920 196624 302932
rect 97408 302892 196624 302920
rect 97408 302880 97414 302892
rect 196618 302880 196624 302892
rect 196676 302880 196682 302932
rect 111150 302404 111156 302456
rect 111208 302444 111214 302456
rect 111610 302444 111616 302456
rect 111208 302416 111616 302444
rect 111208 302404 111214 302416
rect 111610 302404 111616 302416
rect 111668 302444 111674 302456
rect 158070 302444 158076 302456
rect 111668 302416 158076 302444
rect 111668 302404 111674 302416
rect 158070 302404 158076 302416
rect 158128 302404 158134 302456
rect 87598 302336 87604 302388
rect 87656 302376 87662 302388
rect 138750 302376 138756 302388
rect 87656 302348 138756 302376
rect 87656 302336 87662 302348
rect 138750 302336 138756 302348
rect 138808 302336 138814 302388
rect 79134 302268 79140 302320
rect 79192 302308 79198 302320
rect 142890 302308 142896 302320
rect 79192 302280 142896 302308
rect 79192 302268 79198 302280
rect 142890 302268 142896 302280
rect 142948 302268 142954 302320
rect 67358 302200 67364 302252
rect 67416 302240 67422 302252
rect 193122 302240 193128 302252
rect 67416 302212 193128 302240
rect 67416 302200 67422 302212
rect 193122 302200 193128 302212
rect 193180 302240 193186 302252
rect 197354 302240 197360 302252
rect 193180 302212 197360 302240
rect 193180 302200 193186 302212
rect 197354 302200 197360 302212
rect 197412 302200 197418 302252
rect 322474 302200 322480 302252
rect 322532 302240 322538 302252
rect 327074 302240 327080 302252
rect 322532 302212 327080 302240
rect 322532 302200 322538 302212
rect 327074 302200 327080 302212
rect 327132 302200 327138 302252
rect 98546 301588 98552 301640
rect 98604 301628 98610 301640
rect 111058 301628 111064 301640
rect 98604 301600 111064 301628
rect 98604 301588 98610 301600
rect 111058 301588 111064 301600
rect 111116 301588 111122 301640
rect 82078 301520 82084 301572
rect 82136 301560 82142 301572
rect 147030 301560 147036 301572
rect 82136 301532 147036 301560
rect 82136 301520 82142 301532
rect 147030 301520 147036 301532
rect 147088 301520 147094 301572
rect 322198 301520 322204 301572
rect 322256 301560 322262 301572
rect 333974 301560 333980 301572
rect 322256 301532 333980 301560
rect 322256 301520 322262 301532
rect 333974 301520 333980 301532
rect 334032 301520 334038 301572
rect 53650 301452 53656 301504
rect 53708 301492 53714 301504
rect 132586 301492 132592 301504
rect 53708 301464 132592 301492
rect 53708 301452 53714 301464
rect 132586 301452 132592 301464
rect 132644 301452 132650 301504
rect 175090 301452 175096 301504
rect 175148 301492 175154 301504
rect 197262 301492 197268 301504
rect 175148 301464 197268 301492
rect 175148 301452 175154 301464
rect 197262 301452 197268 301464
rect 197320 301452 197326 301504
rect 322842 301452 322848 301504
rect 322900 301492 322906 301504
rect 325050 301492 325056 301504
rect 322900 301464 325056 301492
rect 322900 301452 322906 301464
rect 325050 301452 325056 301464
rect 325108 301492 325114 301504
rect 429194 301492 429200 301504
rect 325108 301464 429200 301492
rect 325108 301452 325114 301464
rect 429194 301452 429200 301464
rect 429252 301452 429258 301504
rect 125778 300976 125784 301028
rect 125836 301016 125842 301028
rect 126238 301016 126244 301028
rect 125836 300988 126244 301016
rect 125836 300976 125842 300988
rect 126238 300976 126244 300988
rect 126296 301016 126302 301028
rect 152550 301016 152556 301028
rect 126296 300988 152556 301016
rect 126296 300976 126302 300988
rect 152550 300976 152556 300988
rect 152608 300976 152614 301028
rect 109678 300908 109684 300960
rect 109736 300948 109742 300960
rect 110322 300948 110328 300960
rect 109736 300920 110328 300948
rect 109736 300908 109742 300920
rect 110322 300908 110328 300920
rect 110380 300948 110386 300960
rect 175090 300948 175096 300960
rect 110380 300920 175096 300948
rect 110380 300908 110386 300920
rect 175090 300908 175096 300920
rect 175148 300908 175154 300960
rect 84194 300840 84200 300892
rect 84252 300880 84258 300892
rect 166258 300880 166264 300892
rect 84252 300852 166264 300880
rect 84252 300840 84258 300852
rect 166258 300840 166264 300852
rect 166316 300840 166322 300892
rect 333974 300840 333980 300892
rect 334032 300880 334038 300892
rect 468478 300880 468484 300892
rect 334032 300852 468484 300880
rect 334032 300840 334038 300852
rect 468478 300840 468484 300852
rect 468536 300840 468542 300892
rect 117866 300772 117872 300824
rect 117924 300812 117930 300824
rect 132770 300812 132776 300824
rect 117924 300784 132776 300812
rect 117924 300772 117930 300784
rect 132770 300772 132776 300784
rect 132828 300812 132834 300824
rect 133782 300812 133788 300824
rect 132828 300784 133788 300812
rect 132828 300772 132834 300784
rect 133782 300772 133788 300784
rect 133840 300772 133846 300824
rect 182174 300772 182180 300824
rect 182232 300812 182238 300824
rect 183462 300812 183468 300824
rect 182232 300784 183468 300812
rect 182232 300772 182238 300784
rect 183462 300772 183468 300784
rect 183520 300772 183526 300824
rect 148502 300268 148508 300280
rect 132466 300240 148508 300268
rect 117958 300160 117964 300212
rect 118016 300200 118022 300212
rect 125778 300200 125784 300212
rect 118016 300172 125784 300200
rect 118016 300160 118022 300172
rect 125778 300160 125784 300172
rect 125836 300160 125842 300212
rect 104986 300092 104992 300144
rect 105044 300132 105050 300144
rect 127158 300132 127164 300144
rect 105044 300104 127164 300132
rect 105044 300092 105050 300104
rect 127158 300092 127164 300104
rect 127216 300132 127222 300144
rect 132466 300132 132494 300240
rect 148502 300228 148508 300240
rect 148560 300228 148566 300280
rect 133782 300160 133788 300212
rect 133840 300200 133846 300212
rect 155310 300200 155316 300212
rect 133840 300172 155316 300200
rect 133840 300160 133846 300172
rect 155310 300160 155316 300172
rect 155368 300160 155374 300212
rect 127216 300104 132494 300132
rect 127216 300092 127222 300104
rect 138014 300092 138020 300144
rect 138072 300132 138078 300144
rect 163590 300132 163596 300144
rect 138072 300104 163596 300132
rect 138072 300092 138078 300104
rect 163590 300092 163596 300104
rect 163648 300092 163654 300144
rect 183462 300092 183468 300144
rect 183520 300132 183526 300144
rect 197354 300132 197360 300144
rect 183520 300104 197360 300132
rect 183520 300092 183526 300104
rect 197354 300092 197360 300104
rect 197412 300092 197418 300144
rect 335262 300092 335268 300144
rect 335320 300132 335326 300144
rect 580350 300132 580356 300144
rect 335320 300104 580356 300132
rect 335320 300092 335326 300104
rect 580350 300092 580356 300104
rect 580408 300092 580414 300144
rect 87506 299684 87512 299736
rect 87564 299724 87570 299736
rect 135990 299724 135996 299736
rect 87564 299696 135996 299724
rect 87564 299684 87570 299696
rect 135990 299684 135996 299696
rect 136048 299684 136054 299736
rect 102134 299616 102140 299668
rect 102192 299656 102198 299668
rect 184290 299656 184296 299668
rect 102192 299628 184296 299656
rect 102192 299616 102198 299628
rect 184290 299616 184296 299628
rect 184348 299616 184354 299668
rect 22738 299548 22744 299600
rect 22796 299588 22802 299600
rect 117958 299588 117964 299600
rect 22796 299560 117964 299588
rect 22796 299548 22802 299560
rect 117958 299548 117964 299560
rect 118016 299548 118022 299600
rect 69014 299480 69020 299532
rect 69072 299520 69078 299532
rect 166442 299520 166448 299532
rect 69072 299492 166448 299520
rect 69072 299480 69078 299492
rect 166442 299480 166448 299492
rect 166500 299480 166506 299532
rect 65518 299412 65524 299464
rect 65576 299452 65582 299464
rect 68646 299452 68652 299464
rect 65576 299424 68652 299452
rect 65576 299412 65582 299424
rect 68646 299412 68652 299424
rect 68704 299412 68710 299464
rect 83458 298732 83464 298784
rect 83516 298772 83522 298784
rect 129918 298772 129924 298784
rect 83516 298744 129924 298772
rect 83516 298732 83522 298744
rect 129918 298732 129924 298744
rect 129976 298732 129982 298784
rect 322474 298732 322480 298784
rect 322532 298772 322538 298784
rect 330478 298772 330484 298784
rect 322532 298744 330484 298772
rect 322532 298732 322538 298744
rect 330478 298732 330484 298744
rect 330536 298732 330542 298784
rect 113818 298392 113824 298444
rect 113876 298432 113882 298444
rect 156690 298432 156696 298444
rect 113876 298404 156696 298432
rect 113876 298392 113882 298404
rect 156690 298392 156696 298404
rect 156748 298392 156754 298444
rect 82262 298324 82268 298376
rect 82320 298364 82326 298376
rect 134610 298364 134616 298376
rect 82320 298336 134616 298364
rect 82320 298324 82326 298336
rect 134610 298324 134616 298336
rect 134668 298324 134674 298376
rect 68646 298256 68652 298308
rect 68704 298296 68710 298308
rect 159634 298296 159640 298308
rect 68704 298268 159640 298296
rect 68704 298256 68710 298268
rect 159634 298256 159640 298268
rect 159692 298256 159698 298308
rect 93854 298188 93860 298240
rect 93912 298228 93918 298240
rect 196710 298228 196716 298240
rect 93912 298200 196716 298228
rect 93912 298188 93918 298200
rect 196710 298188 196716 298200
rect 196768 298188 196774 298240
rect 69106 298120 69112 298172
rect 69164 298160 69170 298172
rect 187234 298160 187240 298172
rect 69164 298132 187240 298160
rect 69164 298120 69170 298132
rect 187234 298120 187240 298132
rect 187292 298120 187298 298172
rect 57238 297480 57244 297492
rect 45526 297452 57244 297480
rect 17218 297372 17224 297424
rect 17276 297412 17282 297424
rect 45526 297412 45554 297452
rect 57238 297440 57244 297452
rect 57296 297480 57302 297492
rect 97074 297480 97080 297492
rect 57296 297452 97080 297480
rect 57296 297440 57302 297452
rect 97074 297440 97080 297452
rect 97132 297440 97138 297492
rect 17276 297384 45554 297412
rect 17276 297372 17282 297384
rect 74994 297372 75000 297424
rect 75052 297412 75058 297424
rect 147858 297412 147864 297424
rect 75052 297384 147864 297412
rect 75052 297372 75058 297384
rect 147858 297372 147864 297384
rect 147916 297412 147922 297424
rect 148134 297412 148140 297424
rect 147916 297384 148140 297412
rect 147916 297372 147922 297384
rect 148134 297372 148140 297384
rect 148192 297372 148198 297424
rect 330478 297372 330484 297424
rect 330536 297412 330542 297424
rect 353386 297412 353392 297424
rect 330536 297384 353392 297412
rect 330536 297372 330542 297384
rect 353386 297372 353392 297384
rect 353444 297412 353450 297424
rect 407758 297412 407764 297424
rect 353444 297384 407764 297412
rect 353444 297372 353450 297384
rect 407758 297372 407764 297384
rect 407816 297372 407822 297424
rect 193030 297168 193036 297220
rect 193088 297208 193094 297220
rect 197354 297208 197360 297220
rect 193088 297180 197360 297208
rect 193088 297168 193094 297180
rect 197354 297168 197360 297180
rect 197412 297168 197418 297220
rect 107286 296964 107292 297016
rect 107344 297004 107350 297016
rect 123754 297004 123760 297016
rect 107344 296976 123760 297004
rect 107344 296964 107350 296976
rect 123754 296964 123760 296976
rect 123812 296964 123818 297016
rect 102870 296896 102876 296948
rect 102928 296936 102934 296948
rect 145558 296936 145564 296948
rect 102928 296908 145564 296936
rect 102928 296896 102934 296908
rect 145558 296896 145564 296908
rect 145616 296896 145622 296948
rect 148134 296896 148140 296948
rect 148192 296936 148198 296948
rect 152458 296936 152464 296948
rect 148192 296908 152464 296936
rect 148192 296896 148198 296908
rect 152458 296896 152464 296908
rect 152516 296896 152522 296948
rect 116670 296828 116676 296880
rect 116728 296868 116734 296880
rect 159542 296868 159548 296880
rect 116728 296840 159548 296868
rect 116728 296828 116734 296840
rect 159542 296828 159548 296840
rect 159600 296828 159606 296880
rect 97074 296760 97080 296812
rect 97132 296800 97138 296812
rect 160830 296800 160836 296812
rect 97132 296772 160836 296800
rect 97132 296760 97138 296772
rect 160830 296760 160836 296772
rect 160888 296760 160894 296812
rect 76466 296692 76472 296744
rect 76524 296732 76530 296744
rect 182910 296732 182916 296744
rect 76524 296704 182916 296732
rect 76524 296692 76530 296704
rect 182910 296692 182916 296704
rect 182968 296692 182974 296744
rect 54754 295944 54760 295996
rect 54812 295984 54818 295996
rect 71774 295984 71780 295996
rect 54812 295956 71780 295984
rect 54812 295944 54818 295956
rect 71774 295944 71780 295956
rect 71832 295944 71838 295996
rect 114462 295944 114468 295996
rect 114520 295984 114526 295996
rect 115290 295984 115296 295996
rect 114520 295956 115296 295984
rect 114520 295944 114526 295956
rect 115290 295944 115296 295956
rect 115348 295944 115354 295996
rect 65978 295672 65984 295724
rect 66036 295712 66042 295724
rect 196618 295712 196624 295724
rect 66036 295684 196624 295712
rect 66036 295672 66042 295684
rect 196618 295672 196624 295684
rect 196676 295672 196682 295724
rect 83550 295604 83556 295656
rect 83608 295644 83614 295656
rect 133230 295644 133236 295656
rect 83608 295616 133236 295644
rect 83608 295604 83614 295616
rect 133230 295604 133236 295616
rect 133288 295604 133294 295656
rect 68922 295536 68928 295588
rect 68980 295576 68986 295588
rect 125042 295576 125048 295588
rect 68980 295548 125048 295576
rect 68980 295536 68986 295548
rect 125042 295536 125048 295548
rect 125100 295536 125106 295588
rect 93210 295468 93216 295520
rect 93268 295508 93274 295520
rect 188430 295508 188436 295520
rect 93268 295480 188436 295508
rect 93268 295468 93274 295480
rect 188430 295468 188436 295480
rect 188488 295468 188494 295520
rect 69198 295400 69204 295452
rect 69256 295440 69262 295452
rect 195882 295440 195888 295452
rect 69256 295412 195888 295440
rect 69256 295400 69262 295412
rect 195882 295400 195888 295412
rect 195940 295440 195946 295452
rect 197446 295440 197452 295452
rect 195940 295412 197452 295440
rect 195940 295400 195946 295412
rect 197446 295400 197452 295412
rect 197504 295400 197510 295452
rect 117222 295332 117228 295384
rect 117280 295372 117286 295384
rect 124858 295372 124864 295384
rect 117280 295344 124864 295372
rect 117280 295332 117286 295344
rect 124858 295332 124864 295344
rect 124916 295332 124922 295384
rect 322474 295332 322480 295384
rect 322532 295372 322538 295384
rect 331214 295372 331220 295384
rect 322532 295344 331220 295372
rect 322532 295332 322538 295344
rect 331214 295332 331220 295344
rect 331272 295332 331278 295384
rect 80330 295264 80336 295316
rect 80388 295304 80394 295316
rect 86218 295304 86224 295316
rect 80388 295276 86224 295304
rect 80388 295264 80394 295276
rect 86218 295264 86224 295276
rect 86276 295264 86282 295316
rect 117038 295264 117044 295316
rect 117096 295304 117102 295316
rect 123478 295304 123484 295316
rect 117096 295276 123484 295304
rect 117096 295264 117102 295276
rect 123478 295264 123484 295276
rect 123536 295264 123542 295316
rect 111242 294924 111248 294976
rect 111300 294964 111306 294976
rect 124950 294964 124956 294976
rect 111300 294936 124956 294964
rect 111300 294924 111306 294936
rect 124950 294924 124956 294936
rect 125008 294924 125014 294976
rect 84838 294856 84844 294908
rect 84896 294896 84902 294908
rect 91738 294896 91744 294908
rect 84896 294868 91744 294896
rect 84896 294856 84902 294868
rect 91738 294856 91744 294868
rect 91796 294856 91802 294908
rect 94498 294856 94504 294908
rect 94556 294896 94562 294908
rect 111150 294896 111156 294908
rect 94556 294868 111156 294896
rect 94556 294856 94562 294868
rect 111150 294856 111156 294868
rect 111208 294856 111214 294908
rect 106734 294788 106740 294840
rect 106792 294828 106798 294840
rect 126330 294828 126336 294840
rect 106792 294800 126336 294828
rect 106792 294788 106798 294800
rect 126330 294788 126336 294800
rect 126388 294788 126394 294840
rect 82906 294720 82912 294772
rect 82964 294760 82970 294772
rect 107286 294760 107292 294772
rect 82964 294732 107292 294760
rect 82964 294720 82970 294732
rect 107286 294720 107292 294732
rect 107344 294720 107350 294772
rect 119614 294720 119620 294772
rect 119672 294760 119678 294772
rect 147766 294760 147772 294772
rect 119672 294732 147772 294760
rect 119672 294720 119678 294732
rect 147766 294720 147772 294732
rect 147824 294720 147830 294772
rect 71314 294652 71320 294704
rect 71372 294692 71378 294704
rect 83458 294692 83464 294704
rect 71372 294664 83464 294692
rect 71372 294652 71378 294664
rect 83458 294652 83464 294664
rect 83516 294652 83522 294704
rect 87414 294652 87420 294704
rect 87472 294692 87478 294704
rect 117222 294692 117228 294704
rect 87472 294664 117228 294692
rect 87472 294652 87478 294664
rect 117222 294652 117228 294664
rect 117280 294652 117286 294704
rect 117682 294652 117688 294704
rect 117740 294692 117746 294704
rect 173250 294692 173256 294704
rect 117740 294664 173256 294692
rect 117740 294652 117746 294664
rect 173250 294652 173256 294664
rect 173308 294652 173314 294704
rect 71958 294584 71964 294636
rect 72016 294624 72022 294636
rect 101398 294624 101404 294636
rect 72016 294596 101404 294624
rect 72016 294584 72022 294596
rect 101398 294584 101404 294596
rect 101456 294584 101462 294636
rect 113818 294584 113824 294636
rect 113876 294624 113882 294636
rect 195330 294624 195336 294636
rect 113876 294596 195336 294624
rect 113876 294584 113882 294596
rect 195330 294584 195336 294596
rect 195388 294584 195394 294636
rect 72602 294516 72608 294568
rect 72660 294556 72666 294568
rect 74994 294556 75000 294568
rect 72660 294528 75000 294556
rect 72660 294516 72666 294528
rect 74994 294516 75000 294528
rect 75052 294516 75058 294568
rect 104894 294312 104900 294364
rect 104952 294352 104958 294364
rect 105814 294352 105820 294364
rect 104952 294324 105820 294352
rect 104952 294312 104958 294324
rect 105814 294312 105820 294324
rect 105872 294312 105878 294364
rect 107654 294312 107660 294364
rect 107712 294352 107718 294364
rect 108390 294352 108396 294364
rect 107712 294324 108396 294352
rect 107712 294312 107718 294324
rect 108390 294312 108396 294324
rect 108448 294312 108454 294364
rect 109310 294312 109316 294364
rect 109368 294352 109374 294364
rect 112438 294352 112444 294364
rect 109368 294324 112444 294352
rect 109368 294312 109374 294324
rect 112438 294312 112444 294324
rect 112496 294312 112502 294364
rect 79042 294176 79048 294228
rect 79100 294216 79106 294228
rect 79226 294216 79232 294228
rect 79100 294188 79232 294216
rect 79100 294176 79106 294188
rect 79226 294176 79232 294188
rect 79284 294176 79290 294228
rect 49602 294108 49608 294160
rect 49660 294148 49666 294160
rect 75178 294148 75184 294160
rect 49660 294120 75184 294148
rect 49660 294108 49666 294120
rect 75178 294108 75184 294120
rect 75236 294108 75242 294160
rect 86126 294108 86132 294160
rect 86184 294148 86190 294160
rect 87598 294148 87604 294160
rect 86184 294120 87604 294148
rect 86184 294108 86190 294120
rect 87598 294108 87604 294120
rect 87656 294108 87662 294160
rect 41230 294040 41236 294092
rect 41288 294080 41294 294092
rect 74534 294080 74540 294092
rect 41288 294052 74540 294080
rect 41288 294040 41294 294052
rect 74534 294040 74540 294052
rect 74592 294040 74598 294092
rect 99282 294040 99288 294092
rect 99340 294080 99346 294092
rect 101582 294080 101588 294092
rect 99340 294052 101588 294080
rect 99340 294040 99346 294052
rect 101582 294040 101588 294052
rect 101640 294040 101646 294092
rect 33778 293972 33784 294024
rect 33836 294012 33842 294024
rect 79042 294012 79048 294024
rect 33836 293984 79048 294012
rect 33836 293972 33842 293984
rect 79042 293972 79048 293984
rect 79100 293972 79106 294024
rect 100938 293972 100944 294024
rect 100996 294012 101002 294024
rect 118694 294012 118700 294024
rect 100996 293984 118700 294012
rect 100996 293972 101002 293984
rect 118694 293972 118700 293984
rect 118752 293972 118758 294024
rect 3418 293836 3424 293888
rect 3476 293876 3482 293888
rect 7558 293876 7564 293888
rect 3476 293848 7564 293876
rect 3476 293836 3482 293848
rect 7558 293836 7564 293848
rect 7616 293836 7622 293888
rect 41322 293224 41328 293276
rect 41380 293264 41386 293276
rect 99282 293264 99288 293276
rect 41380 293236 99288 293264
rect 41380 293224 41386 293236
rect 99282 293224 99288 293236
rect 99340 293224 99346 293276
rect 111702 293224 111708 293276
rect 111760 293264 111766 293276
rect 148318 293264 148324 293276
rect 111760 293236 148324 293264
rect 111760 293224 111766 293236
rect 148318 293224 148324 293236
rect 148376 293224 148382 293276
rect 322842 293224 322848 293276
rect 322900 293264 322906 293276
rect 324314 293264 324320 293276
rect 322900 293236 324320 293264
rect 322900 293224 322906 293236
rect 324314 293224 324320 293236
rect 324372 293264 324378 293276
rect 370498 293264 370504 293276
rect 324372 293236 370504 293264
rect 324372 293224 324378 293236
rect 370498 293224 370504 293236
rect 370556 293224 370562 293276
rect 91922 292816 91928 292868
rect 91980 292856 91986 292868
rect 117498 292856 117504 292868
rect 91980 292828 117504 292856
rect 91980 292816 91986 292828
rect 117498 292816 117504 292828
rect 117556 292816 117562 292868
rect 115198 292748 115204 292800
rect 115256 292788 115262 292800
rect 115750 292788 115756 292800
rect 115256 292760 115756 292788
rect 115256 292748 115262 292760
rect 115750 292748 115756 292760
rect 115808 292788 115814 292800
rect 155402 292788 155408 292800
rect 115808 292760 155408 292788
rect 115808 292748 115814 292760
rect 155402 292748 155408 292760
rect 155460 292748 155466 292800
rect 53098 292680 53104 292732
rect 53156 292720 53162 292732
rect 92566 292720 92572 292732
rect 53156 292692 92572 292720
rect 53156 292680 53162 292692
rect 92566 292680 92572 292692
rect 92624 292720 92630 292732
rect 92934 292720 92940 292732
rect 92624 292692 92940 292720
rect 92624 292680 92630 292692
rect 92934 292680 92940 292692
rect 92992 292680 92998 292732
rect 107378 292680 107384 292732
rect 107436 292720 107442 292732
rect 107562 292720 107568 292732
rect 107436 292692 107568 292720
rect 107436 292680 107442 292692
rect 107562 292680 107568 292692
rect 107620 292720 107626 292732
rect 151354 292720 151360 292732
rect 107620 292692 151360 292720
rect 107620 292680 107626 292692
rect 151354 292680 151360 292692
rect 151412 292680 151418 292732
rect 68738 292612 68744 292664
rect 68796 292652 68802 292664
rect 73798 292652 73804 292664
rect 68796 292624 73804 292652
rect 68796 292612 68802 292624
rect 73798 292612 73804 292624
rect 73856 292612 73862 292664
rect 73890 292612 73896 292664
rect 73948 292652 73954 292664
rect 124122 292652 124128 292664
rect 73948 292624 124128 292652
rect 73948 292612 73954 292624
rect 124122 292612 124128 292624
rect 124180 292612 124186 292664
rect 153470 292612 153476 292664
rect 153528 292652 153534 292664
rect 154666 292652 154672 292664
rect 153528 292624 154672 292652
rect 153528 292612 153534 292624
rect 154666 292612 154672 292624
rect 154724 292612 154730 292664
rect 8202 292544 8208 292596
rect 8260 292584 8266 292596
rect 96430 292584 96436 292596
rect 8260 292556 96436 292584
rect 8260 292544 8266 292556
rect 96430 292544 96436 292556
rect 96488 292544 96494 292596
rect 98362 292544 98368 292596
rect 98420 292584 98426 292596
rect 98730 292584 98736 292596
rect 98420 292556 98736 292584
rect 98420 292544 98426 292556
rect 98730 292544 98736 292556
rect 98788 292584 98794 292596
rect 189810 292584 189816 292596
rect 98788 292556 189816 292584
rect 98788 292544 98794 292556
rect 189810 292544 189816 292556
rect 189868 292544 189874 292596
rect 194042 292544 194048 292596
rect 194100 292584 194106 292596
rect 197446 292584 197452 292596
rect 194100 292556 197452 292584
rect 194100 292544 194106 292556
rect 197446 292544 197452 292556
rect 197504 292544 197510 292596
rect 124122 292476 124128 292528
rect 124180 292516 124186 292528
rect 129826 292516 129832 292528
rect 124180 292488 129832 292516
rect 124180 292476 124186 292488
rect 129826 292476 129832 292488
rect 129884 292476 129890 292528
rect 71682 292340 71688 292392
rect 71740 292380 71746 292392
rect 75362 292380 75368 292392
rect 71740 292352 75368 292380
rect 71740 292340 71746 292352
rect 75362 292340 75368 292352
rect 75420 292340 75426 292392
rect 121454 291932 121460 291984
rect 121512 291972 121518 291984
rect 153470 291972 153476 291984
rect 121512 291944 153476 291972
rect 121512 291932 121518 291944
rect 153470 291932 153476 291944
rect 153528 291972 153534 291984
rect 153930 291972 153936 291984
rect 153528 291944 153936 291972
rect 153528 291932 153534 291944
rect 153930 291932 153936 291944
rect 153988 291932 153994 291984
rect 71038 291904 71044 291916
rect 64846 291876 71044 291904
rect 61838 291796 61844 291848
rect 61896 291836 61902 291848
rect 64846 291836 64874 291876
rect 71038 291864 71044 291876
rect 71096 291864 71102 291916
rect 110874 291864 110880 291916
rect 110932 291864 110938 291916
rect 112806 291864 112812 291916
rect 112864 291904 112870 291916
rect 112864 291876 113174 291904
rect 112864 291864 112870 291876
rect 61896 291808 64874 291836
rect 61896 291796 61902 291808
rect 110892 291224 110920 291864
rect 113146 291292 113174 291876
rect 117498 291864 117504 291916
rect 117556 291864 117562 291916
rect 118694 291864 118700 291916
rect 118752 291904 118758 291916
rect 151170 291904 151176 291916
rect 118752 291876 151176 291904
rect 118752 291864 118758 291876
rect 151170 291864 151176 291876
rect 151228 291864 151234 291916
rect 117516 291836 117544 291864
rect 177390 291836 177396 291848
rect 117516 291808 177396 291836
rect 177390 291796 177396 291808
rect 177448 291796 177454 291848
rect 123662 291292 123668 291304
rect 113146 291264 123668 291292
rect 123662 291252 123668 291264
rect 123720 291252 123726 291304
rect 188522 291224 188528 291236
rect 110892 291196 188528 291224
rect 188522 291184 188528 291196
rect 188580 291184 188586 291236
rect 322842 291184 322848 291236
rect 322900 291224 322906 291236
rect 324314 291224 324320 291236
rect 322900 291196 324320 291224
rect 322900 291184 322906 291196
rect 324314 291184 324320 291196
rect 324372 291224 324378 291236
rect 499666 291224 499672 291236
rect 324372 291196 499672 291224
rect 324372 291184 324378 291196
rect 499666 291184 499672 291196
rect 499724 291184 499730 291236
rect 38102 291116 38108 291168
rect 38160 291156 38166 291168
rect 38470 291156 38476 291168
rect 38160 291128 38476 291156
rect 38160 291116 38166 291128
rect 38470 291116 38476 291128
rect 38528 291156 38534 291168
rect 67634 291156 67640 291168
rect 38528 291128 67640 291156
rect 38528 291116 38534 291128
rect 67634 291116 67640 291128
rect 67692 291116 67698 291168
rect 148410 291116 148416 291168
rect 148468 291156 148474 291168
rect 148594 291156 148600 291168
rect 148468 291128 148600 291156
rect 148468 291116 148474 291128
rect 148594 291116 148600 291128
rect 148652 291116 148658 291168
rect 25498 290436 25504 290488
rect 25556 290476 25562 290488
rect 38102 290476 38108 290488
rect 25556 290448 38108 290476
rect 25556 290436 25562 290448
rect 38102 290436 38108 290448
rect 38160 290436 38166 290488
rect 325050 290436 325056 290488
rect 325108 290476 325114 290488
rect 420914 290476 420920 290488
rect 325108 290448 420920 290476
rect 325108 290436 325114 290448
rect 420914 290436 420920 290448
rect 420972 290436 420978 290488
rect 148594 289960 148600 290012
rect 148652 290000 148658 290012
rect 179230 290000 179236 290012
rect 148652 289972 179236 290000
rect 148652 289960 148658 289972
rect 179230 289960 179236 289972
rect 179288 290000 179294 290012
rect 179288 289972 180794 290000
rect 179288 289960 179294 289972
rect 121546 289892 121552 289944
rect 121604 289932 121610 289944
rect 156598 289932 156604 289944
rect 121604 289904 156604 289932
rect 121604 289892 121610 289904
rect 156598 289892 156604 289904
rect 156656 289892 156662 289944
rect 59078 289824 59084 289876
rect 59136 289864 59142 289876
rect 67634 289864 67640 289876
rect 59136 289836 67640 289864
rect 59136 289824 59142 289836
rect 67634 289824 67640 289836
rect 67692 289824 67698 289876
rect 121454 289824 121460 289876
rect 121512 289864 121518 289876
rect 169202 289864 169208 289876
rect 121512 289836 169208 289864
rect 121512 289824 121518 289836
rect 169202 289824 169208 289836
rect 169260 289824 169266 289876
rect 180766 289864 180794 289972
rect 197446 289864 197452 289876
rect 180766 289836 197452 289864
rect 197446 289824 197452 289836
rect 197504 289824 197510 289876
rect 121546 289756 121552 289808
rect 121604 289796 121610 289808
rect 187050 289796 187056 289808
rect 121604 289768 187056 289796
rect 121604 289756 121610 289768
rect 187050 289756 187056 289768
rect 187108 289756 187114 289808
rect 69014 289144 69020 289196
rect 69072 289184 69078 289196
rect 69750 289184 69756 289196
rect 69072 289156 69756 289184
rect 69072 289144 69078 289156
rect 69750 289144 69756 289156
rect 69808 289144 69814 289196
rect 123570 289144 123576 289196
rect 123628 289184 123634 289196
rect 126422 289184 126428 289196
rect 123628 289156 126428 289184
rect 123628 289144 123634 289156
rect 126422 289144 126428 289156
rect 126480 289184 126486 289196
rect 168282 289184 168288 289196
rect 126480 289156 168288 289184
rect 126480 289144 126486 289156
rect 168282 289144 168288 289156
rect 168340 289144 168346 289196
rect 123662 289076 123668 289128
rect 123720 289116 123726 289128
rect 185762 289116 185768 289128
rect 123720 289088 185768 289116
rect 123720 289076 123726 289088
rect 185762 289076 185768 289088
rect 185820 289076 185826 289128
rect 60366 288396 60372 288448
rect 60424 288436 60430 288448
rect 67634 288436 67640 288448
rect 60424 288408 67640 288436
rect 60424 288396 60430 288408
rect 67634 288396 67640 288408
rect 67692 288396 67698 288448
rect 168282 288396 168288 288448
rect 168340 288436 168346 288448
rect 197446 288436 197452 288448
rect 168340 288408 197452 288436
rect 168340 288396 168346 288408
rect 197446 288396 197452 288408
rect 197504 288396 197510 288448
rect 322842 288396 322848 288448
rect 322900 288436 322906 288448
rect 327258 288436 327264 288448
rect 322900 288408 327264 288436
rect 322900 288396 322906 288408
rect 327258 288396 327264 288408
rect 327316 288396 327322 288448
rect 121454 288328 121460 288380
rect 121512 288368 121518 288380
rect 166350 288368 166356 288380
rect 121512 288340 166356 288368
rect 121512 288328 121518 288340
rect 166350 288328 166356 288340
rect 166408 288328 166414 288380
rect 121546 288260 121552 288312
rect 121604 288300 121610 288312
rect 151998 288300 152004 288312
rect 121604 288272 152004 288300
rect 121604 288260 121610 288272
rect 151998 288260 152004 288272
rect 152056 288300 152062 288312
rect 153102 288300 153108 288312
rect 152056 288272 153108 288300
rect 152056 288260 152062 288272
rect 153102 288260 153108 288272
rect 153160 288260 153166 288312
rect 153102 287648 153108 287700
rect 153160 287688 153166 287700
rect 165062 287688 165068 287700
rect 153160 287660 165068 287688
rect 153160 287648 153166 287660
rect 165062 287648 165068 287660
rect 165120 287648 165126 287700
rect 46750 287036 46756 287088
rect 46808 287076 46814 287088
rect 67634 287076 67640 287088
rect 46808 287048 67640 287076
rect 46808 287036 46814 287048
rect 67634 287036 67640 287048
rect 67692 287036 67698 287088
rect 362954 287036 362960 287088
rect 363012 287076 363018 287088
rect 364242 287076 364248 287088
rect 363012 287048 364248 287076
rect 363012 287036 363018 287048
rect 364242 287036 364248 287048
rect 364300 287076 364306 287088
rect 506474 287076 506480 287088
rect 364300 287048 506480 287076
rect 364300 287036 364306 287048
rect 506474 287036 506480 287048
rect 506532 287036 506538 287088
rect 55122 286968 55128 287020
rect 55180 287008 55186 287020
rect 67726 287008 67732 287020
rect 55180 286980 67732 287008
rect 55180 286968 55186 286980
rect 67726 286968 67732 286980
rect 67784 286968 67790 287020
rect 121546 286968 121552 287020
rect 121604 287008 121610 287020
rect 124214 287008 124220 287020
rect 121604 286980 124220 287008
rect 121604 286968 121610 286980
rect 124214 286968 124220 286980
rect 124272 286968 124278 287020
rect 60550 286900 60556 286952
rect 60608 286940 60614 286952
rect 67634 286940 67640 286952
rect 60608 286912 67640 286940
rect 60608 286900 60614 286912
rect 67634 286900 67640 286912
rect 67692 286900 67698 286952
rect 322198 286288 322204 286340
rect 322256 286328 322262 286340
rect 362954 286328 362960 286340
rect 322256 286300 362960 286328
rect 322256 286288 322262 286300
rect 362954 286288 362960 286300
rect 363012 286288 363018 286340
rect 182082 285744 182088 285796
rect 182140 285784 182146 285796
rect 197446 285784 197452 285796
rect 182140 285756 197452 285784
rect 182140 285744 182146 285756
rect 197446 285744 197452 285756
rect 197504 285744 197510 285796
rect 57514 285676 57520 285728
rect 57572 285716 57578 285728
rect 67818 285716 67824 285728
rect 57572 285688 67824 285716
rect 57572 285676 57578 285688
rect 67818 285676 67824 285688
rect 67876 285676 67882 285728
rect 120718 285676 120724 285728
rect 120776 285716 120782 285728
rect 196802 285716 196808 285728
rect 120776 285688 196808 285716
rect 120776 285676 120782 285688
rect 196802 285676 196808 285688
rect 196860 285676 196866 285728
rect 57790 285608 57796 285660
rect 57848 285648 57854 285660
rect 67634 285648 67640 285660
rect 57848 285620 67640 285648
rect 57848 285608 57854 285620
rect 67634 285608 67640 285620
rect 67692 285608 67698 285660
rect 121454 285608 121460 285660
rect 121512 285648 121518 285660
rect 193950 285648 193956 285660
rect 121512 285620 193956 285648
rect 121512 285608 121518 285620
rect 193950 285608 193956 285620
rect 194008 285608 194014 285660
rect 121546 285540 121552 285592
rect 121604 285580 121610 285592
rect 153194 285580 153200 285592
rect 121604 285552 153200 285580
rect 121604 285540 121610 285552
rect 153194 285540 153200 285552
rect 153252 285540 153258 285592
rect 43806 284316 43812 284368
rect 43864 284356 43870 284368
rect 67634 284356 67640 284368
rect 43864 284328 67640 284356
rect 43864 284316 43870 284328
rect 67634 284316 67640 284328
rect 67692 284316 67698 284368
rect 121454 284248 121460 284300
rect 121512 284288 121518 284300
rect 147122 284288 147128 284300
rect 121512 284260 147128 284288
rect 121512 284248 121518 284260
rect 147122 284248 147128 284260
rect 147180 284248 147186 284300
rect 127066 283568 127072 283620
rect 127124 283608 127130 283620
rect 179414 283608 179420 283620
rect 127124 283580 179420 283608
rect 127124 283568 127130 283580
rect 179414 283568 179420 283580
rect 179472 283568 179478 283620
rect 123570 282956 123576 283008
rect 123628 282996 123634 283008
rect 127066 282996 127072 283008
rect 123628 282968 127072 282996
rect 123628 282956 123634 282968
rect 127066 282956 127072 282968
rect 127124 282956 127130 283008
rect 121454 282888 121460 282940
rect 121512 282928 121518 282940
rect 127710 282928 127716 282940
rect 121512 282900 127716 282928
rect 121512 282888 121518 282900
rect 127710 282888 127716 282900
rect 127768 282888 127774 282940
rect 179414 282888 179420 282940
rect 179472 282928 179478 282940
rect 180702 282928 180708 282940
rect 179472 282900 180708 282928
rect 179472 282888 179478 282900
rect 180702 282888 180708 282900
rect 180760 282928 180766 282940
rect 197446 282928 197452 282940
rect 180760 282900 197452 282928
rect 180760 282888 180766 282900
rect 197446 282888 197452 282900
rect 197504 282888 197510 282940
rect 322474 282888 322480 282940
rect 322532 282928 322538 282940
rect 329926 282928 329932 282940
rect 322532 282900 329932 282928
rect 322532 282888 322538 282900
rect 329926 282888 329932 282900
rect 329984 282888 329990 282940
rect 43990 282820 43996 282872
rect 44048 282860 44054 282872
rect 67634 282860 67640 282872
rect 44048 282832 67640 282860
rect 44048 282820 44054 282832
rect 67634 282820 67640 282832
rect 67692 282820 67698 282872
rect 124950 282140 124956 282192
rect 125008 282180 125014 282192
rect 150618 282180 150624 282192
rect 125008 282152 150624 282180
rect 125008 282140 125014 282152
rect 150618 282140 150624 282152
rect 150676 282140 150682 282192
rect 184750 281596 184756 281648
rect 184808 281636 184814 281648
rect 190454 281636 190460 281648
rect 184808 281608 190460 281636
rect 184808 281596 184814 281608
rect 190454 281596 190460 281608
rect 190512 281636 190518 281648
rect 191742 281636 191748 281648
rect 190512 281608 191748 281636
rect 190512 281596 190518 281608
rect 191742 281596 191748 281608
rect 191800 281596 191806 281648
rect 121454 281528 121460 281580
rect 121512 281568 121518 281580
rect 170398 281568 170404 281580
rect 121512 281540 170404 281568
rect 121512 281528 121518 281540
rect 170398 281528 170404 281540
rect 170456 281528 170462 281580
rect 173342 281528 173348 281580
rect 173400 281568 173406 281580
rect 197446 281568 197452 281580
rect 173400 281540 197452 281568
rect 173400 281528 173406 281540
rect 197446 281528 197452 281540
rect 197504 281528 197510 281580
rect 121546 281460 121552 281512
rect 121604 281500 121610 281512
rect 192478 281500 192484 281512
rect 121604 281472 192484 281500
rect 121604 281460 121610 281472
rect 192478 281460 192484 281472
rect 192536 281460 192542 281512
rect 191742 281392 191748 281444
rect 191800 281432 191806 281444
rect 197446 281432 197452 281444
rect 191800 281404 197452 281432
rect 191800 281392 191806 281404
rect 197446 281392 197452 281404
rect 197504 281392 197510 281444
rect 45462 280168 45468 280220
rect 45520 280208 45526 280220
rect 67634 280208 67640 280220
rect 45520 280180 67640 280208
rect 45520 280168 45526 280180
rect 67634 280168 67640 280180
rect 67692 280168 67698 280220
rect 121454 280168 121460 280220
rect 121512 280208 121518 280220
rect 148410 280208 148416 280220
rect 121512 280180 148416 280208
rect 121512 280168 121518 280180
rect 148410 280168 148416 280180
rect 148468 280168 148474 280220
rect 322474 280168 322480 280220
rect 322532 280208 322538 280220
rect 335998 280208 336004 280220
rect 322532 280180 336004 280208
rect 322532 280168 322538 280180
rect 335998 280168 336004 280180
rect 336056 280168 336062 280220
rect 40862 280100 40868 280152
rect 40920 280140 40926 280152
rect 41138 280140 41144 280152
rect 40920 280112 41144 280140
rect 40920 280100 40926 280112
rect 41138 280100 41144 280112
rect 41196 280140 41202 280152
rect 67726 280140 67732 280152
rect 41196 280112 67732 280140
rect 41196 280100 41202 280112
rect 67726 280100 67732 280112
rect 67784 280100 67790 280152
rect 121546 280100 121552 280152
rect 121604 280140 121610 280152
rect 130378 280140 130384 280152
rect 121604 280112 130384 280140
rect 121604 280100 121610 280112
rect 130378 280100 130384 280112
rect 130436 280100 130442 280152
rect 29638 279420 29644 279472
rect 29696 279460 29702 279472
rect 40862 279460 40868 279472
rect 29696 279432 40868 279460
rect 29696 279420 29702 279432
rect 40862 279420 40868 279432
rect 40920 279420 40926 279472
rect 52270 279420 52276 279472
rect 52328 279460 52334 279472
rect 57790 279460 57796 279472
rect 52328 279432 57796 279460
rect 52328 279420 52334 279432
rect 57790 279420 57796 279432
rect 57848 279460 57854 279472
rect 67634 279460 67640 279472
rect 57848 279432 67640 279460
rect 57848 279420 57854 279432
rect 67634 279420 67640 279432
rect 67692 279420 67698 279472
rect 123754 279420 123760 279472
rect 123812 279460 123818 279472
rect 163682 279460 163688 279472
rect 123812 279432 163688 279460
rect 123812 279420 123818 279432
rect 163682 279420 163688 279432
rect 163740 279420 163746 279472
rect 121454 278740 121460 278792
rect 121512 278780 121518 278792
rect 192478 278780 192484 278792
rect 121512 278752 192484 278780
rect 121512 278740 121518 278752
rect 192478 278740 192484 278752
rect 192536 278740 192542 278792
rect 121546 278672 121552 278724
rect 121604 278712 121610 278724
rect 184842 278712 184848 278724
rect 121604 278684 184848 278712
rect 121604 278672 121610 278684
rect 184842 278672 184848 278684
rect 184900 278672 184906 278724
rect 184842 278196 184848 278248
rect 184900 278236 184906 278248
rect 187050 278236 187056 278248
rect 184900 278208 187056 278236
rect 184900 278196 184906 278208
rect 187050 278196 187056 278208
rect 187108 278196 187114 278248
rect 195790 277448 195796 277500
rect 195848 277488 195854 277500
rect 197446 277488 197452 277500
rect 195848 277460 197452 277488
rect 195848 277448 195854 277460
rect 197446 277448 197452 277460
rect 197504 277448 197510 277500
rect 47946 277380 47952 277432
rect 48004 277420 48010 277432
rect 67634 277420 67640 277432
rect 48004 277392 67640 277420
rect 48004 277380 48010 277392
rect 67634 277380 67640 277392
rect 67692 277380 67698 277432
rect 121454 277312 121460 277364
rect 121512 277352 121518 277364
rect 131114 277352 131120 277364
rect 121512 277324 131120 277352
rect 121512 277312 121518 277324
rect 131114 277312 131120 277324
rect 131172 277312 131178 277364
rect 61838 276632 61844 276684
rect 61896 276672 61902 276684
rect 67634 276672 67640 276684
rect 61896 276644 67640 276672
rect 61896 276632 61902 276644
rect 67634 276632 67640 276644
rect 67692 276632 67698 276684
rect 322198 276088 322204 276140
rect 322256 276128 322262 276140
rect 322256 276100 325694 276128
rect 322256 276088 322262 276100
rect 121454 276020 121460 276072
rect 121512 276060 121518 276072
rect 130562 276060 130568 276072
rect 121512 276032 130568 276060
rect 121512 276020 121518 276032
rect 130562 276020 130568 276032
rect 130620 276020 130626 276072
rect 322842 276020 322848 276072
rect 322900 276060 322906 276072
rect 325050 276060 325056 276072
rect 322900 276032 325056 276060
rect 322900 276020 322906 276032
rect 325050 276020 325056 276032
rect 325108 276020 325114 276072
rect 325666 276060 325694 276100
rect 521654 276060 521660 276072
rect 325666 276032 521660 276060
rect 521654 276020 521660 276032
rect 521712 276020 521718 276072
rect 191742 275408 191748 275460
rect 191800 275448 191806 275460
rect 197354 275448 197360 275460
rect 191800 275420 197360 275448
rect 191800 275408 191806 275420
rect 197354 275408 197360 275420
rect 197412 275408 197418 275460
rect 121546 274796 121552 274848
rect 121604 274836 121610 274848
rect 128262 274836 128268 274848
rect 121604 274808 128268 274836
rect 121604 274796 121610 274808
rect 128262 274796 128268 274808
rect 128320 274836 128326 274848
rect 129918 274836 129924 274848
rect 128320 274808 129924 274836
rect 128320 274796 128326 274808
rect 129918 274796 129924 274808
rect 129976 274796 129982 274848
rect 121454 274728 121460 274780
rect 121512 274768 121518 274780
rect 131850 274768 131856 274780
rect 121512 274740 131856 274768
rect 121512 274728 121518 274740
rect 131850 274728 131856 274740
rect 131908 274728 131914 274780
rect 53650 274660 53656 274712
rect 53708 274700 53714 274712
rect 67634 274700 67640 274712
rect 53708 274672 67640 274700
rect 53708 274660 53714 274672
rect 67634 274660 67640 274672
rect 67692 274660 67698 274712
rect 121546 274660 121552 274712
rect 121604 274700 121610 274712
rect 122098 274700 122104 274712
rect 121604 274672 122104 274700
rect 121604 274660 121610 274672
rect 122098 274660 122104 274672
rect 122156 274700 122162 274712
rect 162394 274700 162400 274712
rect 122156 274672 162400 274700
rect 122156 274660 122162 274672
rect 162394 274660 162400 274672
rect 162452 274660 162458 274712
rect 187142 274660 187148 274712
rect 187200 274700 187206 274712
rect 197354 274700 197360 274712
rect 187200 274672 197360 274700
rect 187200 274660 187206 274672
rect 197354 274660 197360 274672
rect 197412 274660 197418 274712
rect 52086 274592 52092 274644
rect 52144 274632 52150 274644
rect 67726 274632 67732 274644
rect 52144 274604 67732 274632
rect 52144 274592 52150 274604
rect 67726 274592 67732 274604
rect 67784 274592 67790 274644
rect 322382 274592 322388 274644
rect 322440 274632 322446 274644
rect 339586 274632 339592 274644
rect 322440 274604 339592 274632
rect 322440 274592 322446 274604
rect 339586 274592 339592 274604
rect 339644 274592 339650 274644
rect 339586 273912 339592 273964
rect 339644 273952 339650 273964
rect 382918 273952 382924 273964
rect 339644 273924 382924 273952
rect 339644 273912 339650 273924
rect 382918 273912 382924 273924
rect 382976 273912 382982 273964
rect 121454 273300 121460 273352
rect 121512 273340 121518 273352
rect 171870 273340 171876 273352
rect 121512 273312 171876 273340
rect 121512 273300 121518 273312
rect 171870 273300 171876 273312
rect 171928 273300 171934 273352
rect 52270 273232 52276 273284
rect 52328 273272 52334 273284
rect 67634 273272 67640 273284
rect 52328 273244 67640 273272
rect 52328 273232 52334 273244
rect 67634 273232 67640 273244
rect 67692 273232 67698 273284
rect 123478 273232 123484 273284
rect 123536 273272 123542 273284
rect 194502 273272 194508 273284
rect 123536 273244 194508 273272
rect 123536 273232 123542 273244
rect 194502 273232 194508 273244
rect 194560 273272 194566 273284
rect 197354 273272 197360 273284
rect 194560 273244 197360 273272
rect 194560 273232 194566 273244
rect 197354 273232 197360 273244
rect 197412 273232 197418 273284
rect 121454 273164 121460 273216
rect 121512 273204 121518 273216
rect 133874 273204 133880 273216
rect 121512 273176 133880 273204
rect 121512 273164 121518 273176
rect 133874 273164 133880 273176
rect 133932 273164 133938 273216
rect 125134 271872 125140 271924
rect 125192 271912 125198 271924
rect 187142 271912 187148 271924
rect 125192 271884 187148 271912
rect 125192 271872 125198 271884
rect 187142 271872 187148 271884
rect 187200 271872 187206 271924
rect 335998 271872 336004 271924
rect 336056 271912 336062 271924
rect 400858 271912 400864 271924
rect 336056 271884 400864 271912
rect 336056 271872 336062 271884
rect 400858 271872 400864 271884
rect 400916 271872 400922 271924
rect 417418 271872 417424 271924
rect 417476 271912 417482 271924
rect 419534 271912 419540 271924
rect 417476 271884 419540 271912
rect 417476 271872 417482 271884
rect 419534 271872 419540 271884
rect 419592 271912 419598 271924
rect 580166 271912 580172 271924
rect 419592 271884 580172 271912
rect 419592 271872 419598 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 57698 271804 57704 271856
rect 57756 271844 57762 271856
rect 67726 271844 67732 271856
rect 57756 271816 67732 271844
rect 57756 271804 57762 271816
rect 67726 271804 67732 271816
rect 67784 271804 67790 271856
rect 127710 271124 127716 271176
rect 127768 271164 127774 271176
rect 197354 271164 197360 271176
rect 127768 271136 197360 271164
rect 127768 271124 127774 271136
rect 197354 271124 197360 271136
rect 197412 271124 197418 271176
rect 63218 270512 63224 270564
rect 63276 270552 63282 270564
rect 67634 270552 67640 270564
rect 63276 270524 67640 270552
rect 63276 270512 63282 270524
rect 67634 270512 67640 270524
rect 67692 270512 67698 270564
rect 121454 270512 121460 270564
rect 121512 270552 121518 270564
rect 173250 270552 173256 270564
rect 121512 270524 173256 270552
rect 121512 270512 121518 270524
rect 173250 270512 173256 270524
rect 173308 270512 173314 270564
rect 322842 270512 322848 270564
rect 322900 270552 322906 270564
rect 331306 270552 331312 270564
rect 322900 270524 331312 270552
rect 322900 270512 322906 270524
rect 331306 270512 331312 270524
rect 331364 270512 331370 270564
rect 56318 270444 56324 270496
rect 56376 270484 56382 270496
rect 67726 270484 67732 270496
rect 56376 270456 67732 270484
rect 56376 270444 56382 270456
rect 67726 270444 67732 270456
rect 67784 270444 67790 270496
rect 57698 269764 57704 269816
rect 57756 269804 57762 269816
rect 67818 269804 67824 269816
rect 57756 269776 67824 269804
rect 57756 269764 57762 269776
rect 67818 269764 67824 269776
rect 67876 269764 67882 269816
rect 66070 269084 66076 269136
rect 66128 269124 66134 269136
rect 68186 269124 68192 269136
rect 66128 269096 68192 269124
rect 66128 269084 66134 269096
rect 68186 269084 68192 269096
rect 68244 269084 68250 269136
rect 121546 269084 121552 269136
rect 121604 269124 121610 269136
rect 130378 269124 130384 269136
rect 121604 269096 130384 269124
rect 121604 269084 121610 269096
rect 130378 269084 130384 269096
rect 130436 269084 130442 269136
rect 322842 269084 322848 269136
rect 322900 269124 322906 269136
rect 326338 269124 326344 269136
rect 322900 269096 326344 269124
rect 322900 269084 322906 269096
rect 326338 269084 326344 269096
rect 326396 269084 326402 269136
rect 52454 269016 52460 269068
rect 52512 269056 52518 269068
rect 53558 269056 53564 269068
rect 52512 269028 53564 269056
rect 52512 269016 52518 269028
rect 53558 269016 53564 269028
rect 53616 269056 53622 269068
rect 67634 269056 67640 269068
rect 53616 269028 67640 269056
rect 53616 269016 53622 269028
rect 67634 269016 67640 269028
rect 67692 269016 67698 269068
rect 121454 269016 121460 269068
rect 121512 269056 121518 269068
rect 149146 269056 149152 269068
rect 121512 269028 149152 269056
rect 121512 269016 121518 269028
rect 149146 269016 149152 269028
rect 149204 269056 149210 269068
rect 149330 269056 149336 269068
rect 149204 269028 149336 269056
rect 149204 269016 149210 269028
rect 149330 269016 149336 269028
rect 149388 269016 149394 269068
rect 45278 268404 45284 268456
rect 45336 268444 45342 268456
rect 52086 268444 52092 268456
rect 45336 268416 52092 268444
rect 45336 268404 45342 268416
rect 52086 268404 52092 268416
rect 52144 268404 52150 268456
rect 149330 268404 149336 268456
rect 149388 268444 149394 268456
rect 181622 268444 181628 268456
rect 149388 268416 181628 268444
rect 149388 268404 149394 268416
rect 181622 268404 181628 268416
rect 181680 268404 181686 268456
rect 21358 268336 21364 268388
rect 21416 268376 21422 268388
rect 52454 268376 52460 268388
rect 21416 268348 52460 268376
rect 21416 268336 21422 268348
rect 52454 268336 52460 268348
rect 52512 268336 52518 268388
rect 125042 268336 125048 268388
rect 125100 268376 125106 268388
rect 183370 268376 183376 268388
rect 125100 268348 183376 268376
rect 125100 268336 125106 268348
rect 183370 268336 183376 268348
rect 183428 268336 183434 268388
rect 183370 267792 183376 267844
rect 183428 267832 183434 267844
rect 197354 267832 197360 267844
rect 183428 267804 197360 267832
rect 183428 267792 183434 267804
rect 197354 267792 197360 267804
rect 197412 267792 197418 267844
rect 121454 267724 121460 267776
rect 121512 267764 121518 267776
rect 191190 267764 191196 267776
rect 121512 267736 191196 267764
rect 121512 267724 121518 267736
rect 191190 267724 191196 267736
rect 191248 267724 191254 267776
rect 48130 267656 48136 267708
rect 48188 267696 48194 267708
rect 67726 267696 67732 267708
rect 48188 267668 67732 267696
rect 48188 267656 48194 267668
rect 67726 267656 67732 267668
rect 67784 267656 67790 267708
rect 322474 267656 322480 267708
rect 322532 267696 322538 267708
rect 342254 267696 342260 267708
rect 322532 267668 342260 267696
rect 322532 267656 322538 267668
rect 342254 267656 342260 267668
rect 342312 267656 342318 267708
rect 52086 266976 52092 267028
rect 52144 267016 52150 267028
rect 67634 267016 67640 267028
rect 52144 266988 67640 267016
rect 52144 266976 52150 266988
rect 67634 266976 67640 266988
rect 67692 266976 67698 267028
rect 160830 266976 160836 267028
rect 160888 267016 160894 267028
rect 176654 267016 176660 267028
rect 160888 266988 176660 267016
rect 160888 266976 160894 266988
rect 176654 266976 176660 266988
rect 176712 266976 176718 267028
rect 342254 266976 342260 267028
rect 342312 267016 342318 267028
rect 499850 267016 499856 267028
rect 342312 266988 499856 267016
rect 342312 266976 342318 266988
rect 499850 266976 499856 266988
rect 499908 266976 499914 267028
rect 121454 266432 121460 266484
rect 121512 266472 121518 266484
rect 147214 266472 147220 266484
rect 121512 266444 147220 266472
rect 121512 266432 121518 266444
rect 147214 266432 147220 266444
rect 147272 266432 147278 266484
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 54478 266404 54484 266416
rect 3108 266376 54484 266404
rect 3108 266364 3114 266376
rect 54478 266364 54484 266376
rect 54536 266364 54542 266416
rect 121546 266364 121552 266416
rect 121604 266404 121610 266416
rect 149790 266404 149796 266416
rect 121604 266376 149796 266404
rect 121604 266364 121610 266376
rect 149790 266364 149796 266376
rect 149848 266364 149854 266416
rect 176654 266364 176660 266416
rect 176712 266404 176718 266416
rect 177850 266404 177856 266416
rect 176712 266376 177856 266404
rect 176712 266364 176718 266376
rect 177850 266364 177856 266376
rect 177908 266404 177914 266416
rect 197354 266404 197360 266416
rect 177908 266376 197360 266404
rect 177908 266364 177914 266376
rect 197354 266364 197360 266376
rect 197412 266364 197418 266416
rect 54846 266296 54852 266348
rect 54904 266336 54910 266348
rect 67726 266336 67732 266348
rect 54904 266308 67732 266336
rect 54904 266296 54910 266308
rect 67726 266296 67732 266308
rect 67784 266296 67790 266348
rect 121454 265004 121460 265056
rect 121512 265044 121518 265056
rect 152642 265044 152648 265056
rect 121512 265016 152648 265044
rect 121512 265004 121518 265016
rect 152642 265004 152648 265016
rect 152700 265004 152706 265056
rect 54938 264936 54944 264988
rect 54996 264976 55002 264988
rect 67634 264976 67640 264988
rect 54996 264948 67640 264976
rect 54996 264936 55002 264948
rect 67634 264936 67640 264948
rect 67692 264936 67698 264988
rect 68554 264936 68560 264988
rect 68612 264976 68618 264988
rect 68830 264976 68836 264988
rect 68612 264948 68836 264976
rect 68612 264936 68618 264948
rect 68830 264936 68836 264948
rect 68888 264936 68894 264988
rect 121546 264936 121552 264988
rect 121604 264976 121610 264988
rect 158162 264976 158168 264988
rect 121604 264948 158168 264976
rect 121604 264936 121610 264948
rect 158162 264936 158168 264948
rect 158220 264936 158226 264988
rect 322474 264936 322480 264988
rect 322532 264976 322538 264988
rect 330018 264976 330024 264988
rect 322532 264948 330024 264976
rect 322532 264936 322538 264948
rect 330018 264936 330024 264948
rect 330076 264936 330082 264988
rect 14458 264188 14464 264240
rect 14516 264228 14522 264240
rect 43898 264228 43904 264240
rect 14516 264200 43904 264228
rect 14516 264188 14522 264200
rect 43898 264188 43904 264200
rect 43956 264228 43962 264240
rect 55858 264228 55864 264240
rect 43956 264200 55864 264228
rect 43956 264188 43962 264200
rect 55858 264188 55864 264200
rect 55916 264188 55922 264240
rect 124122 264188 124128 264240
rect 124180 264228 124186 264240
rect 195698 264228 195704 264240
rect 124180 264200 195704 264228
rect 124180 264188 124186 264200
rect 195698 264188 195704 264200
rect 195756 264228 195762 264240
rect 197354 264228 197360 264240
rect 195756 264200 197360 264228
rect 195756 264188 195762 264200
rect 197354 264188 197360 264200
rect 197412 264188 197418 264240
rect 56226 263644 56232 263696
rect 56284 263684 56290 263696
rect 67634 263684 67640 263696
rect 56284 263656 67640 263684
rect 56284 263644 56290 263656
rect 67634 263644 67640 263656
rect 67692 263644 67698 263696
rect 55858 263576 55864 263628
rect 55916 263616 55922 263628
rect 56318 263616 56324 263628
rect 55916 263588 56324 263616
rect 55916 263576 55922 263588
rect 56318 263576 56324 263588
rect 56376 263616 56382 263628
rect 67726 263616 67732 263628
rect 56376 263588 67732 263616
rect 56376 263576 56382 263588
rect 67726 263576 67732 263588
rect 67784 263576 67790 263628
rect 121546 263576 121552 263628
rect 121604 263616 121610 263628
rect 134702 263616 134708 263628
rect 121604 263588 134708 263616
rect 121604 263576 121610 263588
rect 134702 263576 134708 263588
rect 134760 263576 134766 263628
rect 335262 263576 335268 263628
rect 335320 263616 335326 263628
rect 490558 263616 490564 263628
rect 335320 263588 490564 263616
rect 335320 263576 335326 263588
rect 490558 263576 490564 263588
rect 490616 263576 490622 263628
rect 56502 263508 56508 263560
rect 56560 263548 56566 263560
rect 67634 263548 67640 263560
rect 56560 263520 67640 263548
rect 56560 263508 56566 263520
rect 67634 263508 67640 263520
rect 67692 263508 67698 263560
rect 121454 263508 121460 263560
rect 121512 263548 121518 263560
rect 136726 263548 136732 263560
rect 121512 263520 136732 263548
rect 121512 263508 121518 263520
rect 136726 263508 136732 263520
rect 136784 263548 136790 263560
rect 137094 263548 137100 263560
rect 136784 263520 137100 263548
rect 136784 263508 136790 263520
rect 137094 263508 137100 263520
rect 137152 263508 137158 263560
rect 332594 263508 332600 263560
rect 332652 263548 332658 263560
rect 335280 263548 335308 263576
rect 332652 263520 335308 263548
rect 332652 263508 332658 263520
rect 68554 262896 68560 262948
rect 68612 262936 68618 262948
rect 68922 262936 68928 262948
rect 68612 262908 68928 262936
rect 68612 262896 68618 262908
rect 68922 262896 68928 262908
rect 68980 262896 68986 262948
rect 137094 262828 137100 262880
rect 137152 262868 137158 262880
rect 178770 262868 178776 262880
rect 137152 262840 178776 262868
rect 137152 262828 137158 262840
rect 178770 262828 178776 262840
rect 178828 262828 178834 262880
rect 121454 262760 121460 262812
rect 121512 262800 121518 262812
rect 125134 262800 125140 262812
rect 121512 262772 125140 262800
rect 121512 262760 121518 262772
rect 125134 262760 125140 262772
rect 125192 262760 125198 262812
rect 56502 262216 56508 262268
rect 56560 262256 56566 262268
rect 67634 262256 67640 262268
rect 56560 262228 67640 262256
rect 56560 262216 56566 262228
rect 67634 262216 67640 262228
rect 67692 262216 67698 262268
rect 322474 262216 322480 262268
rect 322532 262256 322538 262268
rect 332594 262256 332600 262268
rect 322532 262228 332600 262256
rect 322532 262216 322538 262228
rect 332594 262216 332600 262228
rect 332652 262216 332658 262268
rect 65978 262148 65984 262200
rect 66036 262188 66042 262200
rect 67726 262188 67732 262200
rect 66036 262160 67732 262188
rect 66036 262148 66042 262160
rect 67726 262148 67732 262160
rect 67784 262148 67790 262200
rect 121546 262148 121552 262200
rect 121604 262188 121610 262200
rect 126882 262188 126888 262200
rect 121604 262160 126888 262188
rect 121604 262148 121610 262160
rect 126882 262148 126888 262160
rect 126940 262148 126946 262200
rect 121454 261876 121460 261928
rect 121512 261916 121518 261928
rect 123478 261916 123484 261928
rect 121512 261888 123484 261916
rect 121512 261876 121518 261888
rect 123478 261876 123484 261888
rect 123536 261876 123542 261928
rect 126882 261468 126888 261520
rect 126940 261508 126946 261520
rect 160922 261508 160928 261520
rect 126940 261480 160928 261508
rect 126940 261468 126946 261480
rect 160922 261468 160928 261480
rect 160980 261468 160986 261520
rect 140038 260856 140044 260908
rect 140096 260896 140102 260908
rect 190270 260896 190276 260908
rect 140096 260868 190276 260896
rect 140096 260856 140102 260868
rect 190270 260856 190276 260868
rect 190328 260896 190334 260908
rect 197354 260896 197360 260908
rect 190328 260868 197360 260896
rect 190328 260856 190334 260868
rect 197354 260856 197360 260868
rect 197412 260856 197418 260908
rect 56410 260788 56416 260840
rect 56468 260828 56474 260840
rect 67634 260828 67640 260840
rect 56468 260800 67640 260828
rect 56468 260788 56474 260800
rect 67634 260788 67640 260800
rect 67692 260788 67698 260840
rect 121454 260788 121460 260840
rect 121512 260828 121518 260840
rect 139578 260828 139584 260840
rect 121512 260800 139584 260828
rect 121512 260788 121518 260800
rect 139578 260788 139584 260800
rect 139636 260828 139642 260840
rect 140682 260828 140688 260840
rect 139636 260800 140688 260828
rect 139636 260788 139642 260800
rect 140682 260788 140688 260800
rect 140740 260788 140746 260840
rect 370498 260108 370504 260160
rect 370556 260148 370562 260160
rect 548518 260148 548524 260160
rect 370556 260120 548524 260148
rect 370556 260108 370562 260120
rect 548518 260108 548524 260120
rect 548576 260108 548582 260160
rect 139578 259496 139584 259548
rect 139636 259536 139642 259548
rect 144178 259536 144184 259548
rect 139636 259508 144184 259536
rect 139636 259496 139642 259508
rect 144178 259496 144184 259508
rect 144236 259496 144242 259548
rect 121454 259428 121460 259480
rect 121512 259468 121518 259480
rect 170674 259468 170680 259480
rect 121512 259440 170680 259468
rect 121512 259428 121518 259440
rect 170674 259428 170680 259440
rect 170732 259428 170738 259480
rect 179874 259428 179880 259480
rect 179932 259468 179938 259480
rect 197354 259468 197360 259480
rect 179932 259440 197360 259468
rect 179932 259428 179938 259440
rect 197354 259428 197360 259440
rect 197412 259428 197418 259480
rect 322566 259428 322572 259480
rect 322624 259468 322630 259480
rect 327350 259468 327356 259480
rect 322624 259440 327356 259468
rect 322624 259428 322630 259440
rect 327350 259428 327356 259440
rect 327408 259428 327414 259480
rect 121546 259360 121552 259412
rect 121604 259400 121610 259412
rect 143626 259400 143632 259412
rect 121604 259372 143632 259400
rect 121604 259360 121610 259372
rect 143626 259360 143632 259372
rect 143684 259400 143690 259412
rect 144822 259400 144828 259412
rect 143684 259372 144828 259400
rect 143684 259360 143690 259372
rect 144822 259360 144828 259372
rect 144880 259360 144886 259412
rect 144822 258680 144828 258732
rect 144880 258720 144886 258732
rect 166534 258720 166540 258732
rect 144880 258692 166540 258720
rect 144880 258680 144886 258692
rect 166534 258680 166540 258692
rect 166592 258680 166598 258732
rect 548518 258680 548524 258732
rect 548576 258720 548582 258732
rect 579982 258720 579988 258732
rect 548576 258692 579988 258720
rect 548576 258680 548582 258692
rect 579982 258680 579988 258692
rect 580040 258680 580046 258732
rect 61838 258068 61844 258120
rect 61896 258108 61902 258120
rect 67726 258108 67732 258120
rect 61896 258080 67732 258108
rect 61896 258068 61902 258080
rect 67726 258068 67732 258080
rect 67784 258068 67790 258120
rect 121638 258068 121644 258120
rect 121696 258108 121702 258120
rect 154114 258108 154120 258120
rect 121696 258080 154120 258108
rect 121696 258068 121702 258080
rect 154114 258068 154120 258080
rect 154172 258068 154178 258120
rect 324406 258068 324412 258120
rect 324464 258108 324470 258120
rect 425054 258108 425060 258120
rect 324464 258080 425060 258108
rect 324464 258068 324470 258080
rect 425054 258068 425060 258080
rect 425112 258068 425118 258120
rect 34422 258000 34428 258052
rect 34480 258040 34486 258052
rect 67634 258040 67640 258052
rect 34480 258012 67640 258040
rect 34480 258000 34486 258012
rect 67634 258000 67640 258012
rect 67692 258000 67698 258052
rect 121454 258000 121460 258052
rect 121512 258040 121518 258052
rect 154574 258040 154580 258052
rect 121512 258012 154580 258040
rect 121512 258000 121518 258012
rect 154574 258000 154580 258012
rect 154632 258000 154638 258052
rect 15838 257320 15844 257372
rect 15896 257360 15902 257372
rect 34422 257360 34428 257372
rect 15896 257332 34428 257360
rect 15896 257320 15902 257332
rect 34422 257320 34428 257332
rect 34480 257320 34486 257372
rect 131758 257320 131764 257372
rect 131816 257360 131822 257372
rect 197354 257360 197360 257372
rect 131816 257332 197360 257360
rect 131816 257320 131822 257332
rect 197354 257320 197360 257332
rect 197412 257320 197418 257372
rect 65978 256708 65984 256760
rect 66036 256748 66042 256760
rect 68002 256748 68008 256760
rect 66036 256720 68008 256748
rect 66036 256708 66042 256720
rect 68002 256708 68008 256720
rect 68060 256708 68066 256760
rect 121546 256708 121552 256760
rect 121604 256748 121610 256760
rect 134518 256748 134524 256760
rect 121604 256720 134524 256748
rect 121604 256708 121610 256720
rect 134518 256708 134524 256720
rect 134576 256708 134582 256760
rect 121454 256640 121460 256692
rect 121512 256680 121518 256692
rect 148594 256680 148600 256692
rect 121512 256652 148600 256680
rect 121512 256640 121518 256652
rect 148594 256640 148600 256652
rect 148652 256640 148658 256692
rect 121546 256572 121552 256624
rect 121604 256612 121610 256624
rect 133874 256612 133880 256624
rect 121604 256584 133880 256612
rect 121604 256572 121610 256584
rect 133874 256572 133880 256584
rect 133932 256612 133938 256624
rect 135162 256612 135168 256624
rect 133932 256584 135168 256612
rect 133932 256572 133938 256584
rect 135162 256572 135168 256584
rect 135220 256572 135226 256624
rect 135162 255960 135168 256012
rect 135220 256000 135226 256012
rect 166350 256000 166356 256012
rect 135220 255972 166356 256000
rect 135220 255960 135226 255972
rect 166350 255960 166356 255972
rect 166408 255960 166414 256012
rect 178770 255348 178776 255400
rect 178828 255388 178834 255400
rect 180610 255388 180616 255400
rect 178828 255360 180616 255388
rect 178828 255348 178834 255360
rect 180610 255348 180616 255360
rect 180668 255388 180674 255400
rect 180668 255360 180794 255388
rect 180668 255348 180674 255360
rect 53558 255280 53564 255332
rect 53616 255320 53622 255332
rect 67634 255320 67640 255332
rect 53616 255292 67640 255320
rect 53616 255280 53622 255292
rect 67634 255280 67640 255292
rect 67692 255280 67698 255332
rect 176102 255280 176108 255332
rect 176160 255320 176166 255332
rect 179874 255320 179880 255332
rect 176160 255292 179880 255320
rect 176160 255280 176166 255292
rect 179874 255280 179880 255292
rect 179932 255280 179938 255332
rect 180766 255320 180794 255360
rect 197354 255320 197360 255332
rect 180766 255292 197360 255320
rect 197354 255280 197360 255292
rect 197412 255280 197418 255332
rect 50982 255212 50988 255264
rect 51040 255252 51046 255264
rect 67726 255252 67732 255264
rect 51040 255224 67732 255252
rect 51040 255212 51046 255224
rect 67726 255212 67732 255224
rect 67784 255212 67790 255264
rect 143442 255212 143448 255264
rect 143500 255252 143506 255264
rect 194042 255252 194048 255264
rect 143500 255224 194048 255252
rect 143500 255212 143506 255224
rect 194042 255212 194048 255224
rect 194100 255212 194106 255264
rect 52178 255144 52184 255196
rect 52236 255184 52242 255196
rect 67634 255184 67640 255196
rect 52236 255156 67640 255184
rect 52236 255144 52242 255156
rect 67634 255144 67640 255156
rect 67692 255144 67698 255196
rect 142982 254804 142988 254856
rect 143040 254844 143046 254856
rect 143442 254844 143448 254856
rect 143040 254816 143448 254844
rect 143040 254804 143046 254816
rect 143442 254804 143448 254816
rect 143500 254804 143506 254856
rect 121454 253920 121460 253972
rect 121512 253960 121518 253972
rect 161014 253960 161020 253972
rect 121512 253932 161020 253960
rect 121512 253920 121518 253932
rect 161014 253920 161020 253932
rect 161072 253920 161078 253972
rect 48314 253852 48320 253904
rect 48372 253892 48378 253904
rect 48958 253892 48964 253904
rect 48372 253864 48964 253892
rect 48372 253852 48378 253864
rect 48958 253852 48964 253864
rect 49016 253892 49022 253904
rect 67634 253892 67640 253904
rect 49016 253864 67640 253892
rect 49016 253852 49022 253864
rect 67634 253852 67640 253864
rect 67692 253852 67698 253904
rect 32398 253172 32404 253224
rect 32456 253212 32462 253224
rect 48958 253212 48964 253224
rect 32456 253184 48964 253212
rect 32456 253172 32462 253184
rect 48958 253172 48964 253184
rect 49016 253172 49022 253224
rect 121454 252628 121460 252680
rect 121512 252668 121518 252680
rect 126330 252668 126336 252680
rect 121512 252640 126336 252668
rect 121512 252628 121518 252640
rect 126330 252628 126336 252640
rect 126388 252628 126394 252680
rect 121546 252560 121552 252612
rect 121604 252600 121610 252612
rect 155494 252600 155500 252612
rect 121604 252572 155500 252600
rect 121604 252560 121610 252572
rect 155494 252560 155500 252572
rect 155552 252560 155558 252612
rect 191282 252560 191288 252612
rect 191340 252600 191346 252612
rect 197354 252600 197360 252612
rect 191340 252572 197360 252600
rect 191340 252560 191346 252572
rect 197354 252560 197360 252572
rect 197412 252560 197418 252612
rect 121454 252492 121460 252544
rect 121512 252532 121518 252544
rect 155954 252532 155960 252544
rect 121512 252504 155960 252532
rect 121512 252492 121518 252504
rect 155954 252492 155960 252504
rect 156012 252492 156018 252544
rect 322474 251268 322480 251320
rect 322532 251308 322538 251320
rect 325786 251308 325792 251320
rect 322532 251280 325792 251308
rect 322532 251268 322538 251280
rect 325786 251268 325792 251280
rect 325844 251268 325850 251320
rect 61746 251200 61752 251252
rect 61804 251240 61810 251252
rect 67634 251240 67640 251252
rect 61804 251212 67640 251240
rect 61804 251200 61810 251212
rect 67634 251200 67640 251212
rect 67692 251200 67698 251252
rect 121454 251200 121460 251252
rect 121512 251240 121518 251252
rect 188614 251240 188620 251252
rect 121512 251212 188620 251240
rect 121512 251200 121518 251212
rect 188614 251200 188620 251212
rect 188672 251200 188678 251252
rect 66162 251132 66168 251184
rect 66220 251172 66226 251184
rect 67726 251172 67732 251184
rect 66220 251144 67732 251172
rect 66220 251132 66226 251144
rect 67726 251132 67732 251144
rect 67784 251132 67790 251184
rect 120626 251132 120632 251184
rect 120684 251172 120690 251184
rect 140958 251172 140964 251184
rect 120684 251144 140964 251172
rect 120684 251132 120690 251144
rect 140958 251132 140964 251144
rect 141016 251132 141022 251184
rect 121454 249772 121460 249824
rect 121512 249812 121518 249824
rect 137462 249812 137468 249824
rect 121512 249784 137468 249812
rect 121512 249772 121518 249784
rect 137462 249772 137468 249784
rect 137520 249772 137526 249824
rect 121546 249704 121552 249756
rect 121604 249744 121610 249756
rect 129182 249744 129188 249756
rect 121604 249716 129188 249744
rect 121604 249704 121610 249716
rect 129182 249704 129188 249716
rect 129240 249704 129246 249756
rect 39850 249024 39856 249076
rect 39908 249064 39914 249076
rect 57606 249064 57612 249076
rect 39908 249036 57612 249064
rect 39908 249024 39914 249036
rect 57606 249024 57612 249036
rect 57664 249024 57670 249076
rect 189810 249024 189816 249076
rect 189868 249064 189874 249076
rect 194410 249064 194416 249076
rect 189868 249036 194416 249064
rect 189868 249024 189874 249036
rect 194410 249024 194416 249036
rect 194468 249024 194474 249076
rect 194410 248752 194416 248804
rect 194468 248792 194474 248804
rect 197354 248792 197360 248804
rect 194468 248764 197360 248792
rect 194468 248752 194474 248764
rect 197354 248752 197360 248764
rect 197412 248752 197418 248804
rect 57606 248480 57612 248532
rect 57664 248520 57670 248532
rect 67634 248520 67640 248532
rect 57664 248492 67640 248520
rect 57664 248480 57670 248492
rect 67634 248480 67640 248492
rect 67692 248480 67698 248532
rect 120074 248412 120080 248464
rect 120132 248452 120138 248464
rect 176194 248452 176200 248464
rect 120132 248424 176200 248452
rect 120132 248412 120138 248424
rect 176194 248412 176200 248424
rect 176252 248412 176258 248464
rect 320266 248412 320272 248464
rect 320324 248452 320330 248464
rect 434714 248452 434720 248464
rect 320324 248424 434720 248452
rect 320324 248412 320330 248424
rect 434714 248412 434720 248424
rect 434772 248412 434778 248464
rect 121546 248344 121552 248396
rect 121604 248384 121610 248396
rect 146294 248384 146300 248396
rect 121604 248356 146300 248384
rect 121604 248344 121610 248356
rect 146294 248344 146300 248356
rect 146352 248344 146358 248396
rect 121454 247936 121460 247988
rect 121512 247976 121518 247988
rect 123478 247976 123484 247988
rect 121512 247948 123484 247976
rect 121512 247936 121518 247948
rect 123478 247936 123484 247948
rect 123536 247936 123542 247988
rect 134610 247868 134616 247920
rect 134668 247908 134674 247920
rect 147122 247908 147128 247920
rect 134668 247880 147128 247908
rect 134668 247868 134674 247880
rect 147122 247868 147128 247880
rect 147180 247868 147186 247920
rect 146294 247800 146300 247852
rect 146352 247840 146358 247852
rect 173434 247840 173440 247852
rect 146352 247812 173440 247840
rect 146352 247800 146358 247812
rect 173434 247800 173440 247812
rect 173492 247800 173498 247852
rect 122282 247732 122288 247784
rect 122340 247772 122346 247784
rect 160830 247772 160836 247784
rect 122340 247744 160836 247772
rect 122340 247732 122346 247744
rect 160830 247732 160836 247744
rect 160888 247732 160894 247784
rect 122190 247664 122196 247716
rect 122248 247704 122254 247716
rect 164970 247704 164976 247716
rect 122248 247676 164976 247704
rect 122248 247664 122254 247676
rect 164970 247664 164976 247676
rect 165028 247664 165034 247716
rect 65886 247120 65892 247172
rect 65944 247160 65950 247172
rect 67726 247160 67732 247172
rect 65944 247132 67732 247160
rect 65944 247120 65950 247132
rect 67726 247120 67732 247132
rect 67784 247120 67790 247172
rect 60458 247052 60464 247104
rect 60516 247092 60522 247104
rect 67634 247092 67640 247104
rect 60516 247064 67640 247092
rect 60516 247052 60522 247064
rect 67634 247052 67640 247064
rect 67692 247052 67698 247104
rect 120074 246304 120080 246356
rect 120132 246344 120138 246356
rect 135254 246344 135260 246356
rect 120132 246316 135260 246344
rect 120132 246304 120138 246316
rect 135254 246304 135260 246316
rect 135312 246344 135318 246356
rect 192938 246344 192944 246356
rect 135312 246316 192944 246344
rect 135312 246304 135318 246316
rect 192938 246304 192944 246316
rect 192996 246344 193002 246356
rect 197354 246344 197360 246356
rect 192996 246316 197360 246344
rect 192996 246304 193002 246316
rect 197354 246304 197360 246316
rect 197412 246304 197418 246356
rect 121546 245760 121552 245812
rect 121604 245800 121610 245812
rect 123754 245800 123760 245812
rect 121604 245772 123760 245800
rect 121604 245760 121610 245772
rect 123754 245760 123760 245772
rect 123812 245760 123818 245812
rect 64782 245692 64788 245744
rect 64840 245732 64846 245744
rect 67634 245732 67640 245744
rect 64840 245704 67640 245732
rect 64840 245692 64846 245704
rect 67634 245692 67640 245704
rect 67692 245692 67698 245744
rect 56410 245624 56416 245676
rect 56468 245664 56474 245676
rect 67726 245664 67732 245676
rect 56468 245636 67732 245664
rect 56468 245624 56474 245636
rect 67726 245624 67732 245636
rect 67784 245624 67790 245676
rect 121454 245624 121460 245676
rect 121512 245664 121518 245676
rect 151262 245664 151268 245676
rect 121512 245636 151268 245664
rect 121512 245624 121518 245636
rect 151262 245624 151268 245636
rect 151320 245624 151326 245676
rect 320358 245624 320364 245676
rect 320416 245664 320422 245676
rect 374638 245664 374644 245676
rect 320416 245636 374644 245664
rect 320416 245624 320422 245636
rect 374638 245624 374644 245636
rect 374696 245624 374702 245676
rect 50798 245556 50804 245608
rect 50856 245596 50862 245608
rect 67634 245596 67640 245608
rect 50856 245568 67640 245596
rect 50856 245556 50862 245568
rect 67634 245556 67640 245568
rect 67692 245556 67698 245608
rect 121546 245556 121552 245608
rect 121604 245596 121610 245608
rect 138198 245596 138204 245608
rect 121604 245568 138204 245596
rect 121604 245556 121610 245568
rect 138198 245556 138204 245568
rect 138256 245556 138262 245608
rect 46658 245488 46664 245540
rect 46716 245528 46722 245540
rect 55858 245528 55864 245540
rect 46716 245500 55864 245528
rect 46716 245488 46722 245500
rect 55858 245488 55864 245500
rect 55916 245528 55922 245540
rect 56410 245528 56416 245540
rect 55916 245500 56416 245528
rect 55916 245488 55922 245500
rect 56410 245488 56416 245500
rect 56468 245488 56474 245540
rect 121454 244264 121460 244316
rect 121512 244304 121518 244316
rect 154022 244304 154028 244316
rect 121512 244276 154028 244304
rect 121512 244264 121518 244276
rect 154022 244264 154028 244276
rect 154080 244264 154086 244316
rect 322842 244264 322848 244316
rect 322900 244304 322906 244316
rect 324406 244304 324412 244316
rect 322900 244276 324412 244304
rect 322900 244264 322906 244276
rect 324406 244264 324412 244276
rect 324464 244304 324470 244316
rect 378778 244304 378784 244316
rect 324464 244276 378784 244304
rect 324464 244264 324470 244276
rect 378778 244264 378784 244276
rect 378836 244264 378842 244316
rect 37090 244196 37096 244248
rect 37148 244236 37154 244248
rect 67726 244236 67732 244248
rect 37148 244208 67732 244236
rect 37148 244196 37154 244208
rect 67726 244196 67732 244208
rect 67784 244196 67790 244248
rect 45370 244128 45376 244180
rect 45428 244168 45434 244180
rect 67634 244168 67640 244180
rect 45428 244140 67640 244168
rect 45428 244128 45434 244140
rect 67634 244128 67640 244140
rect 67692 244128 67698 244180
rect 68462 243516 68468 243568
rect 68520 243556 68526 243568
rect 68922 243556 68928 243568
rect 68520 243528 68928 243556
rect 68520 243516 68526 243528
rect 68922 243516 68928 243528
rect 68980 243516 68986 243568
rect 137278 242972 137284 243024
rect 137336 243012 137342 243024
rect 184382 243012 184388 243024
rect 137336 242984 184388 243012
rect 137336 242972 137342 242984
rect 184382 242972 184388 242984
rect 184440 242972 184446 243024
rect 121454 242904 121460 242956
rect 121512 242944 121518 242956
rect 185854 242944 185860 242956
rect 121512 242916 185860 242944
rect 121512 242904 121518 242916
rect 185854 242904 185860 242916
rect 185912 242904 185918 242956
rect 321738 242904 321744 242956
rect 321796 242944 321802 242956
rect 449158 242944 449164 242956
rect 321796 242916 449164 242944
rect 321796 242904 321802 242916
rect 449158 242904 449164 242916
rect 449216 242904 449222 242956
rect 121546 242836 121552 242888
rect 121604 242876 121610 242888
rect 137278 242876 137284 242888
rect 121604 242848 137284 242876
rect 121604 242836 121610 242848
rect 137278 242836 137284 242848
rect 137336 242836 137342 242888
rect 121454 242768 121460 242820
rect 121512 242808 121518 242820
rect 132586 242808 132592 242820
rect 121512 242780 132592 242808
rect 121512 242768 121518 242780
rect 132586 242768 132592 242780
rect 132644 242808 132650 242820
rect 133782 242808 133788 242820
rect 132644 242780 133788 242808
rect 132644 242768 132650 242780
rect 133782 242768 133788 242780
rect 133840 242768 133846 242820
rect 196802 242496 196808 242548
rect 196860 242536 196866 242548
rect 197262 242536 197268 242548
rect 196860 242508 197268 242536
rect 196860 242496 196866 242508
rect 197262 242496 197268 242508
rect 197320 242536 197326 242548
rect 198458 242536 198464 242548
rect 197320 242508 198464 242536
rect 197320 242496 197326 242508
rect 198458 242496 198464 242508
rect 198516 242496 198522 242548
rect 154114 242156 154120 242208
rect 154172 242196 154178 242208
rect 189810 242196 189816 242208
rect 154172 242168 189816 242196
rect 154172 242156 154178 242168
rect 189810 242156 189816 242168
rect 189868 242156 189874 242208
rect 3418 241408 3424 241460
rect 3476 241448 3482 241460
rect 34606 241448 34612 241460
rect 3476 241420 34612 241448
rect 3476 241408 3482 241420
rect 34606 241408 34612 241420
rect 34664 241408 34670 241460
rect 34606 240728 34612 240780
rect 34664 240768 34670 240780
rect 35526 240768 35532 240780
rect 34664 240740 35532 240768
rect 34664 240728 34670 240740
rect 35526 240728 35532 240740
rect 35584 240768 35590 240780
rect 58894 240768 58900 240780
rect 35584 240740 58900 240768
rect 35584 240728 35590 240740
rect 58894 240728 58900 240740
rect 58952 240728 58958 240780
rect 158162 240728 158168 240780
rect 158220 240768 158226 240780
rect 194318 240768 194324 240780
rect 158220 240740 194324 240768
rect 158220 240728 158226 240740
rect 194318 240728 194324 240740
rect 194376 240728 194382 240780
rect 536834 240728 536840 240780
rect 536892 240768 536898 240780
rect 580258 240768 580264 240780
rect 536892 240740 580264 240768
rect 536892 240728 536898 240740
rect 580258 240728 580264 240740
rect 580316 240728 580322 240780
rect 121454 240184 121460 240236
rect 121512 240224 121518 240236
rect 126422 240224 126428 240236
rect 121512 240196 126428 240224
rect 121512 240184 121518 240196
rect 126422 240184 126428 240196
rect 126480 240184 126486 240236
rect 325050 240184 325056 240236
rect 325108 240224 325114 240236
rect 502426 240224 502432 240236
rect 325108 240196 502432 240224
rect 325108 240184 325114 240196
rect 502426 240184 502432 240196
rect 502484 240184 502490 240236
rect 119982 240116 119988 240168
rect 120040 240156 120046 240168
rect 199654 240156 199660 240168
rect 120040 240128 199660 240156
rect 120040 240116 120046 240128
rect 199654 240116 199660 240128
rect 199712 240116 199718 240168
rect 320082 240116 320088 240168
rect 320140 240156 320146 240168
rect 536834 240156 536840 240168
rect 320140 240128 536840 240156
rect 320140 240116 320146 240128
rect 536834 240116 536840 240128
rect 536892 240116 536898 240168
rect 3510 240048 3516 240100
rect 3568 240088 3574 240100
rect 39942 240088 39948 240100
rect 3568 240060 39948 240088
rect 3568 240048 3574 240060
rect 39942 240048 39948 240060
rect 40000 240048 40006 240100
rect 55030 240048 55036 240100
rect 55088 240088 55094 240100
rect 68646 240088 68652 240100
rect 55088 240060 68652 240088
rect 55088 240048 55094 240060
rect 68646 240048 68652 240060
rect 68704 240088 68710 240100
rect 68704 240060 71820 240088
rect 68704 240048 68710 240060
rect 71792 239964 71820 240060
rect 120810 240048 120816 240100
rect 120868 240088 120874 240100
rect 329834 240088 329840 240100
rect 120868 240060 329840 240088
rect 120868 240048 120874 240060
rect 329834 240048 329840 240060
rect 329892 240048 329898 240100
rect 130562 239980 130568 240032
rect 130620 240020 130626 240032
rect 327074 240020 327080 240032
rect 130620 239992 327080 240020
rect 130620 239980 130626 239992
rect 327074 239980 327080 239992
rect 327132 239980 327138 240032
rect 71774 239912 71780 239964
rect 71832 239912 71838 239964
rect 201402 239912 201408 239964
rect 201460 239952 201466 239964
rect 320266 239952 320272 239964
rect 201460 239924 320272 239952
rect 201460 239912 201466 239924
rect 320266 239912 320272 239924
rect 320324 239912 320330 239964
rect 70394 239776 70400 239828
rect 70452 239816 70458 239828
rect 71302 239816 71308 239828
rect 70452 239788 71308 239816
rect 70452 239776 70458 239788
rect 71302 239776 71308 239788
rect 71360 239776 71366 239828
rect 75914 239776 75920 239828
rect 75972 239816 75978 239828
rect 77098 239816 77104 239828
rect 75972 239788 77104 239816
rect 75972 239776 75978 239788
rect 77098 239776 77104 239788
rect 77156 239776 77162 239828
rect 77294 239776 77300 239828
rect 77352 239816 77358 239828
rect 78386 239816 78392 239828
rect 77352 239788 78392 239816
rect 77352 239776 77358 239788
rect 78386 239776 78392 239788
rect 78444 239776 78450 239828
rect 84286 239776 84292 239828
rect 84344 239816 84350 239828
rect 85470 239816 85476 239828
rect 84344 239788 85476 239816
rect 84344 239776 84350 239788
rect 85470 239776 85476 239788
rect 85528 239776 85534 239828
rect 86954 239776 86960 239828
rect 87012 239816 87018 239828
rect 88046 239816 88052 239828
rect 87012 239788 88052 239816
rect 87012 239776 87018 239788
rect 88046 239776 88052 239788
rect 88104 239776 88110 239828
rect 92474 239776 92480 239828
rect 92532 239816 92538 239828
rect 93198 239816 93204 239828
rect 92532 239788 93204 239816
rect 92532 239776 92538 239788
rect 93198 239776 93204 239788
rect 93256 239776 93262 239828
rect 95234 239776 95240 239828
rect 95292 239816 95298 239828
rect 96418 239816 96424 239828
rect 95292 239788 96424 239816
rect 95292 239776 95298 239788
rect 96418 239776 96424 239788
rect 96476 239776 96482 239828
rect 99374 239776 99380 239828
rect 99432 239816 99438 239828
rect 100282 239816 100288 239828
rect 99432 239788 100288 239816
rect 99432 239776 99438 239788
rect 100282 239776 100288 239788
rect 100340 239776 100346 239828
rect 100754 239776 100760 239828
rect 100812 239816 100818 239828
rect 101570 239816 101576 239828
rect 100812 239788 101576 239816
rect 100812 239776 100818 239788
rect 101570 239776 101576 239788
rect 101628 239776 101634 239828
rect 102134 239776 102140 239828
rect 102192 239816 102198 239828
rect 102858 239816 102864 239828
rect 102192 239788 102864 239816
rect 102192 239776 102198 239788
rect 102858 239776 102864 239788
rect 102916 239776 102922 239828
rect 110414 239776 110420 239828
rect 110472 239816 110478 239828
rect 111230 239816 111236 239828
rect 110472 239788 111236 239816
rect 110472 239776 110478 239788
rect 111230 239776 111236 239788
rect 111288 239776 111294 239828
rect 114554 239776 114560 239828
rect 114612 239816 114618 239828
rect 115738 239816 115744 239828
rect 114612 239788 115744 239816
rect 114612 239776 114618 239788
rect 115738 239776 115744 239788
rect 115796 239776 115802 239828
rect 238754 239776 238760 239828
rect 238812 239816 238818 239828
rect 239904 239816 239910 239828
rect 238812 239788 239910 239816
rect 238812 239776 238818 239788
rect 239904 239776 239910 239788
rect 239962 239776 239968 239828
rect 247034 239776 247040 239828
rect 247092 239816 247098 239828
rect 248276 239816 248282 239828
rect 247092 239788 248282 239816
rect 247092 239776 247098 239788
rect 248276 239776 248282 239788
rect 248334 239776 248340 239828
rect 258074 239776 258080 239828
rect 258132 239816 258138 239828
rect 259224 239816 259230 239828
rect 258132 239788 259230 239816
rect 258132 239776 258138 239788
rect 259224 239776 259230 239788
rect 259282 239776 259288 239828
rect 266354 239776 266360 239828
rect 266412 239816 266418 239828
rect 267596 239816 267602 239828
rect 266412 239788 267602 239816
rect 266412 239776 266418 239788
rect 267596 239776 267602 239788
rect 267654 239776 267660 239828
rect 285674 239776 285680 239828
rect 285732 239816 285738 239828
rect 286916 239816 286922 239828
rect 285732 239788 286922 239816
rect 285732 239776 285738 239788
rect 286916 239776 286922 239788
rect 286974 239776 286980 239828
rect 195882 239640 195888 239692
rect 195940 239680 195946 239692
rect 200850 239680 200856 239692
rect 195940 239652 200856 239680
rect 195940 239640 195946 239652
rect 200850 239640 200856 239652
rect 200908 239640 200914 239692
rect 193030 239504 193036 239556
rect 193088 239544 193094 239556
rect 201586 239544 201592 239556
rect 193088 239516 201592 239544
rect 193088 239504 193094 239516
rect 201586 239504 201592 239516
rect 201644 239504 201650 239556
rect 69842 239436 69848 239488
rect 69900 239476 69906 239488
rect 76558 239476 76564 239488
rect 69900 239448 76564 239476
rect 69900 239436 69906 239448
rect 76558 239436 76564 239448
rect 76616 239436 76622 239488
rect 187234 239436 187240 239488
rect 187292 239476 187298 239488
rect 196802 239476 196808 239488
rect 187292 239448 196808 239476
rect 187292 239436 187298 239448
rect 196802 239436 196808 239448
rect 196860 239436 196866 239488
rect 65978 239368 65984 239420
rect 66036 239408 66042 239420
rect 82078 239408 82084 239420
rect 66036 239380 82084 239408
rect 66036 239368 66042 239380
rect 82078 239368 82084 239380
rect 82136 239368 82142 239420
rect 153930 239368 153936 239420
rect 153988 239408 153994 239420
rect 195146 239408 195152 239420
rect 153988 239380 195152 239408
rect 153988 239368 153994 239380
rect 195146 239368 195152 239380
rect 195204 239368 195210 239420
rect 512086 239368 512092 239420
rect 512144 239408 512150 239420
rect 580166 239408 580172 239420
rect 512144 239380 580172 239408
rect 512144 239368 512150 239380
rect 580166 239368 580172 239380
rect 580224 239368 580230 239420
rect 117038 238960 117044 239012
rect 117096 239000 117102 239012
rect 125594 239000 125600 239012
rect 117096 238972 125600 239000
rect 117096 238960 117102 238972
rect 125594 238960 125600 238972
rect 125652 238960 125658 239012
rect 85666 238892 85672 238944
rect 85724 238932 85730 238944
rect 86770 238932 86776 238944
rect 85724 238904 86776 238932
rect 85724 238892 85730 238904
rect 86770 238892 86776 238904
rect 86828 238932 86834 238944
rect 123662 238932 123668 238944
rect 86828 238904 123668 238932
rect 86828 238892 86834 238904
rect 123662 238892 123668 238904
rect 123720 238892 123726 238944
rect 82906 238824 82912 238876
rect 82964 238864 82970 238876
rect 120074 238864 120080 238876
rect 82964 238836 120080 238864
rect 82964 238824 82970 238836
rect 120074 238824 120080 238836
rect 120132 238824 120138 238876
rect 121454 238824 121460 238876
rect 121512 238864 121518 238876
rect 304258 238864 304264 238876
rect 121512 238836 304264 238864
rect 121512 238824 121518 238836
rect 304258 238824 304264 238836
rect 304316 238824 304322 238876
rect 39942 238756 39948 238808
rect 40000 238796 40006 238808
rect 111886 238796 111892 238808
rect 40000 238768 111892 238796
rect 40000 238756 40006 238768
rect 111886 238756 111892 238768
rect 111944 238796 111950 238808
rect 112530 238796 112536 238808
rect 111944 238768 112536 238796
rect 111944 238756 111950 238768
rect 112530 238756 112536 238768
rect 112588 238756 112594 238808
rect 114462 238756 114468 238808
rect 114520 238796 114526 238808
rect 131206 238796 131212 238808
rect 114520 238768 131212 238796
rect 114520 238756 114526 238768
rect 131206 238756 131212 238768
rect 131264 238756 131270 238808
rect 252830 238756 252836 238808
rect 252888 238796 252894 238808
rect 512086 238796 512092 238808
rect 252888 238768 512092 238796
rect 252888 238756 252894 238768
rect 512086 238756 512092 238768
rect 512144 238756 512150 238808
rect 53742 238688 53748 238740
rect 53800 238728 53806 238740
rect 82262 238728 82268 238740
rect 53800 238700 82268 238728
rect 53800 238688 53806 238700
rect 82262 238688 82268 238700
rect 82320 238688 82326 238740
rect 83550 238688 83556 238740
rect 83608 238728 83614 238740
rect 149054 238728 149060 238740
rect 83608 238700 149060 238728
rect 83608 238688 83614 238700
rect 149054 238688 149060 238700
rect 149112 238728 149118 238740
rect 316586 238728 316592 238740
rect 149112 238700 316592 238728
rect 149112 238688 149118 238700
rect 316586 238688 316592 238700
rect 316644 238688 316650 238740
rect 48038 238620 48044 238672
rect 48096 238660 48102 238672
rect 72602 238660 72608 238672
rect 48096 238632 72608 238660
rect 48096 238620 48102 238632
rect 72602 238620 72608 238632
rect 72660 238620 72666 238672
rect 88702 238620 88708 238672
rect 88760 238660 88766 238672
rect 241882 238660 241888 238672
rect 88760 238632 241888 238660
rect 88760 238620 88766 238632
rect 241882 238620 241888 238632
rect 241940 238620 241946 238672
rect 299198 238620 299204 238672
rect 299256 238660 299262 238672
rect 320082 238660 320088 238672
rect 299256 238632 320088 238660
rect 299256 238620 299262 238632
rect 320082 238620 320088 238632
rect 320140 238620 320146 238672
rect 118326 238552 118332 238604
rect 118384 238592 118390 238604
rect 143534 238592 143540 238604
rect 118384 238564 143540 238592
rect 118384 238552 118390 238564
rect 143534 238552 143540 238564
rect 143592 238552 143598 238604
rect 304258 238552 304264 238604
rect 304316 238592 304322 238604
rect 312078 238592 312084 238604
rect 304316 238564 312084 238592
rect 304316 238552 304322 238564
rect 312078 238552 312084 238564
rect 312136 238552 312142 238604
rect 115106 238484 115112 238536
rect 115164 238524 115170 238536
rect 144914 238524 144920 238536
rect 115164 238496 144920 238524
rect 115164 238484 115170 238496
rect 144914 238484 144920 238496
rect 144972 238484 144978 238536
rect 69934 238416 69940 238468
rect 69992 238456 69998 238468
rect 119982 238456 119988 238468
rect 69992 238428 119988 238456
rect 69992 238416 69998 238428
rect 119982 238416 119988 238428
rect 120040 238416 120046 238468
rect 71958 238144 71964 238196
rect 72016 238184 72022 238196
rect 78858 238184 78864 238196
rect 72016 238156 78864 238184
rect 72016 238144 72022 238156
rect 78858 238144 78864 238156
rect 78916 238144 78922 238196
rect 194318 238144 194324 238196
rect 194376 238184 194382 238196
rect 204162 238184 204168 238196
rect 194376 238156 204168 238184
rect 194376 238144 194382 238156
rect 204162 238144 204168 238156
rect 204220 238144 204226 238196
rect 60366 238076 60372 238128
rect 60424 238116 60430 238128
rect 72418 238116 72424 238128
rect 60424 238088 72424 238116
rect 60424 238076 60430 238088
rect 72418 238076 72424 238088
rect 72476 238076 72482 238128
rect 73246 238076 73252 238128
rect 73304 238116 73310 238128
rect 83458 238116 83464 238128
rect 73304 238088 83464 238116
rect 73304 238076 73310 238088
rect 83458 238076 83464 238088
rect 83516 238076 83522 238128
rect 159634 238076 159640 238128
rect 159692 238116 159698 238128
rect 201402 238116 201408 238128
rect 159692 238088 201408 238116
rect 159692 238076 159698 238088
rect 201402 238076 201408 238088
rect 201460 238076 201466 238128
rect 314102 238076 314108 238128
rect 314160 238116 314166 238128
rect 320358 238116 320364 238128
rect 314160 238088 320364 238116
rect 314160 238076 314166 238088
rect 320358 238076 320364 238088
rect 320416 238076 320422 238128
rect 64782 238008 64788 238060
rect 64840 238048 64846 238060
rect 88978 238048 88984 238060
rect 64840 238020 88984 238048
rect 64840 238008 64846 238020
rect 88978 238008 88984 238020
rect 89036 238008 89042 238060
rect 155494 238008 155500 238060
rect 155552 238048 155558 238060
rect 204990 238048 204996 238060
rect 155552 238020 204996 238048
rect 155552 238008 155558 238020
rect 204990 238008 204996 238020
rect 205048 238008 205054 238060
rect 316586 238008 316592 238060
rect 316644 238048 316650 238060
rect 438854 238048 438860 238060
rect 316644 238020 438860 238048
rect 316644 238008 316650 238020
rect 438854 238008 438860 238020
rect 438912 238008 438918 238060
rect 323670 237464 323676 237516
rect 323728 237504 323734 237516
rect 332962 237504 332968 237516
rect 323728 237476 332968 237504
rect 323728 237464 323734 237476
rect 332962 237464 332968 237476
rect 333020 237464 333026 237516
rect 80974 237396 80980 237448
rect 81032 237436 81038 237448
rect 86218 237436 86224 237448
rect 81032 237408 86224 237436
rect 81032 237396 81038 237408
rect 86218 237396 86224 237408
rect 86276 237396 86282 237448
rect 199930 237396 199936 237448
rect 199988 237436 199994 237448
rect 202322 237436 202328 237448
rect 199988 237408 202328 237436
rect 199988 237396 199994 237408
rect 202322 237396 202328 237408
rect 202380 237396 202386 237448
rect 218698 237396 218704 237448
rect 218756 237436 218762 237448
rect 220630 237436 220636 237448
rect 218756 237408 220636 237436
rect 218756 237396 218762 237408
rect 220630 237396 220636 237408
rect 220688 237396 220694 237448
rect 228542 237396 228548 237448
rect 228600 237436 228606 237448
rect 229646 237436 229652 237448
rect 228600 237408 229652 237436
rect 228600 237396 228606 237408
rect 229646 237396 229652 237408
rect 229704 237396 229710 237448
rect 235258 237396 235264 237448
rect 235316 237436 235322 237448
rect 236086 237436 236092 237448
rect 235316 237408 236092 237436
rect 235316 237396 235322 237408
rect 236086 237396 236092 237408
rect 236144 237396 236150 237448
rect 244918 237396 244924 237448
rect 244976 237436 244982 237448
rect 246390 237436 246396 237448
rect 244976 237408 246396 237436
rect 244976 237396 244982 237408
rect 246390 237396 246396 237408
rect 246448 237396 246454 237448
rect 251634 237396 251640 237448
rect 251692 237436 251698 237448
rect 254762 237436 254768 237448
rect 251692 237408 254768 237436
rect 251692 237396 251698 237408
rect 254762 237396 254768 237408
rect 254820 237396 254826 237448
rect 283558 237396 283564 237448
rect 283616 237436 283622 237448
rect 284386 237436 284392 237448
rect 283616 237408 284392 237436
rect 283616 237396 283622 237408
rect 284386 237396 284392 237408
rect 284444 237396 284450 237448
rect 312078 237396 312084 237448
rect 312136 237436 312142 237448
rect 312538 237436 312544 237448
rect 312136 237408 312544 237436
rect 312136 237396 312142 237408
rect 312538 237396 312544 237408
rect 312596 237396 312602 237448
rect 318058 237396 318064 237448
rect 318116 237436 318122 237448
rect 318518 237436 318524 237448
rect 318116 237408 318524 237436
rect 318116 237396 318122 237408
rect 318518 237396 318524 237408
rect 318576 237436 318582 237448
rect 498286 237436 498292 237448
rect 318576 237408 498292 237436
rect 318576 237396 318582 237408
rect 498286 237396 498292 237408
rect 498344 237396 498350 237448
rect 57882 237328 57888 237380
rect 57940 237368 57946 237380
rect 86126 237368 86132 237380
rect 57940 237340 86132 237368
rect 57940 237328 57946 237340
rect 86126 237328 86132 237340
rect 86184 237328 86190 237380
rect 128262 237328 128268 237380
rect 128320 237368 128326 237380
rect 322198 237368 322204 237380
rect 128320 237340 322204 237368
rect 128320 237328 128326 237340
rect 322198 237328 322204 237340
rect 322256 237328 322262 237380
rect 107378 237260 107384 237312
rect 107436 237300 107442 237312
rect 132494 237300 132500 237312
rect 107436 237272 132500 237300
rect 107436 237260 107442 237272
rect 132494 237260 132500 237272
rect 132552 237260 132558 237312
rect 162394 237260 162400 237312
rect 162452 237300 162458 237312
rect 332594 237300 332600 237312
rect 162452 237272 332600 237300
rect 162452 237260 162458 237272
rect 332594 237260 332600 237272
rect 332652 237260 332658 237312
rect 95786 237192 95792 237244
rect 95844 237232 95850 237244
rect 128354 237232 128360 237244
rect 95844 237204 128360 237232
rect 95844 237192 95850 237204
rect 128354 237192 128360 237204
rect 128412 237192 128418 237244
rect 166534 237192 166540 237244
rect 166592 237232 166598 237244
rect 319346 237232 319352 237244
rect 166592 237204 319352 237232
rect 166592 237192 166598 237204
rect 319346 237192 319352 237204
rect 319404 237192 319410 237244
rect 201402 237124 201408 237176
rect 201460 237164 201466 237176
rect 303706 237164 303712 237176
rect 201460 237136 303712 237164
rect 201460 237124 201466 237136
rect 303706 237124 303712 237136
rect 303764 237124 303770 237176
rect 181622 237056 181628 237108
rect 181680 237096 181686 237108
rect 276014 237096 276020 237108
rect 181680 237068 276020 237096
rect 181680 237056 181686 237068
rect 276014 237056 276020 237068
rect 276072 237056 276078 237108
rect 195146 236988 195152 237040
rect 195204 237028 195210 237040
rect 210418 237028 210424 237040
rect 195204 237000 210424 237028
rect 195204 236988 195210 237000
rect 210418 236988 210424 237000
rect 210476 236988 210482 237040
rect 276014 235968 276020 236020
rect 276072 236008 276078 236020
rect 276658 236008 276664 236020
rect 276072 235980 276664 236008
rect 276072 235968 276078 235980
rect 276658 235968 276664 235980
rect 276716 235968 276722 236020
rect 303706 235968 303712 236020
rect 303764 236008 303770 236020
rect 304258 236008 304264 236020
rect 303764 235980 304264 236008
rect 303764 235968 303770 235980
rect 304258 235968 304264 235980
rect 304316 235968 304322 236020
rect 326982 235968 326988 236020
rect 327040 236008 327046 236020
rect 349154 236008 349160 236020
rect 327040 235980 349160 236008
rect 327040 235968 327046 235980
rect 349154 235968 349160 235980
rect 349212 235968 349218 236020
rect 48222 235900 48228 235952
rect 48280 235940 48286 235952
rect 98362 235940 98368 235952
rect 48280 235912 98368 235940
rect 48280 235900 48286 235912
rect 98362 235900 98368 235912
rect 98420 235900 98426 235952
rect 106090 235900 106096 235952
rect 106148 235940 106154 235952
rect 173342 235940 173348 235952
rect 106148 235912 173348 235940
rect 106148 235900 106154 235912
rect 173342 235900 173348 235912
rect 173400 235900 173406 235952
rect 195698 235900 195704 235952
rect 195756 235940 195762 235952
rect 504358 235940 504364 235952
rect 195756 235912 504364 235940
rect 195756 235900 195762 235912
rect 504358 235900 504364 235912
rect 504416 235900 504422 235952
rect 54478 235832 54484 235884
rect 54536 235872 54542 235884
rect 85666 235872 85672 235884
rect 54536 235844 85672 235872
rect 54536 235832 54542 235844
rect 85666 235832 85672 235844
rect 85724 235832 85730 235884
rect 89346 235832 89352 235884
rect 89404 235872 89410 235884
rect 142246 235872 142252 235884
rect 89404 235844 142252 235872
rect 89404 235832 89410 235844
rect 142246 235832 142252 235844
rect 142304 235832 142310 235884
rect 149790 235832 149796 235884
rect 149848 235872 149854 235884
rect 321554 235872 321560 235884
rect 149848 235844 321560 235872
rect 149848 235832 149854 235844
rect 321554 235832 321560 235844
rect 321612 235832 321618 235884
rect 97718 235764 97724 235816
rect 97776 235804 97782 235816
rect 251634 235804 251640 235816
rect 97776 235776 251640 235804
rect 97776 235764 97782 235776
rect 251634 235764 251640 235776
rect 251692 235764 251698 235816
rect 58894 235696 58900 235748
rect 58952 235736 58958 235748
rect 103514 235736 103520 235748
rect 58952 235708 103520 235736
rect 58952 235696 58958 235708
rect 103514 235696 103520 235708
rect 103572 235696 103578 235748
rect 113818 235696 113824 235748
rect 113876 235736 113882 235748
rect 131758 235736 131764 235748
rect 113876 235708 131764 235736
rect 113876 235696 113882 235708
rect 131758 235696 131764 235708
rect 131816 235696 131822 235748
rect 165062 235696 165068 235748
rect 165120 235736 165126 235748
rect 301498 235736 301504 235748
rect 165120 235708 301504 235736
rect 165120 235696 165126 235708
rect 301498 235696 301504 235708
rect 301556 235696 301562 235748
rect 91278 235628 91284 235680
rect 91336 235668 91342 235680
rect 124950 235668 124956 235680
rect 91336 235640 124956 235668
rect 91336 235628 91342 235640
rect 124950 235628 124956 235640
rect 125008 235628 125014 235680
rect 191190 235628 191196 235680
rect 191248 235668 191254 235680
rect 326338 235668 326344 235680
rect 191248 235640 326344 235668
rect 191248 235628 191254 235640
rect 326338 235628 326344 235640
rect 326396 235668 326402 235680
rect 326982 235668 326988 235680
rect 326396 235640 326988 235668
rect 326396 235628 326402 235640
rect 326982 235628 326988 235640
rect 327040 235628 327046 235680
rect 118602 235560 118608 235612
rect 118660 235600 118666 235612
rect 129734 235600 129740 235612
rect 118660 235572 129740 235600
rect 118660 235560 118666 235572
rect 129734 235560 129740 235572
rect 129792 235560 129798 235612
rect 185762 235220 185768 235272
rect 185820 235260 185826 235272
rect 268378 235260 268384 235272
rect 185820 235232 268384 235260
rect 185820 235220 185826 235232
rect 268378 235220 268384 235232
rect 268436 235220 268442 235272
rect 503714 234948 503720 235000
rect 503772 234988 503778 235000
rect 504358 234988 504364 235000
rect 503772 234960 504364 234988
rect 503772 234948 503778 234960
rect 504358 234948 504364 234960
rect 504416 234948 504422 235000
rect 117682 234676 117688 234728
rect 117740 234716 117746 234728
rect 118602 234716 118608 234728
rect 117740 234688 118608 234716
rect 117740 234676 117746 234688
rect 118602 234676 118608 234688
rect 118660 234676 118666 234728
rect 321554 234676 321560 234728
rect 321612 234716 321618 234728
rect 322198 234716 322204 234728
rect 321612 234688 322204 234716
rect 321612 234676 321618 234688
rect 322198 234676 322204 234688
rect 322256 234676 322262 234728
rect 288894 234608 288900 234660
rect 288952 234648 288958 234660
rect 289446 234648 289452 234660
rect 288952 234620 289452 234648
rect 288952 234608 288958 234620
rect 289446 234608 289452 234620
rect 289504 234648 289510 234660
rect 432598 234648 432604 234660
rect 289504 234620 432604 234648
rect 289504 234608 289510 234620
rect 432598 234608 432604 234620
rect 432656 234608 432662 234660
rect 61746 234540 61752 234592
rect 61804 234580 61810 234592
rect 256694 234580 256700 234592
rect 61804 234552 256700 234580
rect 61804 234540 61810 234552
rect 256694 234540 256700 234552
rect 256752 234540 256758 234592
rect 50890 234472 50896 234524
rect 50948 234512 50954 234524
rect 91738 234512 91744 234524
rect 50948 234484 91744 234512
rect 50948 234472 50954 234484
rect 91738 234472 91744 234484
rect 91796 234472 91802 234524
rect 95142 234472 95148 234524
rect 95200 234512 95206 234524
rect 170582 234512 170588 234524
rect 95200 234484 170588 234512
rect 95200 234472 95206 234484
rect 170582 234472 170588 234484
rect 170640 234472 170646 234524
rect 81618 234404 81624 234456
rect 81676 234444 81682 234456
rect 123570 234444 123576 234456
rect 81676 234416 123576 234444
rect 81676 234404 81682 234416
rect 123570 234404 123576 234416
rect 123628 234404 123634 234456
rect 151354 234404 151360 234456
rect 151412 234444 151418 234456
rect 211798 234444 211804 234456
rect 151412 234416 211804 234444
rect 151412 234404 151418 234416
rect 211798 234404 211804 234416
rect 211856 234444 211862 234456
rect 212258 234444 212264 234456
rect 211856 234416 212264 234444
rect 211856 234404 211862 234416
rect 212258 234404 212264 234416
rect 212316 234404 212322 234456
rect 106734 234336 106740 234388
rect 106792 234376 106798 234388
rect 140038 234376 140044 234388
rect 106792 234348 140044 234376
rect 106792 234336 106798 234348
rect 140038 234336 140044 234348
rect 140096 234336 140102 234388
rect 256694 234132 256700 234184
rect 256752 234172 256758 234184
rect 257338 234172 257344 234184
rect 256752 234144 257344 234172
rect 256752 234132 256758 234144
rect 257338 234132 257344 234144
rect 257396 234132 257402 234184
rect 196710 233996 196716 234048
rect 196768 234036 196774 234048
rect 224218 234036 224224 234048
rect 196768 234008 224224 234036
rect 196768 233996 196774 234008
rect 224218 233996 224224 234008
rect 224276 233996 224282 234048
rect 84194 233928 84200 233980
rect 84252 233968 84258 233980
rect 84252 233940 84332 233968
rect 84252 233928 84258 233940
rect 74534 233860 74540 233912
rect 74592 233900 74598 233912
rect 75178 233900 75184 233912
rect 74592 233872 75184 233900
rect 74592 233860 74598 233872
rect 75178 233860 75184 233872
rect 75236 233860 75242 233912
rect 84304 233776 84332 233940
rect 171962 233928 171968 233980
rect 172020 233968 172026 233980
rect 228358 233968 228364 233980
rect 172020 233940 228364 233968
rect 172020 233928 172026 233940
rect 228358 233928 228364 233940
rect 228416 233928 228422 233980
rect 318702 233968 318708 233980
rect 316006 233940 318708 233968
rect 118694 233860 118700 233912
rect 118752 233900 118758 233912
rect 119706 233900 119712 233912
rect 118752 233872 119712 233900
rect 118752 233860 118758 233872
rect 119706 233860 119712 233872
rect 119764 233860 119770 233912
rect 188614 233860 188620 233912
rect 188672 233900 188678 233912
rect 316006 233900 316034 233940
rect 318702 233928 318708 233940
rect 318760 233968 318766 233980
rect 321646 233968 321652 233980
rect 318760 233940 321652 233968
rect 318760 233928 318766 233940
rect 321646 233928 321652 233940
rect 321704 233928 321710 233980
rect 188672 233872 316034 233900
rect 188672 233860 188678 233872
rect 316678 233860 316684 233912
rect 316736 233900 316742 233912
rect 319254 233900 319260 233912
rect 316736 233872 319260 233900
rect 316736 233860 316742 233872
rect 319254 233860 319260 233872
rect 319312 233860 319318 233912
rect 84286 233724 84292 233776
rect 84344 233724 84350 233776
rect 205634 233248 205640 233300
rect 205692 233288 205698 233300
rect 205818 233288 205824 233300
rect 205692 233260 205824 233288
rect 205692 233248 205698 233260
rect 205818 233248 205824 233260
rect 205876 233288 205882 233300
rect 307018 233288 307024 233300
rect 205876 233260 307024 233288
rect 205876 233248 205882 233260
rect 307018 233248 307024 233260
rect 307076 233248 307082 233300
rect 56318 233180 56324 233232
rect 56376 233220 56382 233232
rect 324406 233220 324412 233232
rect 56376 233192 324412 233220
rect 56376 233180 56382 233192
rect 324406 233180 324412 233192
rect 324464 233180 324470 233232
rect 161014 233112 161020 233164
rect 161072 233152 161078 233164
rect 325878 233152 325884 233164
rect 161072 233124 325884 233152
rect 161072 233112 161078 233124
rect 325878 233112 325884 233124
rect 325936 233152 325942 233164
rect 333974 233152 333980 233164
rect 325936 233124 333980 233152
rect 325936 233112 325942 233124
rect 333974 233112 333980 233124
rect 334032 233112 334038 233164
rect 53558 233044 53564 233096
rect 53616 233084 53622 233096
rect 176102 233084 176108 233096
rect 53616 233056 176108 233084
rect 53616 233044 53622 233056
rect 176102 233044 176108 233056
rect 176160 233044 176166 233096
rect 189810 233044 189816 233096
rect 189868 233084 189874 233096
rect 331306 233084 331312 233096
rect 189868 233056 331312 233084
rect 189868 233044 189874 233056
rect 331306 233044 331312 233056
rect 331364 233044 331370 233096
rect 155402 232976 155408 233028
rect 155460 233016 155466 233028
rect 218790 233016 218796 233028
rect 155460 232988 218796 233016
rect 155460 232976 155466 232988
rect 218790 232976 218796 232988
rect 218848 232976 218854 233028
rect 183370 232568 183376 232620
rect 183428 232608 183434 232620
rect 206462 232608 206468 232620
rect 183428 232580 206468 232608
rect 183428 232568 183434 232580
rect 206462 232568 206468 232580
rect 206520 232568 206526 232620
rect 67358 232500 67364 232552
rect 67416 232540 67422 232552
rect 106918 232540 106924 232552
rect 67416 232512 106924 232540
rect 67416 232500 67422 232512
rect 106918 232500 106924 232512
rect 106976 232500 106982 232552
rect 198826 232500 198832 232552
rect 198884 232540 198890 232552
rect 324406 232540 324412 232552
rect 198884 232512 324412 232540
rect 198884 232500 198890 232512
rect 324406 232500 324412 232512
rect 324464 232500 324470 232552
rect 418798 231820 418804 231872
rect 418856 231860 418862 231872
rect 580166 231860 580172 231872
rect 418856 231832 580172 231860
rect 418856 231820 418862 231832
rect 580166 231820 580172 231832
rect 580224 231820 580230 231872
rect 99466 231752 99472 231804
rect 99524 231792 99530 231804
rect 269114 231792 269120 231804
rect 99524 231764 269120 231792
rect 99524 231752 99530 231764
rect 269114 231752 269120 231764
rect 269172 231792 269178 231804
rect 269758 231792 269764 231804
rect 269172 231764 269764 231792
rect 269172 231752 269178 231764
rect 269758 231752 269764 231764
rect 269816 231752 269822 231804
rect 54938 231684 54944 231736
rect 54996 231724 55002 231736
rect 205634 231724 205640 231736
rect 54996 231696 205640 231724
rect 54996 231684 55002 231696
rect 205634 231684 205640 231696
rect 205692 231684 205698 231736
rect 109862 231616 109868 231668
rect 109920 231656 109926 231668
rect 136634 231656 136640 231668
rect 109920 231628 136640 231656
rect 109920 231616 109926 231628
rect 136634 231616 136640 231628
rect 136692 231616 136698 231668
rect 204162 231616 204168 231668
rect 204220 231656 204226 231668
rect 329926 231656 329932 231668
rect 204220 231628 329932 231656
rect 204220 231616 204226 231628
rect 329926 231616 329932 231628
rect 329984 231616 329990 231668
rect 152458 231548 152464 231600
rect 152516 231588 152522 231600
rect 277394 231588 277400 231600
rect 152516 231560 277400 231588
rect 152516 231548 152522 231560
rect 277394 231548 277400 231560
rect 277452 231588 277458 231600
rect 278038 231588 278044 231600
rect 277452 231560 278044 231588
rect 277452 231548 277458 231560
rect 278038 231548 278044 231560
rect 278096 231548 278102 231600
rect 182910 231480 182916 231532
rect 182968 231520 182974 231532
rect 244918 231520 244924 231532
rect 182968 231492 244924 231520
rect 182968 231480 182974 231492
rect 244918 231480 244924 231492
rect 244976 231480 244982 231532
rect 69198 231140 69204 231192
rect 69256 231180 69262 231192
rect 104158 231180 104164 231192
rect 69256 231152 104164 231180
rect 69256 231140 69262 231152
rect 104158 231140 104164 231152
rect 104216 231140 104222 231192
rect 103606 231072 103612 231124
rect 103664 231112 103670 231124
rect 190178 231112 190184 231124
rect 103664 231084 190184 231112
rect 103664 231072 103670 231084
rect 190178 231072 190184 231084
rect 190236 231112 190242 231124
rect 191282 231112 191288 231124
rect 190236 231084 191288 231112
rect 190236 231072 190242 231084
rect 191282 231072 191288 231084
rect 191340 231072 191346 231124
rect 192478 231072 192484 231124
rect 192536 231112 192542 231124
rect 226978 231112 226984 231124
rect 192536 231084 226984 231112
rect 192536 231072 192542 231084
rect 226978 231072 226984 231084
rect 227036 231072 227042 231124
rect 76006 230392 76012 230444
rect 76064 230432 76070 230444
rect 126974 230432 126980 230444
rect 76064 230404 126980 230432
rect 76064 230392 76070 230404
rect 126974 230392 126980 230404
rect 127032 230432 127038 230444
rect 280154 230432 280160 230444
rect 127032 230404 280160 230432
rect 127032 230392 127038 230404
rect 280154 230392 280160 230404
rect 280212 230432 280218 230444
rect 281442 230432 281448 230444
rect 280212 230404 281448 230432
rect 280212 230392 280218 230404
rect 281442 230392 281448 230404
rect 281500 230392 281506 230444
rect 78858 230324 78864 230376
rect 78916 230364 78922 230376
rect 202874 230364 202880 230376
rect 78916 230336 202880 230364
rect 78916 230324 78922 230336
rect 202874 230324 202880 230336
rect 202932 230364 202938 230376
rect 203518 230364 203524 230376
rect 202932 230336 203524 230364
rect 202932 230324 202938 230336
rect 203518 230324 203524 230336
rect 203576 230324 203582 230376
rect 211614 230324 211620 230376
rect 211672 230364 211678 230376
rect 327166 230364 327172 230376
rect 211672 230336 327172 230364
rect 211672 230324 211678 230336
rect 327166 230324 327172 230336
rect 327224 230364 327230 230376
rect 328362 230364 328368 230376
rect 327224 230336 328368 230364
rect 327224 230324 327230 230336
rect 328362 230324 328368 230336
rect 328420 230324 328426 230376
rect 188522 229916 188528 229968
rect 188580 229956 188586 229968
rect 213362 229956 213368 229968
rect 188580 229928 213368 229956
rect 188580 229916 188586 229928
rect 213362 229916 213368 229928
rect 213420 229916 213426 229968
rect 61838 229848 61844 229900
rect 61896 229888 61902 229900
rect 119338 229888 119344 229900
rect 61896 229860 119344 229888
rect 61896 229848 61902 229860
rect 119338 229848 119344 229860
rect 119396 229848 119402 229900
rect 196618 229848 196624 229900
rect 196676 229888 196682 229900
rect 233878 229888 233884 229900
rect 196676 229860 233884 229888
rect 196676 229848 196682 229860
rect 233878 229848 233884 229860
rect 233936 229848 233942 229900
rect 111886 229780 111892 229832
rect 111944 229820 111950 229832
rect 262858 229820 262864 229832
rect 111944 229792 262864 229820
rect 111944 229780 111950 229792
rect 262858 229780 262864 229792
rect 262916 229780 262922 229832
rect 328362 229780 328368 229832
rect 328420 229820 328426 229832
rect 340966 229820 340972 229832
rect 328420 229792 340972 229820
rect 328420 229780 328426 229792
rect 340966 229780 340972 229792
rect 341024 229780 341030 229832
rect 4798 229712 4804 229764
rect 4856 229752 4862 229764
rect 83550 229752 83556 229764
rect 4856 229724 83556 229752
rect 4856 229712 4862 229724
rect 83550 229712 83556 229724
rect 83608 229712 83614 229764
rect 90542 229712 90548 229764
rect 90600 229752 90606 229764
rect 255590 229752 255596 229764
rect 90600 229724 255596 229752
rect 90600 229712 90606 229724
rect 255590 229712 255596 229724
rect 255648 229712 255654 229764
rect 281442 229712 281448 229764
rect 281500 229752 281506 229764
rect 334710 229752 334716 229764
rect 281500 229724 334716 229752
rect 281500 229712 281506 229724
rect 334710 229712 334716 229724
rect 334768 229712 334774 229764
rect 43806 229032 43812 229084
rect 43864 229072 43870 229084
rect 327350 229072 327356 229084
rect 43864 229044 327356 229072
rect 43864 229032 43870 229044
rect 327350 229032 327356 229044
rect 327408 229032 327414 229084
rect 118786 228964 118792 229016
rect 118844 229004 118850 229016
rect 143442 229004 143448 229016
rect 118844 228976 143448 229004
rect 118844 228964 118850 228976
rect 143442 228964 143448 228976
rect 143500 228964 143506 229016
rect 173434 228964 173440 229016
rect 173492 229004 173498 229016
rect 324314 229004 324320 229016
rect 173492 228976 324320 229004
rect 173492 228964 173498 228976
rect 324314 228964 324320 228976
rect 324372 228964 324378 229016
rect 77386 228896 77392 228948
rect 77444 228936 77450 228948
rect 216674 228936 216680 228948
rect 77444 228908 216680 228936
rect 77444 228896 77450 228908
rect 216674 228896 216680 228908
rect 216732 228896 216738 228948
rect 185854 228828 185860 228880
rect 185912 228868 185918 228880
rect 321646 228868 321652 228880
rect 185912 228840 321652 228868
rect 185912 228828 185918 228840
rect 321646 228828 321652 228840
rect 321704 228828 321710 228880
rect 162210 228760 162216 228812
rect 162268 228800 162274 228812
rect 262214 228800 262220 228812
rect 162268 228772 262220 228800
rect 162268 228760 162274 228772
rect 262214 228760 262220 228772
rect 262272 228760 262278 228812
rect 59078 228420 59084 228472
rect 59136 228460 59142 228472
rect 166350 228460 166356 228472
rect 59136 228432 166356 228460
rect 59136 228420 59142 228432
rect 166350 228420 166356 228432
rect 166408 228420 166414 228472
rect 327350 228420 327356 228472
rect 327408 228460 327414 228472
rect 343726 228460 343732 228472
rect 327408 228432 343732 228460
rect 327408 228420 327414 228432
rect 343726 228420 343732 228432
rect 343784 228420 343790 228472
rect 143442 228352 143448 228404
rect 143500 228392 143506 228404
rect 495618 228392 495624 228404
rect 143500 228364 495624 228392
rect 143500 228352 143506 228364
rect 495618 228352 495624 228364
rect 495676 228352 495682 228404
rect 216674 227740 216680 227792
rect 216732 227780 216738 227792
rect 217318 227780 217324 227792
rect 216732 227752 217324 227780
rect 216732 227740 216738 227752
rect 217318 227740 217324 227752
rect 217376 227740 217382 227792
rect 262214 227740 262220 227792
rect 262272 227780 262278 227792
rect 262950 227780 262956 227792
rect 262272 227752 262956 227780
rect 262272 227740 262278 227752
rect 262950 227740 262956 227752
rect 263008 227740 263014 227792
rect 110506 227672 110512 227724
rect 110564 227712 110570 227724
rect 140774 227712 140780 227724
rect 110564 227684 140780 227712
rect 110564 227672 110570 227684
rect 140774 227672 140780 227684
rect 140832 227712 140838 227724
rect 140832 227684 142154 227712
rect 140832 227672 140838 227684
rect 142126 227644 142154 227684
rect 170490 227672 170496 227724
rect 170548 227712 170554 227724
rect 418798 227712 418804 227724
rect 170548 227684 418804 227712
rect 170548 227672 170554 227684
rect 418798 227672 418804 227684
rect 418856 227672 418862 227724
rect 335998 227644 336004 227656
rect 142126 227616 336004 227644
rect 335998 227604 336004 227616
rect 336056 227604 336062 227656
rect 87046 227536 87052 227588
rect 87104 227576 87110 227588
rect 235258 227576 235264 227588
rect 87104 227548 235264 227576
rect 87104 227536 87110 227548
rect 235258 227536 235264 227548
rect 235316 227536 235322 227588
rect 204990 227468 204996 227520
rect 205048 227508 205054 227520
rect 330018 227508 330024 227520
rect 205048 227480 330024 227508
rect 205048 227468 205054 227480
rect 330018 227468 330024 227480
rect 330076 227468 330082 227520
rect 190178 227060 190184 227112
rect 190236 227100 190242 227112
rect 202230 227100 202236 227112
rect 190236 227072 202236 227100
rect 190236 227060 190242 227072
rect 202230 227060 202236 227072
rect 202288 227060 202294 227112
rect 96614 226992 96620 227044
rect 96672 227032 96678 227044
rect 252830 227032 252836 227044
rect 96672 227004 252836 227032
rect 96672 226992 96678 227004
rect 252830 226992 252836 227004
rect 252888 226992 252894 227044
rect 305638 226992 305644 227044
rect 305696 227032 305702 227044
rect 340230 227032 340236 227044
rect 305696 227004 340236 227032
rect 305696 226992 305702 227004
rect 340230 226992 340236 227004
rect 340288 226992 340294 227044
rect 110506 226312 110512 226364
rect 110564 226352 110570 226364
rect 111058 226352 111064 226364
rect 110564 226324 111064 226352
rect 110564 226312 110570 226324
rect 111058 226312 111064 226324
rect 111116 226312 111122 226364
rect 80054 226244 80060 226296
rect 80112 226284 80118 226296
rect 222194 226284 222200 226296
rect 80112 226256 222200 226284
rect 80112 226244 80118 226256
rect 222194 226244 222200 226256
rect 222252 226244 222258 226296
rect 155310 226176 155316 226228
rect 155368 226216 155374 226228
rect 289814 226216 289820 226228
rect 155368 226188 289820 226216
rect 155368 226176 155374 226188
rect 289814 226176 289820 226188
rect 289872 226176 289878 226228
rect 74626 226108 74632 226160
rect 74684 226148 74690 226160
rect 201586 226148 201592 226160
rect 74684 226120 201592 226148
rect 74684 226108 74690 226120
rect 201586 226108 201592 226120
rect 201644 226148 201650 226160
rect 202782 226148 202788 226160
rect 201644 226120 202788 226148
rect 201644 226108 201650 226120
rect 202782 226108 202788 226120
rect 202840 226108 202846 226160
rect 194410 225768 194416 225820
rect 194468 225808 194474 225820
rect 213270 225808 213276 225820
rect 194468 225780 213276 225808
rect 194468 225768 194474 225780
rect 213270 225768 213276 225780
rect 213328 225768 213334 225820
rect 196802 225700 196808 225752
rect 196860 225740 196866 225752
rect 314010 225740 314016 225752
rect 196860 225712 314016 225740
rect 196860 225700 196866 225712
rect 314010 225700 314016 225712
rect 314068 225700 314074 225752
rect 202782 225632 202788 225684
rect 202840 225672 202846 225684
rect 342254 225672 342260 225684
rect 202840 225644 342260 225672
rect 202840 225632 202846 225644
rect 342254 225632 342260 225644
rect 342312 225632 342318 225684
rect 3418 225564 3424 225616
rect 3476 225604 3482 225616
rect 120166 225604 120172 225616
rect 3476 225576 120172 225604
rect 3476 225564 3482 225576
rect 120166 225564 120172 225576
rect 120224 225564 120230 225616
rect 210418 225564 210424 225616
rect 210476 225604 210482 225616
rect 485038 225604 485044 225616
rect 210476 225576 485044 225604
rect 210476 225564 210482 225576
rect 485038 225564 485044 225576
rect 485096 225564 485102 225616
rect 222194 224952 222200 225004
rect 222252 224992 222258 225004
rect 222930 224992 222936 225004
rect 222252 224964 222936 224992
rect 222252 224952 222258 224964
rect 222930 224952 222936 224964
rect 222988 224952 222994 225004
rect 289814 224952 289820 225004
rect 289872 224992 289878 225004
rect 290458 224992 290464 225004
rect 289872 224964 290464 224992
rect 289872 224952 289878 224964
rect 290458 224952 290464 224964
rect 290516 224952 290522 225004
rect 52086 224884 52092 224936
rect 52144 224924 52150 224936
rect 318058 224924 318064 224936
rect 52144 224896 318064 224924
rect 52144 224884 52150 224896
rect 318058 224884 318064 224896
rect 318116 224884 318122 224936
rect 55858 224816 55864 224868
rect 55916 224856 55922 224868
rect 258074 224856 258080 224868
rect 55916 224828 258080 224856
rect 55916 224816 55922 224828
rect 258074 224816 258080 224828
rect 258132 224856 258138 224868
rect 258718 224856 258724 224868
rect 258132 224828 258724 224856
rect 258132 224816 258138 224828
rect 258718 224816 258724 224828
rect 258776 224816 258782 224868
rect 296714 224856 296720 224868
rect 277366 224828 296720 224856
rect 141510 224748 141516 224800
rect 141568 224788 141574 224800
rect 277366 224788 277394 224828
rect 296714 224816 296720 224828
rect 296772 224856 296778 224868
rect 297358 224856 297364 224868
rect 296772 224828 297364 224856
rect 296772 224816 296778 224828
rect 297358 224816 297364 224828
rect 297416 224816 297422 224868
rect 141568 224760 277394 224788
rect 141568 224748 141574 224760
rect 75914 224680 75920 224732
rect 75972 224720 75978 224732
rect 213914 224720 213920 224732
rect 75972 224692 213920 224720
rect 75972 224680 75978 224692
rect 213914 224680 213920 224692
rect 213972 224680 213978 224732
rect 213914 224408 213920 224460
rect 213972 224448 213978 224460
rect 214650 224448 214656 224460
rect 213972 224420 214656 224448
rect 213972 224408 213978 224420
rect 214650 224408 214656 224420
rect 214708 224408 214714 224460
rect 126422 224272 126428 224324
rect 126480 224312 126486 224324
rect 231118 224312 231124 224324
rect 126480 224284 231124 224312
rect 126480 224272 126486 224284
rect 231118 224272 231124 224284
rect 231176 224272 231182 224324
rect 100846 224204 100852 224256
rect 100904 224244 100910 224256
rect 255406 224244 255412 224256
rect 100904 224216 255412 224244
rect 100904 224204 100910 224216
rect 255406 224204 255412 224216
rect 255464 224204 255470 224256
rect 276658 224204 276664 224256
rect 276716 224244 276722 224256
rect 478874 224244 478880 224256
rect 276716 224216 478880 224244
rect 276716 224204 276722 224216
rect 478874 224204 478880 224216
rect 478932 224204 478938 224256
rect 82078 223524 82084 223576
rect 82136 223564 82142 223576
rect 313274 223564 313280 223576
rect 82136 223536 313280 223564
rect 82136 223524 82142 223536
rect 313274 223524 313280 223536
rect 313332 223564 313338 223576
rect 313918 223564 313924 223576
rect 313332 223536 313924 223564
rect 313332 223524 313338 223536
rect 313918 223524 313924 223536
rect 313976 223524 313982 223576
rect 70486 223456 70492 223508
rect 70544 223496 70550 223508
rect 201494 223496 201500 223508
rect 70544 223468 201500 223496
rect 70544 223456 70550 223468
rect 201494 223456 201500 223468
rect 201552 223496 201558 223508
rect 202414 223496 202420 223508
rect 201552 223468 202420 223496
rect 201552 223456 201558 223468
rect 202414 223456 202420 223468
rect 202472 223456 202478 223508
rect 148502 223388 148508 223440
rect 148560 223428 148566 223440
rect 238754 223428 238760 223440
rect 148560 223400 238760 223428
rect 148560 223388 148566 223400
rect 238754 223388 238760 223400
rect 238812 223428 238818 223440
rect 239398 223428 239404 223440
rect 238812 223400 239404 223428
rect 238812 223388 238818 223400
rect 239398 223388 239404 223400
rect 239456 223388 239462 223440
rect 177390 222980 177396 223032
rect 177448 223020 177454 223032
rect 232498 223020 232504 223032
rect 177448 222992 232504 223020
rect 177448 222980 177454 222992
rect 232498 222980 232504 222992
rect 232556 222980 232562 223032
rect 122098 222912 122104 222964
rect 122156 222952 122162 222964
rect 254026 222952 254032 222964
rect 122156 222924 254032 222952
rect 122156 222912 122162 222924
rect 254026 222912 254032 222924
rect 254084 222912 254090 222964
rect 301498 222912 301504 222964
rect 301556 222952 301562 222964
rect 495710 222952 495716 222964
rect 301556 222924 495716 222952
rect 301556 222912 301562 222924
rect 495710 222912 495716 222924
rect 495768 222912 495774 222964
rect 60458 222844 60464 222896
rect 60516 222884 60522 222896
rect 162210 222884 162216 222896
rect 60516 222856 162216 222884
rect 60516 222844 60522 222856
rect 162210 222844 162216 222856
rect 162268 222844 162274 222896
rect 195790 222844 195796 222896
rect 195848 222884 195854 222896
rect 471238 222884 471244 222896
rect 195848 222856 471244 222884
rect 195848 222844 195854 222856
rect 471238 222844 471244 222856
rect 471296 222844 471302 222896
rect 154022 222096 154028 222148
rect 154080 222136 154086 222148
rect 309134 222136 309140 222148
rect 154080 222108 309140 222136
rect 154080 222096 154086 222108
rect 309134 222096 309140 222108
rect 309192 222136 309198 222148
rect 309870 222136 309876 222148
rect 309192 222108 309876 222136
rect 309192 222096 309198 222108
rect 309870 222096 309876 222108
rect 309928 222096 309934 222148
rect 79226 222028 79232 222080
rect 79284 222068 79290 222080
rect 218698 222068 218704 222080
rect 79284 222040 218704 222068
rect 79284 222028 79290 222040
rect 218698 222028 218704 222040
rect 218756 222028 218762 222080
rect 73798 221960 73804 222012
rect 73856 222000 73862 222012
rect 182082 222000 182088 222012
rect 73856 221972 182088 222000
rect 73856 221960 73862 221972
rect 182082 221960 182088 221972
rect 182140 221960 182146 222012
rect 158070 221892 158076 221944
rect 158128 221932 158134 221944
rect 237374 221932 237380 221944
rect 158128 221904 237380 221932
rect 158128 221892 158134 221904
rect 237374 221892 237380 221904
rect 237432 221892 237438 221944
rect 92566 221552 92572 221604
rect 92624 221592 92630 221604
rect 228450 221592 228456 221604
rect 92624 221564 228456 221592
rect 92624 221552 92630 221564
rect 228450 221552 228456 221564
rect 228508 221552 228514 221604
rect 182082 221484 182088 221536
rect 182140 221524 182146 221536
rect 347866 221524 347872 221536
rect 182140 221496 347872 221524
rect 182140 221484 182146 221496
rect 347866 221484 347872 221496
rect 347924 221484 347930 221536
rect 192938 221416 192944 221468
rect 192996 221456 193002 221468
rect 510706 221456 510712 221468
rect 192996 221428 510712 221456
rect 192996 221416 193002 221428
rect 510706 221416 510712 221428
rect 510764 221416 510770 221468
rect 247034 220804 247040 220856
rect 247092 220844 247098 220856
rect 323670 220844 323676 220856
rect 247092 220816 323676 220844
rect 247092 220804 247098 220816
rect 323670 220804 323676 220816
rect 323728 220804 323734 220856
rect 156690 220736 156696 220788
rect 156748 220776 156754 220788
rect 314102 220776 314108 220788
rect 156748 220748 314108 220776
rect 156748 220736 156754 220748
rect 314102 220736 314108 220748
rect 314160 220736 314166 220788
rect 429838 220736 429844 220788
rect 429896 220776 429902 220788
rect 431218 220776 431224 220788
rect 429896 220748 431224 220776
rect 429896 220736 429902 220748
rect 431218 220736 431224 220748
rect 431276 220736 431282 220788
rect 93946 220668 93952 220720
rect 94004 220708 94010 220720
rect 247034 220708 247040 220720
rect 94004 220680 247040 220708
rect 94004 220668 94010 220680
rect 247034 220668 247040 220680
rect 247092 220668 247098 220720
rect 84378 220600 84384 220652
rect 84436 220640 84442 220652
rect 230474 220640 230480 220652
rect 84436 220612 230480 220640
rect 84436 220600 84442 220612
rect 230474 220600 230480 220612
rect 230532 220640 230538 220652
rect 231210 220640 231216 220652
rect 230532 220612 231216 220640
rect 230532 220600 230538 220612
rect 231210 220600 231216 220612
rect 231268 220600 231274 220652
rect 163682 220192 163688 220244
rect 163740 220232 163746 220244
rect 259454 220232 259460 220244
rect 163740 220204 259460 220232
rect 163740 220192 163746 220204
rect 259454 220192 259460 220204
rect 259512 220192 259518 220244
rect 167730 220124 167736 220176
rect 167788 220164 167794 220176
rect 289078 220164 289084 220176
rect 167788 220136 289084 220164
rect 167788 220124 167794 220136
rect 289078 220124 289084 220136
rect 289136 220124 289142 220176
rect 68922 220056 68928 220108
rect 68980 220096 68986 220108
rect 253934 220096 253940 220108
rect 68980 220068 253940 220096
rect 68980 220056 68986 220068
rect 253934 220056 253940 220068
rect 253992 220056 253998 220108
rect 293218 220056 293224 220108
rect 293276 220096 293282 220108
rect 429838 220096 429844 220108
rect 293276 220068 429844 220096
rect 293276 220056 293282 220068
rect 429838 220056 429844 220068
rect 429896 220056 429902 220108
rect 88978 219376 88984 219428
rect 89036 219416 89042 219428
rect 266354 219416 266360 219428
rect 89036 219388 266360 219416
rect 89036 219376 89042 219388
rect 266354 219376 266360 219388
rect 266412 219376 266418 219428
rect 84286 219308 84292 219360
rect 84344 219348 84350 219360
rect 228542 219348 228548 219360
rect 84344 219320 228548 219348
rect 84344 219308 84350 219320
rect 228542 219308 228548 219320
rect 228600 219308 228606 219360
rect 172422 218900 172428 218952
rect 172480 218940 172486 218952
rect 227070 218940 227076 218952
rect 172480 218912 227076 218940
rect 172480 218900 172486 218912
rect 227070 218900 227076 218912
rect 227128 218900 227134 218952
rect 134702 218832 134708 218884
rect 134760 218872 134766 218884
rect 236638 218872 236644 218884
rect 134760 218844 236644 218872
rect 134760 218832 134766 218844
rect 236638 218832 236644 218844
rect 236696 218832 236702 218884
rect 138750 218764 138756 218816
rect 138808 218804 138814 218816
rect 263594 218804 263600 218816
rect 138808 218776 263600 218804
rect 138808 218764 138814 218776
rect 263594 218764 263600 218776
rect 263652 218764 263658 218816
rect 147122 218696 147128 218748
rect 147180 218736 147186 218748
rect 278774 218736 278780 218748
rect 147180 218708 278780 218736
rect 147180 218696 147186 218708
rect 278774 218696 278780 218708
rect 278832 218696 278838 218748
rect 520918 218696 520924 218748
rect 520976 218736 520982 218748
rect 579798 218736 579804 218748
rect 520976 218708 579804 218736
rect 520976 218696 520982 218708
rect 579798 218696 579804 218708
rect 579856 218696 579862 218748
rect 266354 218016 266360 218068
rect 266412 218056 266418 218068
rect 266998 218056 267004 218068
rect 266412 218028 267004 218056
rect 266412 218016 266418 218028
rect 266998 218016 267004 218028
rect 267056 218016 267062 218068
rect 107746 217948 107752 218000
rect 107804 217988 107810 218000
rect 283558 217988 283564 218000
rect 107804 217960 283564 217988
rect 107804 217948 107810 217960
rect 283558 217948 283564 217960
rect 283616 217948 283622 218000
rect 131850 217540 131856 217592
rect 131908 217580 131914 217592
rect 238202 217580 238208 217592
rect 131908 217552 238208 217580
rect 131908 217540 131914 217552
rect 238202 217540 238208 217552
rect 238260 217540 238266 217592
rect 93854 217472 93860 217524
rect 93912 217512 93918 217524
rect 249886 217512 249892 217524
rect 93912 217484 249892 217512
rect 93912 217472 93918 217484
rect 249886 217472 249892 217484
rect 249944 217472 249950 217524
rect 77294 217404 77300 217456
rect 77352 217444 77358 217456
rect 249058 217444 249064 217456
rect 77352 217416 249064 217444
rect 77352 217404 77358 217416
rect 249058 217404 249064 217416
rect 249116 217404 249122 217456
rect 237374 217336 237380 217388
rect 237432 217376 237438 217388
rect 483014 217376 483020 217388
rect 237432 217348 483020 217376
rect 237432 217336 237438 217348
rect 483014 217336 483020 217348
rect 483072 217336 483078 217388
rect 177850 217268 177856 217320
rect 177908 217308 177914 217320
rect 436094 217308 436100 217320
rect 177908 217280 436100 217308
rect 177908 217268 177914 217280
rect 436094 217268 436100 217280
rect 436152 217268 436158 217320
rect 191742 216656 191748 216708
rect 191800 216696 191806 216708
rect 198182 216696 198188 216708
rect 191800 216668 198188 216696
rect 191800 216656 191806 216668
rect 198182 216656 198188 216668
rect 198240 216656 198246 216708
rect 114554 216588 114560 216640
rect 114612 216628 114618 216640
rect 295334 216628 295340 216640
rect 114612 216600 295340 216628
rect 114612 216588 114618 216600
rect 295334 216588 295340 216600
rect 295392 216588 295398 216640
rect 57606 216520 57612 216572
rect 57664 216560 57670 216572
rect 233234 216560 233240 216572
rect 57664 216532 233240 216560
rect 57664 216520 57670 216532
rect 233234 216520 233240 216532
rect 233292 216520 233298 216572
rect 198642 215976 198648 216028
rect 198700 216016 198706 216028
rect 325878 216016 325884 216028
rect 198700 215988 325884 216016
rect 198700 215976 198706 215988
rect 325878 215976 325884 215988
rect 325936 215976 325942 216028
rect 175090 215908 175096 215960
rect 175148 215948 175154 215960
rect 497458 215948 497464 215960
rect 175148 215920 497464 215948
rect 175148 215908 175154 215920
rect 497458 215908 497464 215920
rect 497516 215908 497522 215960
rect 295334 215296 295340 215348
rect 295392 215336 295398 215348
rect 295978 215336 295984 215348
rect 295392 215308 295984 215336
rect 295392 215296 295398 215308
rect 295978 215296 295984 215308
rect 296036 215296 296042 215348
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 14458 215268 14464 215280
rect 3384 215240 14464 215268
rect 3384 215228 3390 215240
rect 14458 215228 14464 215240
rect 14516 215228 14522 215280
rect 103698 215228 103704 215280
rect 103756 215268 103762 215280
rect 271874 215268 271880 215280
rect 103756 215240 271880 215268
rect 103756 215228 103762 215240
rect 271874 215228 271880 215240
rect 271932 215228 271938 215280
rect 83458 215160 83464 215212
rect 83516 215200 83522 215212
rect 208394 215200 208400 215212
rect 83516 215172 208400 215200
rect 83516 215160 83522 215172
rect 208394 215160 208400 215172
rect 208452 215160 208458 215212
rect 208394 214820 208400 214872
rect 208452 214860 208458 214872
rect 209038 214860 209044 214872
rect 208452 214832 209044 214860
rect 208452 214820 208458 214832
rect 209038 214820 209044 214832
rect 209096 214820 209102 214872
rect 166258 214752 166264 214804
rect 166316 214792 166322 214804
rect 240778 214792 240784 214804
rect 166316 214764 240784 214792
rect 166316 214752 166322 214764
rect 240778 214752 240784 214764
rect 240836 214752 240842 214804
rect 271874 214752 271880 214804
rect 271932 214792 271938 214804
rect 272518 214792 272524 214804
rect 271932 214764 272524 214792
rect 271932 214752 271938 214764
rect 272518 214752 272524 214764
rect 272576 214752 272582 214804
rect 184750 214684 184756 214736
rect 184808 214724 184814 214736
rect 389818 214724 389824 214736
rect 184808 214696 389824 214724
rect 184808 214684 184814 214696
rect 389818 214684 389824 214696
rect 389876 214684 389882 214736
rect 41230 214616 41236 214668
rect 41288 214656 41294 214668
rect 270494 214656 270500 214668
rect 41288 214628 270500 214656
rect 41288 214616 41294 214628
rect 270494 214616 270500 214628
rect 270552 214616 270558 214668
rect 157978 214548 157984 214600
rect 158036 214588 158042 214600
rect 216030 214588 216036 214600
rect 158036 214560 216036 214588
rect 158036 214548 158042 214560
rect 216030 214548 216036 214560
rect 216088 214548 216094 214600
rect 233234 214548 233240 214600
rect 233292 214588 233298 214600
rect 486418 214588 486424 214600
rect 233292 214560 486424 214588
rect 233292 214548 233298 214560
rect 486418 214548 486424 214560
rect 486476 214548 486482 214600
rect 102226 213868 102232 213920
rect 102284 213908 102290 213920
rect 273254 213908 273260 213920
rect 102284 213880 273260 213908
rect 102284 213868 102290 213880
rect 273254 213868 273260 213880
rect 273312 213908 273318 213920
rect 273898 213908 273904 213920
rect 273312 213880 273904 213908
rect 273312 213868 273318 213880
rect 273898 213868 273904 213880
rect 273956 213868 273962 213920
rect 176010 213392 176016 213444
rect 176068 213432 176074 213444
rect 291838 213432 291844 213444
rect 176068 213404 291844 213432
rect 176068 213392 176074 213404
rect 291838 213392 291844 213404
rect 291896 213392 291902 213444
rect 74534 213324 74540 213376
rect 74592 213364 74598 213376
rect 246298 213364 246304 213376
rect 74592 213336 246304 213364
rect 74592 213324 74598 213336
rect 246298 213324 246304 213336
rect 246356 213324 246362 213376
rect 56502 213256 56508 213308
rect 56560 213296 56566 213308
rect 258258 213296 258264 213308
rect 56560 213268 258264 213296
rect 56560 213256 56566 213268
rect 258258 213256 258264 213268
rect 258316 213256 258322 213308
rect 190270 213188 190276 213240
rect 190328 213228 190334 213240
rect 393958 213228 393964 213240
rect 190328 213200 393964 213228
rect 190328 213188 190334 213200
rect 393958 213188 393964 213200
rect 394016 213188 394022 213240
rect 184290 211896 184296 211948
rect 184348 211936 184354 211948
rect 256970 211936 256976 211948
rect 184348 211908 256976 211936
rect 184348 211896 184354 211908
rect 256970 211896 256976 211908
rect 257028 211896 257034 211948
rect 258718 211896 258724 211948
rect 258776 211936 258782 211948
rect 342898 211936 342904 211948
rect 258776 211908 342904 211936
rect 258776 211896 258782 211908
rect 342898 211896 342904 211908
rect 342956 211896 342962 211948
rect 106918 211828 106924 211880
rect 106976 211868 106982 211880
rect 274634 211868 274640 211880
rect 106976 211840 274640 211868
rect 106976 211828 106982 211840
rect 274634 211828 274640 211840
rect 274692 211828 274698 211880
rect 118694 211760 118700 211812
rect 118752 211800 118758 211812
rect 307754 211800 307760 211812
rect 118752 211772 307760 211800
rect 118752 211760 118758 211772
rect 307754 211760 307760 211772
rect 307812 211760 307818 211812
rect 432598 211080 432604 211132
rect 432656 211120 432662 211132
rect 446398 211120 446404 211132
rect 432656 211092 446404 211120
rect 432656 211080 432662 211092
rect 446398 211080 446404 211092
rect 446456 211080 446462 211132
rect 431954 210672 431960 210724
rect 432012 210712 432018 210724
rect 432598 210712 432604 210724
rect 432012 210684 432604 210712
rect 432012 210672 432018 210684
rect 432598 210672 432604 210684
rect 432656 210672 432662 210724
rect 115934 210536 115940 210588
rect 115992 210576 115998 210588
rect 245010 210576 245016 210588
rect 115992 210548 245016 210576
rect 115992 210536 115998 210548
rect 245010 210536 245016 210548
rect 245068 210536 245074 210588
rect 86218 210468 86224 210520
rect 86276 210508 86282 210520
rect 224954 210508 224960 210520
rect 86276 210480 224960 210508
rect 86276 210468 86282 210480
rect 224954 210468 224960 210480
rect 225012 210468 225018 210520
rect 304258 210468 304264 210520
rect 304316 210508 304322 210520
rect 498378 210508 498384 210520
rect 304316 210480 498384 210508
rect 304316 210468 304322 210480
rect 498378 210468 498384 210480
rect 498436 210468 498442 210520
rect 179230 210400 179236 210452
rect 179288 210440 179294 210452
rect 417418 210440 417424 210452
rect 179288 210412 417424 210440
rect 179288 210400 179294 210412
rect 417418 210400 417424 210412
rect 417476 210400 417482 210452
rect 447778 210400 447784 210452
rect 447836 210440 447842 210452
rect 480254 210440 480260 210452
rect 447836 210412 480260 210440
rect 447836 210400 447842 210412
rect 480254 210400 480260 210412
rect 480312 210400 480318 210452
rect 104894 209720 104900 209772
rect 104952 209760 104958 209772
rect 281534 209760 281540 209772
rect 104952 209732 281540 209760
rect 104952 209720 104958 209732
rect 281534 209720 281540 209732
rect 281592 209720 281598 209772
rect 113174 209652 113180 209704
rect 113232 209692 113238 209704
rect 179322 209692 179328 209704
rect 113232 209664 179328 209692
rect 113232 209652 113238 209664
rect 179322 209652 179328 209664
rect 179380 209652 179386 209704
rect 133230 209244 133236 209296
rect 133288 209284 133294 209296
rect 240870 209284 240876 209296
rect 133288 209256 240876 209284
rect 133288 209244 133294 209256
rect 240870 209244 240876 209256
rect 240928 209244 240934 209296
rect 179322 209176 179328 209228
rect 179380 209216 179386 209228
rect 338114 209216 338120 209228
rect 179380 209188 338120 209216
rect 179380 209176 179386 209188
rect 338114 209176 338120 209188
rect 338172 209176 338178 209228
rect 169662 209108 169668 209160
rect 169720 209148 169726 209160
rect 367738 209148 367744 209160
rect 169720 209120 367744 209148
rect 169720 209108 169726 209120
rect 367738 209108 367744 209120
rect 367796 209108 367802 209160
rect 11698 209040 11704 209092
rect 11756 209080 11762 209092
rect 111058 209080 111064 209092
rect 11756 209052 111064 209080
rect 11756 209040 11762 209052
rect 111058 209040 111064 209052
rect 111116 209040 111122 209092
rect 218790 209040 218796 209092
rect 218848 209080 218854 209092
rect 494238 209080 494244 209092
rect 218848 209052 494244 209080
rect 218848 209040 218854 209052
rect 494238 209040 494244 209052
rect 494296 209040 494302 209092
rect 281534 208360 281540 208412
rect 281592 208400 281598 208412
rect 282270 208400 282276 208412
rect 281592 208372 282276 208400
rect 281592 208360 281598 208372
rect 282270 208360 282276 208372
rect 282328 208360 282334 208412
rect 95234 208292 95240 208344
rect 95292 208332 95298 208344
rect 260834 208332 260840 208344
rect 95292 208304 260840 208332
rect 95292 208292 95298 208304
rect 260834 208292 260840 208304
rect 260892 208292 260898 208344
rect 197262 207952 197268 208004
rect 197320 207992 197326 208004
rect 238018 207992 238024 208004
rect 197320 207964 238024 207992
rect 197320 207952 197326 207964
rect 238018 207952 238024 207964
rect 238076 207952 238082 208004
rect 165522 207884 165528 207936
rect 165580 207924 165586 207936
rect 222838 207924 222844 207936
rect 165580 207896 222844 207924
rect 165580 207884 165586 207896
rect 222838 207884 222844 207896
rect 222896 207884 222902 207936
rect 214650 207816 214656 207868
rect 214708 207856 214714 207868
rect 329926 207856 329932 207868
rect 214708 207828 329932 207856
rect 214708 207816 214714 207828
rect 329926 207816 329932 207828
rect 329984 207816 329990 207868
rect 89714 207748 89720 207800
rect 89772 207788 89778 207800
rect 252738 207788 252744 207800
rect 89772 207760 252744 207788
rect 89772 207748 89778 207760
rect 252738 207748 252744 207760
rect 252796 207748 252802 207800
rect 135898 207680 135904 207732
rect 135956 207720 135962 207732
rect 360194 207720 360200 207732
rect 135956 207692 360200 207720
rect 135956 207680 135962 207692
rect 360194 207680 360200 207692
rect 360252 207680 360258 207732
rect 46750 207612 46756 207664
rect 46808 207652 46814 207664
rect 214558 207652 214564 207664
rect 46808 207624 214564 207652
rect 46808 207612 46814 207624
rect 214558 207612 214564 207624
rect 214616 207612 214622 207664
rect 239398 207612 239404 207664
rect 239456 207652 239462 207664
rect 514754 207652 514760 207664
rect 239456 207624 514760 207652
rect 239456 207612 239462 207624
rect 514754 207612 514760 207624
rect 514812 207612 514818 207664
rect 260834 207068 260840 207120
rect 260892 207108 260898 207120
rect 261478 207108 261484 207120
rect 260892 207080 261484 207108
rect 260892 207068 260898 207080
rect 261478 207068 261484 207080
rect 261536 207068 261542 207120
rect 346486 207040 346492 207052
rect 250824 207012 346492 207040
rect 92474 206932 92480 206984
rect 92532 206972 92538 206984
rect 249794 206972 249800 206984
rect 92532 206944 249800 206972
rect 92532 206932 92538 206944
rect 249794 206932 249800 206944
rect 249852 206972 249858 206984
rect 250824 206972 250852 207012
rect 346486 207000 346492 207012
rect 346544 207000 346550 207052
rect 249852 206944 250852 206972
rect 249852 206932 249858 206944
rect 100754 206388 100760 206440
rect 100812 206428 100818 206440
rect 255498 206428 255504 206440
rect 100812 206400 255504 206428
rect 100812 206388 100818 206400
rect 255498 206388 255504 206400
rect 255556 206388 255562 206440
rect 63310 206320 63316 206372
rect 63368 206360 63374 206372
rect 282178 206360 282184 206372
rect 63368 206332 282184 206360
rect 63368 206320 63374 206332
rect 282178 206320 282184 206332
rect 282236 206320 282242 206372
rect 180702 206252 180708 206304
rect 180760 206292 180766 206304
rect 505094 206292 505100 206304
rect 180760 206264 505100 206292
rect 180760 206252 180766 206264
rect 505094 206252 505100 206264
rect 505152 206252 505158 206304
rect 514754 206252 514760 206304
rect 514812 206292 514818 206304
rect 515398 206292 515404 206304
rect 514812 206264 515404 206292
rect 514812 206252 514818 206264
rect 515398 206252 515404 206264
rect 515456 206292 515462 206304
rect 580166 206292 580172 206304
rect 515456 206264 580172 206292
rect 515456 206252 515462 206264
rect 580166 206252 580172 206264
rect 580224 206252 580230 206304
rect 107654 205572 107660 205624
rect 107712 205612 107718 205624
rect 285674 205612 285680 205624
rect 107712 205584 285680 205612
rect 107712 205572 107718 205584
rect 285674 205572 285680 205584
rect 285732 205572 285738 205624
rect 285674 205096 285680 205148
rect 285732 205136 285738 205148
rect 286410 205136 286416 205148
rect 285732 205108 286416 205136
rect 285732 205096 285738 205108
rect 286410 205096 286416 205108
rect 286468 205096 286474 205148
rect 222930 204960 222936 205012
rect 222988 205000 222994 205012
rect 320910 205000 320916 205012
rect 222988 204972 320916 205000
rect 222988 204960 222994 204972
rect 320910 204960 320916 204972
rect 320968 204960 320974 205012
rect 65886 204892 65892 204944
rect 65944 204932 65950 204944
rect 240962 204932 240968 204944
rect 65944 204904 240968 204932
rect 65944 204892 65950 204904
rect 240962 204892 240968 204904
rect 241020 204892 241026 204944
rect 262950 204892 262956 204944
rect 263008 204932 263014 204944
rect 494146 204932 494152 204944
rect 263008 204904 494152 204932
rect 263008 204892 263014 204904
rect 494146 204892 494152 204904
rect 494204 204892 494210 204944
rect 97994 204212 98000 204264
rect 98052 204252 98058 204264
rect 146938 204252 146944 204264
rect 98052 204224 146944 204252
rect 98052 204212 98058 204224
rect 146938 204212 146944 204224
rect 146996 204212 147002 204264
rect 156598 203736 156604 203788
rect 156656 203776 156662 203788
rect 266354 203776 266360 203788
rect 156656 203748 266360 203776
rect 156656 203736 156662 203748
rect 266354 203736 266360 203748
rect 266412 203736 266418 203788
rect 149698 203668 149704 203720
rect 149756 203708 149762 203720
rect 280798 203708 280804 203720
rect 149756 203680 280804 203708
rect 149756 203668 149762 203680
rect 280798 203668 280804 203680
rect 280856 203668 280862 203720
rect 99374 203600 99380 203652
rect 99432 203640 99438 203652
rect 254118 203640 254124 203652
rect 99432 203612 254124 203640
rect 99432 203600 99438 203612
rect 254118 203600 254124 203612
rect 254176 203600 254182 203652
rect 146938 203532 146944 203584
rect 146996 203572 147002 203584
rect 392578 203572 392584 203584
rect 146996 203544 392584 203572
rect 146996 203532 147002 203544
rect 392578 203532 392584 203544
rect 392636 203532 392642 203584
rect 217318 202376 217324 202428
rect 217376 202416 217382 202428
rect 321554 202416 321560 202428
rect 217376 202388 321560 202416
rect 217376 202376 217382 202388
rect 321554 202376 321560 202388
rect 321612 202376 321618 202428
rect 123754 202308 123760 202360
rect 123812 202348 123818 202360
rect 262214 202348 262220 202360
rect 123812 202320 262220 202348
rect 123812 202308 123818 202320
rect 262214 202308 262220 202320
rect 262272 202308 262278 202360
rect 45462 202240 45468 202292
rect 45520 202280 45526 202292
rect 232590 202280 232596 202292
rect 45520 202252 232596 202280
rect 45520 202240 45526 202252
rect 232590 202240 232596 202252
rect 232648 202240 232654 202292
rect 69106 202172 69112 202224
rect 69164 202212 69170 202224
rect 280154 202212 280160 202224
rect 69164 202184 280160 202212
rect 69164 202172 69170 202184
rect 280154 202172 280160 202184
rect 280212 202172 280218 202224
rect 322198 202172 322204 202224
rect 322256 202212 322262 202224
rect 328638 202212 328644 202224
rect 322256 202184 328644 202212
rect 322256 202172 322262 202184
rect 328638 202172 328644 202184
rect 328696 202172 328702 202224
rect 159542 202104 159548 202156
rect 159600 202144 159606 202156
rect 381538 202144 381544 202156
rect 159600 202116 381544 202144
rect 159600 202104 159606 202116
rect 381538 202104 381544 202116
rect 381596 202104 381602 202156
rect 126330 200880 126336 200932
rect 126388 200920 126394 200932
rect 242250 200920 242256 200932
rect 126388 200892 242256 200920
rect 126388 200880 126394 200892
rect 242250 200880 242256 200892
rect 242308 200880 242314 200932
rect 269758 200880 269764 200932
rect 269816 200920 269822 200932
rect 327258 200920 327264 200932
rect 269816 200892 327264 200920
rect 269816 200880 269822 200892
rect 327258 200880 327264 200892
rect 327316 200880 327322 200932
rect 86954 200812 86960 200864
rect 87012 200852 87018 200864
rect 274726 200852 274732 200864
rect 87012 200824 274732 200852
rect 87012 200812 87018 200824
rect 274726 200812 274732 200824
rect 274784 200812 274790 200864
rect 144178 200744 144184 200796
rect 144236 200784 144242 200796
rect 509326 200784 509332 200796
rect 144236 200756 509332 200784
rect 144236 200744 144242 200756
rect 509326 200744 509332 200756
rect 509384 200744 509390 200796
rect 145650 199588 145656 199640
rect 145708 199628 145714 199640
rect 276658 199628 276664 199640
rect 145708 199600 276664 199628
rect 145708 199588 145714 199600
rect 276658 199588 276664 199600
rect 276716 199588 276722 199640
rect 104158 199520 104164 199572
rect 104216 199560 104222 199572
rect 260926 199560 260932 199572
rect 104216 199532 260932 199560
rect 104216 199520 104222 199532
rect 260926 199520 260932 199532
rect 260984 199520 260990 199572
rect 53650 199452 53656 199504
rect 53708 199492 53714 199504
rect 238110 199492 238116 199504
rect 53708 199464 238116 199492
rect 53708 199452 53714 199464
rect 238110 199452 238116 199464
rect 238168 199452 238174 199504
rect 261478 199452 261484 199504
rect 261536 199492 261542 199504
rect 321830 199492 321836 199504
rect 261536 199464 321836 199492
rect 261536 199452 261542 199464
rect 321830 199452 321836 199464
rect 321888 199452 321894 199504
rect 211798 199384 211804 199436
rect 211856 199424 211862 199436
rect 514754 199424 514760 199436
rect 211856 199396 514760 199424
rect 211856 199384 211862 199396
rect 514754 199384 514760 199396
rect 514812 199384 514818 199436
rect 181530 198228 181536 198280
rect 181588 198268 181594 198280
rect 213178 198268 213184 198280
rect 181588 198240 213184 198268
rect 181588 198228 181594 198240
rect 213178 198228 213184 198240
rect 213236 198228 213242 198280
rect 162210 198160 162216 198212
rect 162268 198200 162274 198212
rect 262306 198200 262312 198212
rect 162268 198172 262312 198200
rect 162268 198160 162274 198172
rect 262306 198160 262312 198172
rect 262364 198160 262370 198212
rect 102134 198092 102140 198144
rect 102192 198132 102198 198144
rect 250070 198132 250076 198144
rect 102192 198104 250076 198132
rect 102192 198092 102198 198104
rect 250070 198092 250076 198104
rect 250128 198092 250134 198144
rect 67450 198024 67456 198076
rect 67508 198064 67514 198076
rect 251174 198064 251180 198076
rect 67508 198036 251180 198064
rect 67508 198024 67514 198036
rect 251174 198024 251180 198036
rect 251232 198024 251238 198076
rect 127618 197956 127624 198008
rect 127676 197996 127682 198008
rect 195330 197996 195336 198008
rect 127676 197968 195336 197996
rect 127676 197956 127682 197968
rect 195330 197956 195336 197968
rect 195388 197956 195394 198008
rect 213270 197956 213276 198008
rect 213328 197996 213334 198008
rect 451274 197996 451280 198008
rect 213328 197968 451280 197996
rect 213328 197956 213334 197968
rect 451274 197956 451280 197968
rect 451332 197956 451338 198008
rect 238202 196800 238208 196852
rect 238260 196840 238266 196852
rect 271966 196840 271972 196852
rect 238260 196812 271972 196840
rect 238260 196800 238266 196812
rect 271966 196800 271972 196812
rect 272024 196800 272030 196852
rect 126238 196732 126244 196784
rect 126296 196772 126302 196784
rect 184290 196772 184296 196784
rect 126296 196744 184296 196772
rect 126296 196732 126302 196744
rect 184290 196732 184296 196744
rect 184348 196732 184354 196784
rect 242158 196732 242164 196784
rect 242216 196772 242222 196784
rect 328730 196772 328736 196784
rect 242216 196744 328736 196772
rect 242216 196732 242222 196744
rect 328730 196732 328736 196744
rect 328788 196732 328794 196784
rect 142890 196664 142896 196716
rect 142948 196704 142954 196716
rect 243538 196704 243544 196716
rect 142948 196676 243544 196704
rect 142948 196664 142954 196676
rect 243538 196664 243544 196676
rect 243596 196664 243602 196716
rect 160922 196596 160928 196648
rect 160980 196636 160986 196648
rect 502334 196636 502340 196648
rect 160980 196608 502340 196636
rect 160980 196596 160986 196608
rect 502334 196596 502340 196608
rect 502392 196596 502398 196648
rect 129090 195508 129096 195560
rect 129148 195548 129154 195560
rect 213270 195548 213276 195560
rect 129148 195520 213276 195548
rect 129148 195508 129154 195520
rect 213270 195508 213276 195520
rect 213328 195508 213334 195560
rect 194502 195440 194508 195492
rect 194560 195480 194566 195492
rect 336918 195480 336924 195492
rect 194560 195452 336924 195480
rect 194560 195440 194566 195452
rect 336918 195440 336924 195452
rect 336976 195440 336982 195492
rect 70394 195372 70400 195424
rect 70452 195412 70458 195424
rect 254210 195412 254216 195424
rect 70452 195384 254216 195412
rect 70452 195372 70458 195384
rect 254210 195372 254216 195384
rect 254268 195372 254274 195424
rect 138658 195304 138664 195356
rect 138716 195344 138722 195356
rect 352006 195344 352012 195356
rect 138716 195316 352012 195344
rect 138716 195304 138722 195316
rect 352006 195304 352012 195316
rect 352064 195304 352070 195356
rect 78674 195236 78680 195288
rect 78732 195276 78738 195288
rect 267734 195276 267740 195288
rect 78732 195248 267740 195276
rect 78732 195236 78738 195248
rect 267734 195236 267740 195248
rect 267792 195236 267798 195288
rect 290458 195236 290464 195288
rect 290516 195276 290522 195288
rect 507946 195276 507952 195288
rect 290516 195248 507952 195276
rect 290516 195236 290522 195248
rect 507946 195236 507952 195248
rect 508004 195236 508010 195288
rect 151078 193944 151084 193996
rect 151136 193984 151142 193996
rect 286318 193984 286324 193996
rect 151136 193956 286324 193984
rect 151136 193944 151142 193956
rect 286318 193944 286324 193956
rect 286376 193944 286382 193996
rect 323578 193944 323584 193996
rect 323636 193984 323642 193996
rect 341058 193984 341064 193996
rect 323636 193956 341064 193984
rect 323636 193944 323642 193956
rect 341058 193944 341064 193956
rect 341116 193944 341122 193996
rect 111794 193876 111800 193928
rect 111852 193916 111858 193928
rect 252646 193916 252652 193928
rect 111852 193888 252652 193916
rect 111852 193876 111858 193888
rect 252646 193876 252652 193888
rect 252704 193876 252710 193928
rect 286410 193876 286416 193928
rect 286468 193916 286474 193928
rect 330110 193916 330116 193928
rect 286468 193888 330116 193916
rect 286468 193876 286474 193888
rect 330110 193876 330116 193888
rect 330168 193876 330174 193928
rect 128998 193808 129004 193860
rect 129056 193848 129062 193860
rect 369854 193848 369860 193860
rect 129056 193820 369860 193848
rect 129056 193808 129062 193820
rect 369854 193808 369860 193820
rect 369912 193808 369918 193860
rect 188430 192720 188436 192772
rect 188488 192760 188494 192772
rect 245102 192760 245108 192772
rect 188488 192732 245108 192760
rect 188488 192720 188494 192732
rect 245102 192720 245108 192732
rect 245160 192720 245166 192772
rect 224862 192652 224868 192704
rect 224920 192692 224926 192704
rect 318058 192692 318064 192704
rect 224920 192664 318064 192692
rect 224920 192652 224926 192664
rect 318058 192652 318064 192664
rect 318116 192652 318122 192704
rect 130378 192584 130384 192636
rect 130436 192624 130442 192636
rect 264974 192624 264980 192636
rect 130436 192596 264980 192624
rect 130436 192584 130442 192596
rect 264974 192584 264980 192596
rect 265032 192584 265038 192636
rect 272518 192584 272524 192636
rect 272576 192624 272582 192636
rect 325786 192624 325792 192636
rect 272576 192596 325792 192624
rect 272576 192584 272582 192596
rect 325786 192584 325792 192596
rect 325844 192584 325850 192636
rect 176102 192516 176108 192568
rect 176160 192556 176166 192568
rect 343818 192556 343824 192568
rect 176160 192528 343824 192556
rect 176160 192516 176166 192528
rect 343818 192516 343824 192528
rect 343876 192516 343882 192568
rect 137370 192448 137376 192500
rect 137428 192488 137434 192500
rect 357526 192488 357532 192500
rect 137428 192460 357532 192488
rect 137428 192448 137434 192460
rect 357526 192448 357532 192460
rect 357584 192448 357590 192500
rect 360838 192448 360844 192500
rect 360896 192488 360902 192500
rect 517514 192488 517520 192500
rect 360896 192460 517520 192488
rect 360896 192448 360902 192460
rect 517514 192448 517520 192460
rect 517572 192448 517578 192500
rect 134518 191156 134524 191208
rect 134576 191196 134582 191208
rect 269114 191196 269120 191208
rect 134576 191168 269120 191196
rect 134576 191156 134582 191168
rect 269114 191156 269120 191168
rect 269172 191156 269178 191208
rect 72418 191088 72424 191140
rect 72476 191128 72482 191140
rect 273438 191128 273444 191140
rect 72476 191100 273444 191128
rect 72476 191088 72482 191100
rect 273438 191088 273444 191100
rect 273496 191088 273502 191140
rect 133138 190068 133144 190120
rect 133196 190108 133202 190120
rect 200758 190108 200764 190120
rect 133196 190080 200764 190108
rect 133196 190068 133202 190080
rect 200758 190068 200764 190080
rect 200816 190068 200822 190120
rect 228542 190068 228548 190120
rect 228600 190108 228606 190120
rect 309778 190108 309784 190120
rect 228600 190080 309784 190108
rect 228600 190068 228606 190080
rect 309778 190068 309784 190080
rect 309836 190068 309842 190120
rect 164970 190000 164976 190052
rect 165028 190040 165034 190052
rect 258166 190040 258172 190052
rect 165028 190012 258172 190040
rect 165028 190000 165034 190012
rect 258166 190000 258172 190012
rect 258224 190000 258230 190052
rect 193122 189932 193128 189984
rect 193180 189972 193186 189984
rect 335630 189972 335636 189984
rect 193180 189944 335636 189972
rect 193180 189932 193186 189944
rect 335630 189932 335636 189944
rect 335688 189932 335694 189984
rect 76558 189864 76564 189916
rect 76616 189904 76622 189916
rect 260834 189904 260840 189916
rect 76616 189876 260840 189904
rect 76616 189864 76622 189876
rect 260834 189864 260840 189876
rect 260892 189864 260898 189916
rect 52270 189796 52276 189848
rect 52328 189836 52334 189848
rect 267826 189836 267832 189848
rect 52328 189808 267832 189836
rect 52328 189796 52334 189808
rect 267826 189796 267832 189808
rect 267884 189796 267890 189848
rect 297358 189796 297364 189848
rect 297416 189836 297422 189848
rect 501138 189836 501144 189848
rect 297416 189808 501144 189836
rect 297416 189796 297422 189808
rect 501138 189796 501144 189808
rect 501196 189796 501202 189848
rect 183462 189728 183468 189780
rect 183520 189768 183526 189780
rect 460106 189768 460112 189780
rect 183520 189740 460112 189768
rect 183520 189728 183526 189740
rect 460106 189728 460112 189740
rect 460164 189728 460170 189780
rect 268378 189048 268384 189100
rect 268436 189088 268442 189100
rect 269206 189088 269212 189100
rect 268436 189060 269212 189088
rect 268436 189048 268442 189060
rect 269206 189048 269212 189060
rect 269264 189048 269270 189100
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 53098 189020 53104 189032
rect 3476 188992 53104 189020
rect 3476 188980 3482 188992
rect 53098 188980 53104 188992
rect 53156 188980 53162 189032
rect 151170 188504 151176 188556
rect 151228 188544 151234 188556
rect 270678 188544 270684 188556
rect 151228 188516 270684 188544
rect 151228 188504 151234 188516
rect 270678 188504 270684 188516
rect 270736 188504 270742 188556
rect 142798 188436 142804 188488
rect 142856 188476 142862 188488
rect 196618 188476 196624 188488
rect 142856 188448 196624 188476
rect 142856 188436 142862 188448
rect 196618 188436 196624 188448
rect 196676 188436 196682 188488
rect 218698 188436 218704 188488
rect 218756 188476 218762 188488
rect 339586 188476 339592 188488
rect 218756 188448 339592 188476
rect 218756 188436 218762 188448
rect 339586 188436 339592 188448
rect 339644 188436 339650 188488
rect 84194 188368 84200 188420
rect 84252 188408 84258 188420
rect 249978 188408 249984 188420
rect 84252 188380 249984 188408
rect 84252 188368 84258 188380
rect 249978 188368 249984 188380
rect 250036 188368 250042 188420
rect 320818 188368 320824 188420
rect 320876 188408 320882 188420
rect 334066 188408 334072 188420
rect 320876 188380 334072 188408
rect 320876 188368 320882 188380
rect 334066 188368 334072 188380
rect 334124 188368 334130 188420
rect 47946 188300 47952 188352
rect 48004 188340 48010 188352
rect 256786 188340 256792 188352
rect 48004 188312 256792 188340
rect 48004 188300 48010 188312
rect 256786 188300 256792 188312
rect 256844 188300 256850 188352
rect 265618 188300 265624 188352
rect 265676 188340 265682 188352
rect 494330 188340 494336 188352
rect 265676 188312 494336 188340
rect 265676 188300 265682 188312
rect 494330 188300 494336 188312
rect 494388 188300 494394 188352
rect 235258 187280 235264 187332
rect 235316 187320 235322 187332
rect 308398 187320 308404 187332
rect 235316 187292 308404 187320
rect 235316 187280 235322 187292
rect 308398 187280 308404 187292
rect 308456 187280 308462 187332
rect 173250 187212 173256 187264
rect 173308 187252 173314 187264
rect 261018 187252 261024 187264
rect 173308 187224 261024 187252
rect 173308 187212 173314 187224
rect 261018 187212 261024 187224
rect 261076 187212 261082 187264
rect 147030 187144 147036 187196
rect 147088 187184 147094 187196
rect 189810 187184 189816 187196
rect 147088 187156 189816 187184
rect 147088 187144 147094 187156
rect 189810 187144 189816 187156
rect 189868 187144 189874 187196
rect 231210 187144 231216 187196
rect 231268 187184 231274 187196
rect 335538 187184 335544 187196
rect 231268 187156 335544 187184
rect 231268 187144 231274 187156
rect 335538 187144 335544 187156
rect 335596 187144 335602 187196
rect 110414 187076 110420 187128
rect 110472 187116 110478 187128
rect 249794 187116 249800 187128
rect 110472 187088 249800 187116
rect 110472 187076 110478 187088
rect 249794 187076 249800 187088
rect 249852 187076 249858 187128
rect 124858 187008 124864 187060
rect 124916 187048 124922 187060
rect 270586 187048 270592 187060
rect 124916 187020 270592 187048
rect 124916 187008 124922 187020
rect 270586 187008 270592 187020
rect 270644 187008 270650 187060
rect 173342 186940 173348 186992
rect 173400 186980 173406 186992
rect 342346 186980 342352 186992
rect 173400 186952 342352 186980
rect 173400 186940 173406 186952
rect 342346 186940 342352 186952
rect 342404 186940 342410 186992
rect 358078 186940 358084 186992
rect 358136 186980 358142 186992
rect 513374 186980 513380 186992
rect 358136 186952 513380 186980
rect 358136 186940 358142 186952
rect 513374 186940 513380 186952
rect 513432 186940 513438 186992
rect 148318 185784 148324 185836
rect 148376 185824 148382 185836
rect 210418 185824 210424 185836
rect 148376 185796 210424 185824
rect 148376 185784 148382 185796
rect 210418 185784 210424 185796
rect 210476 185784 210482 185836
rect 213362 185784 213368 185836
rect 213420 185824 213426 185836
rect 259546 185824 259552 185836
rect 213420 185796 259552 185824
rect 213420 185784 213426 185796
rect 259546 185784 259552 185796
rect 259604 185784 259610 185836
rect 177942 185716 177948 185768
rect 178000 185756 178006 185768
rect 345198 185756 345204 185768
rect 178000 185728 345204 185756
rect 178000 185716 178006 185728
rect 345198 185716 345204 185728
rect 345256 185716 345262 185768
rect 141418 185648 141424 185700
rect 141476 185688 141482 185700
rect 351178 185688 351184 185700
rect 141476 185660 351184 185688
rect 141476 185648 141482 185660
rect 351178 185648 351184 185660
rect 351236 185648 351242 185700
rect 422938 185648 422944 185700
rect 422996 185688 423002 185700
rect 450538 185688 450544 185700
rect 422996 185660 450544 185688
rect 422996 185648 423002 185660
rect 450538 185648 450544 185660
rect 450596 185648 450602 185700
rect 119338 185580 119344 185632
rect 119396 185620 119402 185632
rect 273346 185620 273352 185632
rect 119396 185592 273352 185620
rect 119396 185580 119402 185592
rect 273346 185580 273352 185592
rect 273404 185580 273410 185632
rect 278038 185580 278044 185632
rect 278096 185620 278102 185632
rect 503898 185620 503904 185632
rect 278096 185592 503904 185620
rect 278096 185580 278102 185592
rect 503898 185580 503904 185592
rect 503956 185580 503962 185632
rect 318610 185512 318616 185564
rect 318668 185552 318674 185564
rect 320174 185552 320180 185564
rect 318668 185524 320180 185552
rect 318668 185512 318674 185524
rect 320174 185512 320180 185524
rect 320232 185512 320238 185564
rect 102042 184968 102048 185020
rect 102100 185008 102106 185020
rect 169018 185008 169024 185020
rect 102100 184980 169024 185008
rect 102100 184968 102106 184980
rect 169018 184968 169024 184980
rect 169076 184968 169082 185020
rect 100662 184900 100668 184952
rect 100720 184940 100726 184952
rect 173158 184940 173164 184952
rect 100720 184912 173164 184940
rect 100720 184900 100726 184912
rect 173158 184900 173164 184912
rect 173216 184900 173222 184952
rect 232590 184424 232596 184476
rect 232648 184464 232654 184476
rect 266538 184464 266544 184476
rect 232648 184436 266544 184464
rect 232648 184424 232654 184436
rect 266538 184424 266544 184436
rect 266596 184424 266602 184476
rect 145558 184356 145564 184408
rect 145616 184396 145622 184408
rect 273254 184396 273260 184408
rect 145616 184368 273260 184396
rect 145616 184356 145622 184368
rect 273254 184356 273260 184368
rect 273312 184356 273318 184408
rect 140130 184288 140136 184340
rect 140188 184328 140194 184340
rect 278038 184328 278044 184340
rect 140188 184300 278044 184328
rect 140188 184288 140194 184300
rect 278038 184288 278044 184300
rect 278096 184288 278102 184340
rect 345658 184288 345664 184340
rect 345716 184328 345722 184340
rect 443914 184328 443920 184340
rect 345716 184300 443920 184328
rect 345716 184288 345722 184300
rect 443914 184288 443920 184300
rect 443972 184288 443978 184340
rect 468478 184288 468484 184340
rect 468536 184328 468542 184340
rect 510798 184328 510804 184340
rect 468536 184300 510804 184328
rect 468536 184288 468542 184300
rect 510798 184288 510804 184300
rect 510856 184288 510862 184340
rect 171778 184220 171784 184272
rect 171836 184260 171842 184272
rect 345290 184260 345296 184272
rect 171836 184232 345296 184260
rect 171836 184220 171842 184232
rect 345290 184220 345296 184232
rect 345348 184220 345354 184272
rect 400858 184220 400864 184272
rect 400916 184260 400922 184272
rect 505186 184260 505192 184272
rect 400916 184232 505192 184260
rect 400916 184220 400922 184232
rect 505186 184220 505192 184232
rect 505244 184220 505250 184272
rect 155218 184152 155224 184204
rect 155276 184192 155282 184204
rect 202138 184192 202144 184204
rect 155276 184164 202144 184192
rect 155276 184152 155282 184164
rect 202138 184152 202144 184164
rect 202196 184152 202202 184204
rect 227070 184152 227076 184204
rect 227128 184192 227134 184204
rect 507854 184192 507860 184204
rect 227128 184164 507860 184192
rect 227128 184152 227134 184164
rect 507854 184152 507860 184164
rect 507912 184152 507918 184204
rect 128262 183608 128268 183660
rect 128320 183648 128326 183660
rect 180242 183648 180248 183660
rect 128320 183620 180248 183648
rect 128320 183608 128326 183620
rect 180242 183608 180248 183620
rect 180300 183608 180306 183660
rect 107562 183540 107568 183592
rect 107620 183580 107626 183592
rect 196710 183580 196716 183592
rect 107620 183552 196716 183580
rect 107620 183540 107626 183552
rect 196710 183540 196716 183552
rect 196768 183540 196774 183592
rect 403618 183472 403624 183524
rect 403676 183512 403682 183524
rect 404262 183512 404268 183524
rect 403676 183484 404268 183512
rect 403676 183472 403682 183484
rect 404262 183472 404268 183484
rect 404320 183472 404326 183524
rect 236638 183132 236644 183184
rect 236696 183172 236702 183184
rect 263778 183172 263784 183184
rect 236696 183144 263784 183172
rect 236696 183132 236702 183144
rect 263778 183132 263784 183144
rect 263836 183132 263842 183184
rect 228358 183064 228364 183116
rect 228416 183104 228422 183116
rect 265066 183104 265072 183116
rect 228416 183076 265072 183104
rect 228416 183064 228422 183076
rect 265066 183064 265072 183076
rect 265124 183064 265130 183116
rect 251910 182996 251916 183048
rect 251968 183036 251974 183048
rect 345014 183036 345020 183048
rect 251968 183008 345020 183036
rect 251968 182996 251974 183008
rect 345014 182996 345020 183008
rect 345072 182996 345078 183048
rect 195238 182928 195244 182980
rect 195296 182968 195302 182980
rect 313826 182968 313832 182980
rect 195296 182940 313832 182968
rect 195296 182928 195302 182940
rect 313826 182928 313832 182940
rect 313884 182928 313890 182980
rect 200850 182860 200856 182912
rect 200908 182900 200914 182912
rect 338298 182900 338304 182912
rect 200908 182872 338304 182900
rect 200908 182860 200914 182872
rect 338298 182860 338304 182872
rect 338356 182860 338362 182912
rect 57698 182792 57704 182844
rect 57756 182832 57762 182844
rect 262398 182832 262404 182844
rect 57756 182804 262404 182832
rect 57756 182792 57762 182804
rect 262398 182792 262404 182804
rect 262456 182792 262462 182844
rect 314010 182792 314016 182844
rect 314068 182832 314074 182844
rect 331490 182832 331496 182844
rect 314068 182804 331496 182832
rect 314068 182792 314074 182804
rect 331490 182792 331496 182804
rect 331548 182792 331554 182844
rect 419350 182792 419356 182844
rect 419408 182832 419414 182844
rect 580350 182832 580356 182844
rect 419408 182804 580356 182832
rect 419408 182792 419414 182804
rect 580350 182792 580356 182804
rect 580408 182792 580414 182844
rect 132402 182452 132408 182504
rect 132460 182492 132466 182504
rect 164970 182492 164976 182504
rect 132460 182464 164976 182492
rect 132460 182452 132466 182464
rect 164970 182452 164976 182464
rect 165028 182452 165034 182504
rect 105722 182384 105728 182436
rect 105780 182424 105786 182436
rect 170766 182424 170772 182436
rect 105780 182396 170772 182424
rect 105780 182384 105786 182396
rect 170766 182384 170772 182396
rect 170824 182384 170830 182436
rect 119706 182316 119712 182368
rect 119764 182356 119770 182368
rect 204990 182356 204996 182368
rect 119764 182328 204996 182356
rect 119764 182316 119770 182328
rect 204990 182316 204996 182328
rect 205048 182316 205054 182368
rect 489178 182316 489184 182368
rect 489236 182356 489242 182368
rect 490558 182356 490564 182368
rect 489236 182328 490564 182356
rect 489236 182316 489242 182328
rect 490558 182316 490564 182328
rect 490616 182316 490622 182368
rect 110690 182248 110696 182300
rect 110748 182288 110754 182300
rect 196802 182288 196808 182300
rect 110748 182260 196808 182288
rect 110748 182248 110754 182260
rect 196802 182248 196808 182260
rect 196860 182248 196866 182300
rect 400858 182248 400864 182300
rect 400916 182288 400922 182300
rect 494054 182288 494060 182300
rect 400916 182260 494060 182288
rect 400916 182248 400922 182260
rect 494054 182248 494060 182260
rect 494112 182248 494118 182300
rect 123294 182180 123300 182232
rect 123352 182220 123358 182232
rect 214650 182220 214656 182232
rect 123352 182192 214656 182220
rect 123352 182180 123358 182192
rect 214650 182180 214656 182192
rect 214708 182180 214714 182232
rect 404262 182180 404268 182232
rect 404320 182220 404326 182232
rect 580258 182220 580264 182232
rect 404320 182192 580264 182220
rect 404320 182180 404326 182192
rect 580258 182180 580264 182192
rect 580316 182180 580322 182232
rect 454678 182112 454684 182164
rect 454736 182152 454742 182164
rect 455598 182152 455604 182164
rect 454736 182124 455604 182152
rect 454736 182112 454742 182124
rect 455598 182112 455604 182124
rect 455656 182112 455662 182164
rect 461578 182112 461584 182164
rect 461636 182152 461642 182164
rect 462590 182152 462596 182164
rect 461636 182124 462596 182152
rect 461636 182112 461642 182124
rect 462590 182112 462596 182124
rect 462648 182112 462654 182164
rect 471238 182112 471244 182164
rect 471296 182152 471302 182164
rect 476574 182152 476580 182164
rect 471296 182124 476580 182152
rect 471296 182112 471302 182124
rect 476574 182112 476580 182124
rect 476632 182112 476638 182164
rect 485038 182112 485044 182164
rect 485096 182152 485102 182164
rect 485774 182152 485780 182164
rect 485096 182124 485780 182152
rect 485096 182112 485102 182124
rect 485774 182112 485780 182124
rect 485832 182112 485838 182164
rect 245010 181772 245016 181824
rect 245068 181812 245074 181824
rect 263686 181812 263692 181824
rect 245068 181784 263692 181812
rect 245068 181772 245074 181784
rect 263686 181772 263692 181784
rect 263744 181772 263750 181824
rect 486418 181772 486424 181824
rect 486476 181812 486482 181824
rect 492858 181812 492864 181824
rect 486476 181784 492864 181812
rect 486476 181772 486482 181784
rect 492858 181772 492864 181784
rect 492916 181772 492922 181824
rect 168282 181704 168288 181756
rect 168340 181744 168346 181756
rect 216122 181744 216128 181756
rect 168340 181716 216128 181744
rect 168340 181704 168346 181716
rect 216122 181704 216128 181716
rect 216180 181704 216186 181756
rect 228450 181704 228456 181756
rect 228508 181744 228514 181756
rect 259730 181744 259736 181756
rect 228508 181716 259736 181744
rect 228508 181704 228514 181716
rect 259730 181704 259736 181716
rect 259788 181704 259794 181756
rect 307018 181704 307024 181756
rect 307076 181744 307082 181756
rect 336734 181744 336740 181756
rect 307076 181716 336740 181744
rect 307076 181704 307082 181716
rect 336734 181704 336740 181716
rect 336792 181704 336798 181756
rect 475378 181704 475384 181756
rect 475436 181744 475442 181756
rect 488626 181744 488632 181756
rect 475436 181716 488632 181744
rect 475436 181704 475442 181716
rect 488626 181704 488632 181716
rect 488684 181704 488690 181756
rect 170674 181636 170680 181688
rect 170732 181676 170738 181688
rect 251266 181676 251272 181688
rect 170732 181648 251272 181676
rect 170732 181636 170738 181648
rect 251266 181636 251272 181648
rect 251324 181636 251330 181688
rect 251818 181636 251824 181688
rect 251876 181676 251882 181688
rect 341150 181676 341156 181688
rect 251876 181648 341156 181676
rect 251876 181636 251882 181648
rect 341150 181636 341156 181648
rect 341208 181636 341214 181688
rect 414658 181636 414664 181688
rect 414716 181676 414722 181688
rect 441614 181676 441620 181688
rect 414716 181648 441620 181676
rect 414716 181636 414722 181648
rect 441614 181636 441620 181648
rect 441672 181636 441678 181688
rect 457438 181636 457444 181688
rect 457496 181676 457502 181688
rect 474182 181676 474188 181688
rect 457496 181648 474188 181676
rect 457496 181636 457502 181648
rect 474182 181636 474188 181648
rect 474240 181636 474246 181688
rect 482278 181636 482284 181688
rect 482336 181676 482342 181688
rect 505278 181676 505284 181688
rect 482336 181648 505284 181676
rect 482336 181636 482342 181648
rect 505278 181636 505284 181648
rect 505336 181636 505342 181688
rect 159358 181568 159364 181620
rect 159416 181608 159422 181620
rect 209038 181608 209044 181620
rect 159416 181580 209044 181608
rect 159416 181568 159422 181580
rect 209038 181568 209044 181580
rect 209096 181568 209102 181620
rect 233878 181568 233884 181620
rect 233936 181608 233942 181620
rect 334158 181608 334164 181620
rect 233936 181580 334164 181608
rect 233936 181568 233942 181580
rect 334158 181568 334164 181580
rect 334216 181568 334222 181620
rect 352558 181568 352564 181620
rect 352616 181608 352622 181620
rect 448606 181608 448612 181620
rect 352616 181580 448612 181608
rect 352616 181568 352622 181580
rect 448606 181568 448612 181580
rect 448664 181568 448670 181620
rect 464338 181568 464344 181620
rect 464396 181608 464402 181620
rect 503990 181608 503996 181620
rect 464396 181580 503996 181608
rect 464396 181568 464402 181580
rect 503990 181568 503996 181580
rect 504048 181568 504054 181620
rect 137462 181500 137468 181552
rect 137520 181540 137526 181552
rect 249150 181540 249156 181552
rect 137520 181512 249156 181540
rect 137520 181500 137526 181512
rect 249150 181500 249156 181512
rect 249208 181500 249214 181552
rect 262858 181500 262864 181552
rect 262916 181540 262922 181552
rect 446398 181540 446404 181552
rect 262916 181512 446404 181540
rect 262916 181500 262922 181512
rect 446398 181500 446404 181512
rect 446456 181500 446462 181552
rect 449158 181500 449164 181552
rect 449216 181540 449222 181552
rect 502610 181540 502616 181552
rect 449216 181512 502616 181540
rect 449216 181500 449222 181512
rect 502610 181500 502616 181512
rect 502668 181500 502674 181552
rect 180610 181432 180616 181484
rect 180668 181472 180674 181484
rect 496998 181472 497004 181484
rect 180668 181444 497004 181472
rect 180668 181432 180674 181444
rect 496998 181432 497004 181444
rect 497056 181432 497062 181484
rect 130930 181024 130936 181076
rect 130988 181064 130994 181076
rect 166534 181064 166540 181076
rect 130988 181036 166540 181064
rect 130988 181024 130994 181036
rect 166534 181024 166540 181036
rect 166592 181024 166598 181076
rect 129458 180956 129464 181008
rect 129516 180996 129522 181008
rect 167914 180996 167920 181008
rect 129516 180968 167920 180996
rect 129516 180956 129522 180968
rect 167914 180956 167920 180968
rect 167972 180956 167978 181008
rect 121178 180888 121184 180940
rect 121236 180928 121242 180940
rect 167822 180928 167828 180940
rect 121236 180900 167828 180928
rect 121236 180888 121242 180900
rect 167822 180888 167828 180900
rect 167880 180888 167886 180940
rect 116946 180820 116952 180872
rect 117004 180860 117010 180872
rect 170858 180860 170864 180872
rect 117004 180832 170864 180860
rect 117004 180820 117010 180832
rect 170858 180820 170864 180832
rect 170916 180820 170922 180872
rect 246298 180412 246304 180464
rect 246356 180452 246362 180464
rect 272058 180452 272064 180464
rect 246356 180424 272064 180452
rect 246356 180412 246362 180424
rect 272058 180412 272064 180424
rect 272116 180412 272122 180464
rect 169202 180344 169208 180396
rect 169260 180384 169266 180396
rect 251358 180384 251364 180396
rect 169260 180356 251364 180384
rect 169260 180344 169266 180356
rect 251358 180344 251364 180356
rect 251416 180344 251422 180396
rect 151262 180276 151268 180328
rect 151320 180316 151326 180328
rect 266446 180316 266452 180328
rect 151320 180288 266452 180316
rect 151320 180276 151326 180288
rect 266446 180276 266452 180288
rect 266504 180276 266510 180328
rect 273898 180276 273904 180328
rect 273956 180316 273962 180328
rect 332870 180316 332876 180328
rect 273956 180288 332876 180316
rect 273956 180276 273962 180288
rect 332870 180276 332876 180288
rect 332928 180276 332934 180328
rect 490650 180276 490656 180328
rect 490708 180316 490714 180328
rect 501230 180316 501236 180328
rect 490708 180288 501236 180316
rect 490708 180276 490714 180288
rect 501230 180276 501236 180288
rect 501288 180276 501294 180328
rect 187050 180208 187056 180260
rect 187108 180248 187114 180260
rect 324498 180248 324504 180260
rect 187108 180220 324504 180248
rect 187108 180208 187114 180220
rect 324498 180208 324504 180220
rect 324556 180208 324562 180260
rect 411898 180208 411904 180260
rect 411956 180248 411962 180260
rect 506566 180248 506572 180260
rect 411956 180220 506572 180248
rect 411956 180208 411962 180220
rect 506566 180208 506572 180220
rect 506624 180208 506630 180260
rect 187142 180140 187148 180192
rect 187200 180180 187206 180192
rect 349246 180180 349252 180192
rect 187200 180152 349252 180180
rect 187200 180140 187206 180152
rect 349246 180140 349252 180152
rect 349304 180140 349310 180192
rect 359458 180140 359464 180192
rect 359516 180180 359522 180192
rect 509234 180180 509240 180192
rect 359516 180152 509240 180180
rect 359516 180140 359522 180152
rect 509234 180140 509240 180152
rect 509292 180140 509298 180192
rect 160738 180072 160744 180124
rect 160796 180112 160802 180124
rect 195238 180112 195244 180124
rect 160796 180084 195244 180112
rect 160796 180072 160802 180084
rect 195238 180072 195244 180084
rect 195296 180072 195302 180124
rect 222838 180072 222844 180124
rect 222896 180112 222902 180124
rect 503806 180112 503812 180124
rect 222896 180084 503812 180112
rect 222896 180072 222902 180084
rect 503806 180072 503812 180084
rect 503864 180072 503870 180124
rect 134702 179596 134708 179648
rect 134760 179636 134766 179648
rect 165430 179636 165436 179648
rect 134760 179608 165436 179636
rect 134760 179596 134766 179608
rect 165430 179596 165436 179608
rect 165488 179596 165494 179648
rect 126054 179528 126060 179580
rect 126112 179568 126118 179580
rect 168006 179568 168012 179580
rect 126112 179540 168012 179568
rect 126112 179528 126118 179540
rect 168006 179528 168012 179540
rect 168064 179528 168070 179580
rect 115842 179460 115848 179512
rect 115900 179500 115906 179512
rect 166258 179500 166264 179512
rect 115900 179472 166264 179500
rect 115900 179460 115906 179472
rect 166258 179460 166264 179472
rect 166316 179460 166322 179512
rect 109954 179392 109960 179444
rect 110012 179432 110018 179444
rect 169294 179432 169300 179444
rect 110012 179404 169300 179432
rect 110012 179392 110018 179404
rect 169294 179392 169300 179404
rect 169352 179392 169358 179444
rect 309870 178984 309876 179036
rect 309928 179024 309934 179036
rect 325970 179024 325976 179036
rect 309928 178996 325976 179024
rect 309928 178984 309934 178996
rect 325970 178984 325976 178996
rect 326028 178984 326034 179036
rect 170398 178916 170404 178968
rect 170456 178956 170462 178968
rect 251450 178956 251456 178968
rect 170456 178928 251456 178956
rect 170456 178916 170462 178928
rect 251450 178916 251456 178928
rect 251508 178916 251514 178968
rect 313918 178916 313924 178968
rect 313976 178956 313982 178968
rect 332686 178956 332692 178968
rect 313976 178928 332692 178956
rect 313976 178916 313982 178928
rect 332686 178916 332692 178928
rect 332744 178916 332750 178968
rect 244918 178848 244924 178900
rect 244976 178888 244982 178900
rect 336826 178888 336832 178900
rect 244976 178860 336832 178888
rect 244976 178848 244982 178860
rect 336826 178848 336832 178860
rect 336884 178848 336890 178900
rect 166350 178780 166356 178832
rect 166408 178820 166414 178832
rect 267918 178820 267924 178832
rect 166408 178792 267924 178820
rect 166408 178780 166414 178792
rect 267918 178780 267924 178792
rect 267976 178780 267982 178832
rect 295978 178780 295984 178832
rect 296036 178820 296042 178832
rect 327166 178820 327172 178832
rect 296036 178792 327172 178820
rect 296036 178780 296042 178792
rect 327166 178780 327172 178792
rect 327224 178780 327230 178832
rect 123478 178712 123484 178764
rect 123536 178752 123542 178764
rect 249334 178752 249340 178764
rect 123536 178724 249340 178752
rect 123536 178712 123542 178724
rect 249334 178712 249340 178724
rect 249392 178712 249398 178764
rect 257338 178712 257344 178764
rect 257396 178752 257402 178764
rect 346578 178752 346584 178764
rect 257396 178724 346584 178752
rect 257396 178712 257402 178724
rect 346578 178712 346584 178724
rect 346636 178712 346642 178764
rect 162118 178644 162124 178696
rect 162176 178684 162182 178696
rect 197998 178684 198004 178696
rect 162176 178656 198004 178684
rect 162176 178644 162182 178656
rect 197998 178644 198004 178656
rect 198056 178644 198062 178696
rect 202322 178644 202328 178696
rect 202380 178684 202386 178696
rect 339678 178684 339684 178696
rect 202380 178656 339684 178684
rect 202380 178644 202386 178656
rect 339678 178644 339684 178656
rect 339736 178644 339742 178696
rect 497458 178644 497464 178696
rect 497516 178684 497522 178696
rect 502518 178684 502524 178696
rect 497516 178656 502524 178684
rect 497516 178644 497522 178656
rect 502518 178644 502524 178656
rect 502576 178684 502582 178696
rect 503622 178684 503628 178696
rect 502576 178656 503628 178684
rect 502576 178644 502582 178656
rect 503622 178644 503628 178656
rect 503680 178644 503686 178696
rect 148226 178236 148232 178288
rect 148284 178276 148290 178288
rect 170490 178276 170496 178288
rect 148284 178248 170496 178276
rect 148284 178236 148290 178248
rect 170490 178236 170496 178248
rect 170548 178236 170554 178288
rect 114370 178168 114376 178220
rect 114428 178208 114434 178220
rect 166442 178208 166448 178220
rect 114428 178180 166448 178208
rect 114428 178168 114434 178180
rect 166442 178168 166448 178180
rect 166500 178168 166506 178220
rect 112254 178100 112260 178152
rect 112312 178140 112318 178152
rect 171962 178140 171968 178152
rect 112312 178112 171968 178140
rect 112312 178100 112318 178112
rect 171962 178100 171968 178112
rect 172020 178100 172026 178152
rect 97810 178032 97816 178084
rect 97868 178072 97874 178084
rect 177390 178072 177396 178084
rect 97868 178044 177396 178072
rect 97868 178032 97874 178044
rect 177390 178032 177396 178044
rect 177448 178032 177454 178084
rect 347038 178032 347044 178084
rect 347096 178072 347102 178084
rect 416774 178072 416780 178084
rect 347096 178044 416780 178072
rect 347096 178032 347102 178044
rect 416774 178032 416780 178044
rect 416832 178032 416838 178084
rect 503622 178032 503628 178084
rect 503680 178072 503686 178084
rect 580166 178072 580172 178084
rect 503680 178044 580172 178072
rect 503680 178032 503686 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 323670 177964 323676 178016
rect 323728 178004 323734 178016
rect 327074 178004 327080 178016
rect 323728 177976 327080 178004
rect 323728 177964 323734 177976
rect 327074 177964 327080 177976
rect 327132 177964 327138 178016
rect 242250 177624 242256 177676
rect 242308 177664 242314 177676
rect 256878 177664 256884 177676
rect 242308 177636 256884 177664
rect 242308 177624 242314 177636
rect 256878 177624 256884 177636
rect 256936 177624 256942 177676
rect 312538 177624 312544 177676
rect 312596 177664 312602 177676
rect 321738 177664 321744 177676
rect 312596 177636 321744 177664
rect 312596 177624 312602 177636
rect 321738 177624 321744 177636
rect 321796 177624 321802 177676
rect 226978 177556 226984 177608
rect 227036 177596 227042 177608
rect 249242 177596 249248 177608
rect 227036 177568 249248 177596
rect 227036 177556 227042 177568
rect 249242 177556 249248 177568
rect 249300 177556 249306 177608
rect 318702 177556 318708 177608
rect 318760 177596 318766 177608
rect 331398 177596 331404 177608
rect 318760 177568 331404 177596
rect 318760 177556 318766 177568
rect 331398 177556 331404 177568
rect 331456 177556 331462 177608
rect 231118 177488 231124 177540
rect 231176 177528 231182 177540
rect 258350 177528 258356 177540
rect 231176 177500 258356 177528
rect 231176 177488 231182 177500
rect 258350 177488 258356 177500
rect 258408 177488 258414 177540
rect 283558 177488 283564 177540
rect 283616 177528 283622 177540
rect 350626 177528 350632 177540
rect 283616 177500 350632 177528
rect 283616 177488 283622 177500
rect 350626 177488 350632 177500
rect 350684 177488 350690 177540
rect 190362 177420 190368 177472
rect 190420 177460 190426 177472
rect 294690 177460 294696 177472
rect 190420 177432 294696 177460
rect 190420 177420 190426 177432
rect 294690 177420 294696 177432
rect 294748 177420 294754 177472
rect 318058 177420 318064 177472
rect 318116 177460 318122 177472
rect 332778 177460 332784 177472
rect 318116 177432 332784 177460
rect 318116 177420 318122 177432
rect 332778 177420 332784 177432
rect 332836 177420 332842 177472
rect 202414 177352 202420 177404
rect 202472 177392 202478 177404
rect 323118 177392 323124 177404
rect 202472 177364 323124 177392
rect 202472 177352 202478 177364
rect 323118 177352 323124 177364
rect 323176 177352 323182 177404
rect 14458 177284 14464 177336
rect 14516 177324 14522 177336
rect 109678 177324 109684 177336
rect 14516 177296 109684 177324
rect 14516 177284 14522 177296
rect 109678 177284 109684 177296
rect 109736 177284 109742 177336
rect 203518 177284 203524 177336
rect 203576 177324 203582 177336
rect 338206 177324 338212 177336
rect 203576 177296 338212 177324
rect 203576 177284 203582 177296
rect 338206 177284 338212 177296
rect 338264 177284 338270 177336
rect 128170 177012 128176 177064
rect 128228 177052 128234 177064
rect 160094 177052 160100 177064
rect 128228 177024 160100 177052
rect 128228 177012 128234 177024
rect 160094 177012 160100 177024
rect 160152 177012 160158 177064
rect 124490 176944 124496 176996
rect 124548 176984 124554 176996
rect 165246 176984 165252 176996
rect 124548 176956 165252 176984
rect 124548 176944 124554 176956
rect 165246 176944 165252 176956
rect 165304 176944 165310 176996
rect 158898 176876 158904 176928
rect 158956 176916 158962 176928
rect 214742 176916 214748 176928
rect 158956 176888 214748 176916
rect 158956 176876 158962 176888
rect 214742 176876 214748 176888
rect 214800 176876 214806 176928
rect 108114 176808 108120 176860
rect 108172 176848 108178 176860
rect 169110 176848 169116 176860
rect 108172 176820 169116 176848
rect 108172 176808 108178 176820
rect 169110 176808 169116 176820
rect 169168 176808 169174 176860
rect 136082 176740 136088 176792
rect 136140 176780 136146 176792
rect 201586 176780 201592 176792
rect 136140 176752 201592 176780
rect 136140 176740 136146 176752
rect 201586 176740 201592 176752
rect 201644 176740 201650 176792
rect 496906 176740 496912 176792
rect 496964 176780 496970 176792
rect 501046 176780 501052 176792
rect 496964 176752 501052 176780
rect 496964 176740 496970 176752
rect 501046 176740 501052 176752
rect 501104 176740 501110 176792
rect 133138 176672 133144 176724
rect 133196 176712 133202 176724
rect 205634 176712 205640 176724
rect 133196 176684 205640 176712
rect 133196 176672 133202 176684
rect 205634 176672 205640 176684
rect 205692 176672 205698 176724
rect 342990 176672 342996 176724
rect 343048 176712 343054 176724
rect 416774 176712 416780 176724
rect 343048 176684 416780 176712
rect 343048 176672 343054 176684
rect 416774 176672 416780 176684
rect 416832 176672 416838 176724
rect 496814 176672 496820 176724
rect 496872 176712 496878 176724
rect 499758 176712 499764 176724
rect 496872 176684 499764 176712
rect 496872 176672 496878 176684
rect 499758 176672 499764 176684
rect 499816 176672 499822 176724
rect 201586 176604 201592 176656
rect 201644 176644 201650 176656
rect 213914 176644 213920 176656
rect 201644 176616 213920 176644
rect 201644 176604 201650 176616
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 313826 176604 313832 176656
rect 313884 176644 313890 176656
rect 321462 176644 321468 176656
rect 313884 176616 321468 176644
rect 313884 176604 313890 176616
rect 321462 176604 321468 176616
rect 321520 176604 321526 176656
rect 118418 176264 118424 176316
rect 118476 176304 118482 176316
rect 166350 176304 166356 176316
rect 118476 176276 166356 176304
rect 118476 176264 118482 176276
rect 166350 176264 166356 176276
rect 166408 176264 166414 176316
rect 163498 176196 163504 176248
rect 163556 176236 163562 176248
rect 211798 176236 211804 176248
rect 163556 176208 211804 176236
rect 163556 176196 163562 176208
rect 211798 176196 211804 176208
rect 211856 176196 211862 176248
rect 160094 176128 160100 176180
rect 160152 176168 160158 176180
rect 214098 176168 214104 176180
rect 160152 176140 214104 176168
rect 160152 176128 160158 176140
rect 214098 176128 214104 176140
rect 214156 176128 214162 176180
rect 102042 176060 102048 176112
rect 102100 176100 102106 176112
rect 171778 176100 171784 176112
rect 102100 176072 171784 176100
rect 102100 176060 102106 176072
rect 171778 176060 171784 176072
rect 171836 176060 171842 176112
rect 238110 176060 238116 176112
rect 238168 176100 238174 176112
rect 256694 176100 256700 176112
rect 238168 176072 256700 176100
rect 238168 176060 238174 176072
rect 256694 176060 256700 176072
rect 256752 176060 256758 176112
rect 307662 176060 307668 176112
rect 307720 176100 307726 176112
rect 349338 176100 349344 176112
rect 307720 176072 349344 176100
rect 307720 176060 307726 176072
rect 349338 176060 349344 176072
rect 349396 176060 349402 176112
rect 98362 175992 98368 176044
rect 98420 176032 98426 176044
rect 170398 176032 170404 176044
rect 98420 176004 170404 176032
rect 98420 175992 98426 176004
rect 170398 175992 170404 176004
rect 170456 175992 170462 176044
rect 171870 175992 171876 176044
rect 171928 176032 171934 176044
rect 258074 176032 258080 176044
rect 171928 176004 258080 176032
rect 171928 175992 171934 176004
rect 258074 175992 258080 176004
rect 258132 175992 258138 176044
rect 266998 175992 267004 176044
rect 267056 176032 267062 176044
rect 323026 176032 323032 176044
rect 267056 176004 323032 176032
rect 267056 175992 267062 176004
rect 323026 175992 323032 176004
rect 323084 175992 323090 176044
rect 121914 175924 121920 175976
rect 121972 175964 121978 175976
rect 195422 175964 195428 175976
rect 121972 175936 195428 175964
rect 121972 175924 121978 175936
rect 195422 175924 195428 175936
rect 195480 175924 195486 175976
rect 238018 175924 238024 175976
rect 238076 175964 238082 175976
rect 396718 175964 396724 175976
rect 238076 175936 396724 175964
rect 238076 175924 238082 175936
rect 396718 175924 396724 175936
rect 396776 175924 396782 175976
rect 240778 175788 240784 175840
rect 240836 175828 240842 175840
rect 248046 175828 248052 175840
rect 240836 175800 248052 175828
rect 240836 175788 240842 175800
rect 248046 175788 248052 175800
rect 248104 175788 248110 175840
rect 496814 175584 496820 175636
rect 496872 175624 496878 175636
rect 498470 175624 498476 175636
rect 496872 175596 498476 175624
rect 496872 175584 496878 175596
rect 498470 175584 498476 175596
rect 498528 175584 498534 175636
rect 165430 175176 165436 175228
rect 165488 175216 165494 175228
rect 213914 175216 213920 175228
rect 165488 175188 213920 175216
rect 165488 175176 165494 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 205634 175108 205640 175160
rect 205692 175148 205698 175160
rect 214006 175148 214012 175160
rect 205692 175120 214012 175148
rect 205692 175108 205698 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 252462 175108 252468 175160
rect 252520 175148 252526 175160
rect 258166 175148 258172 175160
rect 252520 175120 258172 175148
rect 252520 175108 252526 175120
rect 258166 175108 258172 175120
rect 258224 175108 258230 175160
rect 165246 174496 165252 174548
rect 165304 174536 165310 174548
rect 214926 174536 214932 174548
rect 165304 174508 214932 174536
rect 165304 174496 165310 174508
rect 214926 174496 214932 174508
rect 214984 174496 214990 174548
rect 284938 174020 284944 174072
rect 284996 174060 285002 174072
rect 307570 174060 307576 174072
rect 284996 174032 307576 174060
rect 284996 174020 285002 174032
rect 307570 174020 307576 174032
rect 307628 174020 307634 174072
rect 265802 173952 265808 174004
rect 265860 173992 265866 174004
rect 307662 173992 307668 174004
rect 265860 173964 307668 173992
rect 265860 173952 265866 173964
rect 307662 173952 307668 173964
rect 307720 173952 307726 174004
rect 263042 173884 263048 173936
rect 263100 173924 263106 173936
rect 307478 173924 307484 173936
rect 263100 173896 307484 173924
rect 263100 173884 263106 173896
rect 307478 173884 307484 173896
rect 307536 173884 307542 173936
rect 358078 173884 358084 173936
rect 358136 173924 358142 173936
rect 416774 173924 416780 173936
rect 358136 173896 416780 173924
rect 358136 173884 358142 173896
rect 416774 173884 416780 173896
rect 416832 173884 416838 173936
rect 164970 173816 164976 173868
rect 165028 173856 165034 173868
rect 213914 173856 213920 173868
rect 165028 173828 213920 173856
rect 165028 173816 165034 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 252462 173816 252468 173868
rect 252520 173856 252526 173868
rect 262398 173856 262404 173868
rect 252520 173828 262404 173856
rect 252520 173816 252526 173828
rect 262398 173816 262404 173828
rect 262456 173816 262462 173868
rect 166534 173748 166540 173800
rect 166592 173788 166598 173800
rect 214006 173788 214012 173800
rect 166592 173760 214012 173788
rect 166592 173748 166598 173760
rect 214006 173748 214012 173760
rect 214064 173748 214070 173800
rect 302878 172660 302884 172712
rect 302936 172700 302942 172712
rect 307478 172700 307484 172712
rect 302936 172672 307484 172700
rect 302936 172660 302942 172672
rect 307478 172660 307484 172672
rect 307536 172660 307542 172712
rect 298738 172592 298744 172644
rect 298796 172632 298802 172644
rect 307662 172632 307668 172644
rect 298796 172604 307668 172632
rect 298796 172592 298802 172604
rect 307662 172592 307668 172604
rect 307720 172592 307726 172644
rect 276750 172524 276756 172576
rect 276808 172564 276814 172576
rect 307294 172564 307300 172576
rect 276808 172536 307300 172564
rect 276808 172524 276814 172536
rect 307294 172524 307300 172536
rect 307352 172524 307358 172576
rect 167914 172456 167920 172508
rect 167972 172496 167978 172508
rect 213914 172496 213920 172508
rect 167972 172468 213920 172496
rect 167972 172456 167978 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 252370 172456 252376 172508
rect 252428 172496 252434 172508
rect 261018 172496 261024 172508
rect 252428 172468 261024 172496
rect 252428 172456 252434 172468
rect 261018 172456 261024 172468
rect 261076 172456 261082 172508
rect 252462 172116 252468 172168
rect 252520 172156 252526 172168
rect 258074 172156 258080 172168
rect 252520 172128 258080 172156
rect 252520 172116 252526 172128
rect 258074 172116 258080 172128
rect 258132 172116 258138 172168
rect 261478 171776 261484 171828
rect 261536 171816 261542 171828
rect 307386 171816 307392 171828
rect 261536 171788 307392 171816
rect 261536 171776 261542 171788
rect 307386 171776 307392 171788
rect 307444 171776 307450 171828
rect 278222 171164 278228 171216
rect 278280 171204 278286 171216
rect 307662 171204 307668 171216
rect 278280 171176 307668 171204
rect 278280 171164 278286 171176
rect 307662 171164 307668 171176
rect 307720 171164 307726 171216
rect 265710 171096 265716 171148
rect 265768 171136 265774 171148
rect 307110 171136 307116 171148
rect 265768 171108 307116 171136
rect 265768 171096 265774 171108
rect 307110 171096 307116 171108
rect 307168 171096 307174 171148
rect 324958 171096 324964 171148
rect 325016 171136 325022 171148
rect 327074 171136 327080 171148
rect 325016 171108 327080 171136
rect 325016 171096 325022 171108
rect 327074 171096 327080 171108
rect 327132 171096 327138 171148
rect 353938 171096 353944 171148
rect 353996 171136 354002 171148
rect 416774 171136 416780 171148
rect 353996 171108 416780 171136
rect 353996 171096 354002 171108
rect 416774 171096 416780 171108
rect 416832 171096 416838 171148
rect 168006 171028 168012 171080
rect 168064 171068 168070 171080
rect 214006 171068 214012 171080
rect 168064 171040 214012 171068
rect 168064 171028 168070 171040
rect 214006 171028 214012 171040
rect 214064 171028 214070 171080
rect 252462 171028 252468 171080
rect 252520 171068 252526 171080
rect 263594 171068 263600 171080
rect 252520 171040 263600 171068
rect 252520 171028 252526 171040
rect 263594 171028 263600 171040
rect 263652 171028 263658 171080
rect 180242 170960 180248 171012
rect 180300 171000 180306 171012
rect 213914 171000 213920 171012
rect 180300 170972 213920 171000
rect 180300 170960 180306 170972
rect 213914 170960 213920 170972
rect 213972 170960 213978 171012
rect 252370 170960 252376 171012
rect 252428 171000 252434 171012
rect 262306 171000 262312 171012
rect 252428 170972 262312 171000
rect 252428 170960 252434 170972
rect 262306 170960 262312 170972
rect 262364 170960 262370 171012
rect 252462 170552 252468 170604
rect 252520 170592 252526 170604
rect 256694 170592 256700 170604
rect 252520 170564 256700 170592
rect 252520 170552 252526 170564
rect 256694 170552 256700 170564
rect 256752 170552 256758 170604
rect 297450 169872 297456 169924
rect 297508 169912 297514 169924
rect 306742 169912 306748 169924
rect 297508 169884 306748 169912
rect 297508 169872 297514 169884
rect 306742 169872 306748 169884
rect 306800 169872 306806 169924
rect 267182 169804 267188 169856
rect 267240 169844 267246 169856
rect 307662 169844 307668 169856
rect 267240 169816 307668 169844
rect 267240 169804 267246 169816
rect 307662 169804 307668 169816
rect 307720 169804 307726 169856
rect 261662 169736 261668 169788
rect 261720 169776 261726 169788
rect 307478 169776 307484 169788
rect 261720 169748 307484 169776
rect 261720 169736 261726 169748
rect 307478 169736 307484 169748
rect 307536 169736 307542 169788
rect 324314 169668 324320 169720
rect 324372 169708 324378 169720
rect 335630 169708 335636 169720
rect 324372 169680 335636 169708
rect 324372 169668 324378 169680
rect 335630 169668 335636 169680
rect 335688 169668 335694 169720
rect 300302 168444 300308 168496
rect 300360 168484 300366 168496
rect 307662 168484 307668 168496
rect 300360 168456 307668 168484
rect 300360 168444 300366 168456
rect 307662 168444 307668 168456
rect 307720 168444 307726 168496
rect 258994 168376 259000 168428
rect 259052 168416 259058 168428
rect 307570 168416 307576 168428
rect 259052 168388 307576 168416
rect 259052 168376 259058 168388
rect 307570 168376 307576 168388
rect 307628 168376 307634 168428
rect 414658 168376 414664 168428
rect 414716 168416 414722 168428
rect 416774 168416 416780 168428
rect 414716 168388 416780 168416
rect 414716 168376 414722 168388
rect 416774 168376 416780 168388
rect 416832 168376 416838 168428
rect 167822 168308 167828 168360
rect 167880 168348 167886 168360
rect 214006 168348 214012 168360
rect 167880 168320 214012 168348
rect 167880 168308 167886 168320
rect 214006 168308 214012 168320
rect 214064 168308 214070 168360
rect 252370 168308 252376 168360
rect 252428 168348 252434 168360
rect 256878 168348 256884 168360
rect 252428 168320 256884 168348
rect 252428 168308 252434 168320
rect 256878 168308 256884 168320
rect 256936 168308 256942 168360
rect 324314 168308 324320 168360
rect 324372 168348 324378 168360
rect 357434 168348 357440 168360
rect 324372 168320 357440 168348
rect 324372 168308 324378 168320
rect 357434 168308 357440 168320
rect 357492 168308 357498 168360
rect 496814 168308 496820 168360
rect 496872 168348 496878 168360
rect 502426 168348 502432 168360
rect 496872 168320 502432 168348
rect 496872 168308 496878 168320
rect 502426 168308 502432 168320
rect 502484 168348 502490 168360
rect 503622 168348 503628 168360
rect 502484 168320 503628 168348
rect 502484 168308 502490 168320
rect 503622 168308 503628 168320
rect 503680 168308 503686 168360
rect 195422 168240 195428 168292
rect 195480 168280 195486 168292
rect 213914 168280 213920 168292
rect 195480 168252 213920 168280
rect 195480 168240 195486 168252
rect 213914 168240 213920 168252
rect 213972 168240 213978 168292
rect 252462 168036 252468 168088
rect 252520 168076 252526 168088
rect 259454 168076 259460 168088
rect 252520 168048 259460 168076
rect 252520 168036 252526 168048
rect 259454 168036 259460 168048
rect 259512 168036 259518 168088
rect 291930 167628 291936 167680
rect 291988 167668 291994 167680
rect 306558 167668 306564 167680
rect 291988 167640 306564 167668
rect 291988 167628 291994 167640
rect 306558 167628 306564 167640
rect 306616 167628 306622 167680
rect 338758 167628 338764 167680
rect 338816 167668 338822 167680
rect 348418 167668 348424 167680
rect 338816 167640 348424 167668
rect 338816 167628 338822 167640
rect 348418 167628 348424 167640
rect 348476 167628 348482 167680
rect 503622 167628 503628 167680
rect 503680 167668 503686 167680
rect 542998 167668 543004 167680
rect 503680 167640 543004 167668
rect 503680 167628 503686 167640
rect 542998 167628 543004 167640
rect 543056 167628 543062 167680
rect 251266 167220 251272 167272
rect 251324 167260 251330 167272
rect 251542 167260 251548 167272
rect 251324 167232 251548 167260
rect 251324 167220 251330 167232
rect 251542 167220 251548 167232
rect 251600 167220 251606 167272
rect 268378 167084 268384 167136
rect 268436 167124 268442 167136
rect 307662 167124 307668 167136
rect 268436 167096 307668 167124
rect 268436 167084 268442 167096
rect 307662 167084 307668 167096
rect 307720 167084 307726 167136
rect 264422 167016 264428 167068
rect 264480 167056 264486 167068
rect 307294 167056 307300 167068
rect 264480 167028 307300 167056
rect 264480 167016 264486 167028
rect 307294 167016 307300 167028
rect 307352 167016 307358 167068
rect 166350 166948 166356 167000
rect 166408 166988 166414 167000
rect 214098 166988 214104 167000
rect 166408 166960 214104 166988
rect 166408 166948 166414 166960
rect 214098 166948 214104 166960
rect 214156 166948 214162 167000
rect 170858 166880 170864 166932
rect 170916 166920 170922 166932
rect 214006 166920 214012 166932
rect 170916 166892 214012 166920
rect 170916 166880 170922 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 204990 166812 204996 166864
rect 205048 166852 205054 166864
rect 213914 166852 213920 166864
rect 205048 166824 213920 166852
rect 205048 166812 205054 166824
rect 213914 166812 213920 166824
rect 213972 166812 213978 166864
rect 252370 166676 252376 166728
rect 252428 166716 252434 166728
rect 258258 166716 258264 166728
rect 252428 166688 258264 166716
rect 252428 166676 252434 166688
rect 258258 166676 258264 166688
rect 258316 166676 258322 166728
rect 252462 166608 252468 166660
rect 252520 166648 252526 166660
rect 258350 166648 258356 166660
rect 252520 166620 258356 166648
rect 252520 166608 252526 166620
rect 258350 166608 258356 166620
rect 258408 166608 258414 166660
rect 295978 166336 295984 166388
rect 296036 166376 296042 166388
rect 306650 166376 306656 166388
rect 296036 166348 306656 166376
rect 296036 166336 296042 166348
rect 306650 166336 306656 166348
rect 306708 166336 306714 166388
rect 264330 166268 264336 166320
rect 264388 166308 264394 166320
rect 306926 166308 306932 166320
rect 264388 166280 306932 166308
rect 264388 166268 264394 166280
rect 306926 166268 306932 166280
rect 306984 166268 306990 166320
rect 496814 166268 496820 166320
rect 496872 166308 496878 166320
rect 504082 166308 504088 166320
rect 496872 166280 504088 166308
rect 496872 166268 496878 166280
rect 504082 166268 504088 166280
rect 504140 166268 504146 166320
rect 252462 166064 252468 166116
rect 252520 166104 252526 166116
rect 259730 166104 259736 166116
rect 252520 166076 259736 166104
rect 252520 166064 252526 166076
rect 259730 166064 259736 166076
rect 259788 166064 259794 166116
rect 271138 165588 271144 165640
rect 271196 165628 271202 165640
rect 306742 165628 306748 165640
rect 271196 165600 306748 165628
rect 271196 165588 271202 165600
rect 306742 165588 306748 165600
rect 306800 165588 306806 165640
rect 338758 165588 338764 165640
rect 338816 165628 338822 165640
rect 416774 165628 416780 165640
rect 338816 165600 416780 165628
rect 338816 165588 338822 165600
rect 416774 165588 416780 165600
rect 416832 165588 416838 165640
rect 504082 165588 504088 165640
rect 504140 165628 504146 165640
rect 525058 165628 525064 165640
rect 504140 165600 525064 165628
rect 504140 165588 504146 165600
rect 525058 165588 525064 165600
rect 525116 165588 525122 165640
rect 535454 165588 535460 165640
rect 535512 165628 535518 165640
rect 580166 165628 580172 165640
rect 535512 165600 580172 165628
rect 535512 165588 535518 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 166258 165520 166264 165572
rect 166316 165560 166322 165572
rect 213914 165560 213920 165572
rect 166316 165532 213920 165560
rect 166316 165520 166322 165532
rect 213914 165520 213920 165532
rect 213972 165520 213978 165572
rect 252462 165520 252468 165572
rect 252520 165560 252526 165572
rect 259546 165560 259552 165572
rect 252520 165532 259552 165560
rect 252520 165520 252526 165532
rect 259546 165520 259552 165532
rect 259604 165520 259610 165572
rect 324314 165520 324320 165572
rect 324372 165560 324378 165572
rect 339678 165560 339684 165572
rect 324372 165532 339684 165560
rect 324372 165520 324378 165532
rect 339678 165520 339684 165532
rect 339736 165520 339742 165572
rect 166442 165452 166448 165504
rect 166500 165492 166506 165504
rect 214006 165492 214012 165504
rect 166500 165464 214012 165492
rect 166500 165452 166506 165464
rect 214006 165452 214012 165464
rect 214064 165452 214070 165504
rect 252370 165452 252376 165504
rect 252428 165492 252434 165504
rect 256786 165492 256792 165504
rect 252428 165464 256792 165492
rect 252428 165452 252434 165464
rect 256786 165452 256792 165464
rect 256844 165452 256850 165504
rect 324406 165452 324412 165504
rect 324464 165492 324470 165504
rect 332870 165492 332876 165504
rect 324464 165464 332876 165492
rect 324464 165452 324470 165464
rect 332870 165452 332876 165464
rect 332928 165452 332934 165504
rect 258718 164840 258724 164892
rect 258776 164880 258782 164892
rect 307478 164880 307484 164892
rect 258776 164852 307484 164880
rect 258776 164840 258782 164852
rect 307478 164840 307484 164852
rect 307536 164840 307542 164892
rect 496814 164840 496820 164892
rect 496872 164880 496878 164892
rect 503990 164880 503996 164892
rect 496872 164852 503996 164880
rect 496872 164840 496878 164852
rect 503990 164840 503996 164852
rect 504048 164840 504054 164892
rect 301590 164296 301596 164348
rect 301648 164336 301654 164348
rect 307110 164336 307116 164348
rect 301648 164308 307116 164336
rect 301648 164296 301654 164308
rect 307110 164296 307116 164308
rect 307168 164296 307174 164348
rect 269850 164228 269856 164280
rect 269908 164268 269914 164280
rect 307662 164268 307668 164280
rect 269908 164240 307668 164268
rect 269908 164228 269914 164240
rect 307662 164228 307668 164240
rect 307720 164228 307726 164280
rect 359458 164228 359464 164280
rect 359516 164268 359522 164280
rect 416774 164268 416780 164280
rect 359516 164240 416780 164268
rect 359516 164228 359522 164240
rect 416774 164228 416780 164240
rect 416832 164228 416838 164280
rect 496354 164228 496360 164280
rect 496412 164268 496418 164280
rect 530578 164268 530584 164280
rect 496412 164240 530584 164268
rect 496412 164228 496418 164240
rect 530578 164228 530584 164240
rect 530636 164228 530642 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 33778 164200 33784 164212
rect 3292 164172 33784 164200
rect 3292 164160 3298 164172
rect 33778 164160 33784 164172
rect 33836 164160 33842 164212
rect 171962 164160 171968 164212
rect 172020 164200 172026 164212
rect 213914 164200 213920 164212
rect 172020 164172 213920 164200
rect 172020 164160 172026 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 252462 164160 252468 164212
rect 252520 164200 252526 164212
rect 270494 164200 270500 164212
rect 252520 164172 270500 164200
rect 252520 164160 252526 164172
rect 270494 164160 270500 164172
rect 270552 164160 270558 164212
rect 324314 164160 324320 164212
rect 324372 164200 324378 164212
rect 334158 164200 334164 164212
rect 324372 164172 334164 164200
rect 324372 164160 324378 164172
rect 334158 164160 334164 164172
rect 334216 164160 334222 164212
rect 496814 164160 496820 164212
rect 496872 164200 496878 164212
rect 509326 164200 509332 164212
rect 496872 164172 509332 164200
rect 496872 164160 496878 164172
rect 509326 164160 509332 164172
rect 509384 164200 509390 164212
rect 535454 164200 535460 164212
rect 509384 164172 535460 164200
rect 509384 164160 509390 164172
rect 535454 164160 535460 164172
rect 535512 164160 535518 164212
rect 252370 164092 252376 164144
rect 252428 164132 252434 164144
rect 263778 164132 263784 164144
rect 252428 164104 263784 164132
rect 252428 164092 252434 164104
rect 263778 164092 263784 164104
rect 263836 164092 263842 164144
rect 324406 164092 324412 164144
rect 324464 164132 324470 164144
rect 331490 164132 331496 164144
rect 324464 164104 331496 164132
rect 324464 164092 324470 164104
rect 331490 164092 331496 164104
rect 331548 164092 331554 164144
rect 272518 163548 272524 163600
rect 272576 163588 272582 163600
rect 306558 163588 306564 163600
rect 272576 163560 306564 163588
rect 272576 163548 272582 163560
rect 306558 163548 306564 163560
rect 306616 163548 306622 163600
rect 257614 163480 257620 163532
rect 257672 163520 257678 163532
rect 307570 163520 307576 163532
rect 257672 163492 307576 163520
rect 257672 163480 257678 163492
rect 307570 163480 307576 163492
rect 307628 163480 307634 163532
rect 293310 162868 293316 162920
rect 293368 162908 293374 162920
rect 307662 162908 307668 162920
rect 293368 162880 307668 162908
rect 293368 162868 293374 162880
rect 307662 162868 307668 162880
rect 307720 162868 307726 162920
rect 340138 162868 340144 162920
rect 340196 162908 340202 162920
rect 416774 162908 416780 162920
rect 340196 162880 416780 162908
rect 340196 162868 340202 162880
rect 416774 162868 416780 162880
rect 416832 162868 416838 162920
rect 169294 162800 169300 162852
rect 169352 162840 169358 162852
rect 214006 162840 214012 162852
rect 169352 162812 214012 162840
rect 169352 162800 169358 162812
rect 214006 162800 214012 162812
rect 214064 162800 214070 162852
rect 252370 162800 252376 162852
rect 252428 162840 252434 162852
rect 266538 162840 266544 162852
rect 252428 162812 266544 162840
rect 252428 162800 252434 162812
rect 266538 162800 266544 162812
rect 266596 162800 266602 162852
rect 324314 162800 324320 162852
rect 324372 162840 324378 162852
rect 334066 162840 334072 162852
rect 324372 162812 334072 162840
rect 324372 162800 324378 162812
rect 334066 162800 334072 162812
rect 334124 162800 334130 162852
rect 496814 162800 496820 162852
rect 496872 162840 496878 162852
rect 515398 162840 515404 162852
rect 496872 162812 515404 162840
rect 496872 162800 496878 162812
rect 515398 162800 515404 162812
rect 515456 162800 515462 162852
rect 196802 162732 196808 162784
rect 196860 162772 196866 162784
rect 213914 162772 213920 162784
rect 196860 162744 213920 162772
rect 196860 162732 196866 162744
rect 213914 162732 213920 162744
rect 213972 162732 213978 162784
rect 252462 162732 252468 162784
rect 252520 162772 252526 162784
rect 264974 162772 264980 162784
rect 252520 162744 264980 162772
rect 252520 162732 252526 162744
rect 264974 162732 264980 162744
rect 265032 162732 265038 162784
rect 302970 161644 302976 161696
rect 303028 161684 303034 161696
rect 307386 161684 307392 161696
rect 303028 161656 307392 161684
rect 303028 161644 303034 161656
rect 307386 161644 307392 161656
rect 307444 161644 307450 161696
rect 299014 161576 299020 161628
rect 299072 161616 299078 161628
rect 307478 161616 307484 161628
rect 299072 161588 307484 161616
rect 299072 161576 299078 161588
rect 307478 161576 307484 161588
rect 307536 161576 307542 161628
rect 269942 161508 269948 161560
rect 270000 161548 270006 161560
rect 307570 161548 307576 161560
rect 270000 161520 307576 161548
rect 270000 161508 270006 161520
rect 307570 161508 307576 161520
rect 307628 161508 307634 161560
rect 262858 161440 262864 161492
rect 262916 161480 262922 161492
rect 307662 161480 307668 161492
rect 262916 161452 307668 161480
rect 262916 161440 262922 161452
rect 307662 161440 307668 161452
rect 307720 161440 307726 161492
rect 334802 161440 334808 161492
rect 334860 161480 334866 161492
rect 416774 161480 416780 161492
rect 334860 161452 416780 161480
rect 334860 161440 334866 161452
rect 416774 161440 416780 161452
rect 416832 161440 416838 161492
rect 169110 161372 169116 161424
rect 169168 161412 169174 161424
rect 213914 161412 213920 161424
rect 169168 161384 213920 161412
rect 169168 161372 169174 161384
rect 213914 161372 213920 161384
rect 213972 161372 213978 161424
rect 252462 161372 252468 161424
rect 252520 161412 252526 161424
rect 263686 161412 263692 161424
rect 252520 161384 263692 161412
rect 252520 161372 252526 161384
rect 263686 161372 263692 161384
rect 263744 161372 263750 161424
rect 496906 161372 496912 161424
rect 496964 161412 496970 161424
rect 512086 161412 512092 161424
rect 496964 161384 512092 161412
rect 496964 161372 496970 161384
rect 512086 161372 512092 161384
rect 512144 161372 512150 161424
rect 196710 161304 196716 161356
rect 196768 161344 196774 161356
rect 214006 161344 214012 161356
rect 196768 161316 214012 161344
rect 196768 161304 196774 161316
rect 214006 161304 214012 161316
rect 214064 161304 214070 161356
rect 252370 160488 252376 160540
rect 252428 160528 252434 160540
rect 259638 160528 259644 160540
rect 252428 160500 259644 160528
rect 252428 160488 252434 160500
rect 259638 160488 259644 160500
rect 259696 160488 259702 160540
rect 287974 160216 287980 160268
rect 288032 160256 288038 160268
rect 307570 160256 307576 160268
rect 288032 160228 307576 160256
rect 288032 160216 288038 160228
rect 307570 160216 307576 160228
rect 307628 160216 307634 160268
rect 260466 160148 260472 160200
rect 260524 160188 260530 160200
rect 307662 160188 307668 160200
rect 260524 160160 307668 160188
rect 260524 160148 260530 160160
rect 307662 160148 307668 160160
rect 307720 160148 307726 160200
rect 260098 160080 260104 160132
rect 260156 160120 260162 160132
rect 306558 160120 306564 160132
rect 260156 160092 306564 160120
rect 260156 160080 260162 160092
rect 306558 160080 306564 160092
rect 306616 160080 306622 160132
rect 167730 160012 167736 160064
rect 167788 160052 167794 160064
rect 214006 160052 214012 160064
rect 167788 160024 214012 160052
rect 167788 160012 167794 160024
rect 214006 160012 214012 160024
rect 214064 160012 214070 160064
rect 252462 160012 252468 160064
rect 252520 160052 252526 160064
rect 273438 160052 273444 160064
rect 252520 160024 273444 160052
rect 252520 160012 252526 160024
rect 273438 160012 273444 160024
rect 273496 160012 273502 160064
rect 496906 160012 496912 160064
rect 496964 160052 496970 160064
rect 536834 160052 536840 160064
rect 496964 160024 536840 160052
rect 496964 160012 496970 160024
rect 536834 160012 536840 160024
rect 536892 160012 536898 160064
rect 170766 159944 170772 159996
rect 170824 159984 170830 159996
rect 213914 159984 213920 159996
rect 170824 159956 213920 159984
rect 170824 159944 170830 159956
rect 213914 159944 213920 159956
rect 213972 159944 213978 159996
rect 496998 159944 497004 159996
rect 497056 159984 497062 159996
rect 503714 159984 503720 159996
rect 497056 159956 503720 159984
rect 497056 159944 497062 159956
rect 503714 159944 503720 159956
rect 503772 159944 503778 159996
rect 273898 158856 273904 158908
rect 273956 158896 273962 158908
rect 306926 158896 306932 158908
rect 273956 158868 306932 158896
rect 273956 158856 273962 158868
rect 306926 158856 306932 158868
rect 306984 158856 306990 158908
rect 264514 158788 264520 158840
rect 264572 158828 264578 158840
rect 307662 158828 307668 158840
rect 264572 158800 307668 158828
rect 264572 158788 264578 158800
rect 307662 158788 307668 158800
rect 307720 158788 307726 158840
rect 260374 158720 260380 158772
rect 260432 158760 260438 158772
rect 307570 158760 307576 158772
rect 260432 158732 307576 158760
rect 260432 158720 260438 158732
rect 307570 158720 307576 158732
rect 307628 158720 307634 158772
rect 344278 158720 344284 158772
rect 344336 158760 344342 158772
rect 416774 158760 416780 158772
rect 344336 158732 416780 158760
rect 344336 158720 344342 158732
rect 416774 158720 416780 158732
rect 416832 158720 416838 158772
rect 171778 158652 171784 158704
rect 171836 158692 171842 158704
rect 213914 158692 213920 158704
rect 171836 158664 213920 158692
rect 171836 158652 171842 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 252462 158652 252468 158704
rect 252520 158692 252526 158704
rect 260926 158692 260932 158704
rect 252520 158664 260932 158692
rect 252520 158652 252526 158664
rect 260926 158652 260932 158664
rect 260984 158652 260990 158704
rect 324406 158652 324412 158704
rect 324464 158692 324470 158704
rect 335446 158692 335452 158704
rect 324464 158664 335452 158692
rect 324464 158652 324470 158664
rect 335446 158652 335452 158664
rect 335504 158652 335510 158704
rect 496906 158652 496912 158704
rect 496964 158692 496970 158704
rect 517606 158692 517612 158704
rect 496964 158664 517612 158692
rect 496964 158652 496970 158664
rect 517606 158652 517612 158664
rect 517664 158692 517670 158704
rect 544378 158692 544384 158704
rect 517664 158664 544384 158692
rect 517664 158652 517670 158664
rect 544378 158652 544384 158664
rect 544436 158652 544442 158704
rect 324314 158516 324320 158568
rect 324372 158556 324378 158568
rect 327442 158556 327448 158568
rect 324372 158528 327448 158556
rect 324372 158516 324378 158528
rect 327442 158516 327448 158528
rect 327500 158516 327506 158568
rect 253382 157972 253388 158024
rect 253440 158012 253446 158024
rect 307202 158012 307208 158024
rect 253440 157984 307208 158012
rect 253440 157972 253446 157984
rect 307202 157972 307208 157984
rect 307260 157972 307266 158024
rect 283558 157428 283564 157480
rect 283616 157468 283622 157480
rect 307478 157468 307484 157480
rect 283616 157440 307484 157468
rect 283616 157428 283622 157440
rect 307478 157428 307484 157440
rect 307536 157428 307542 157480
rect 257338 157360 257344 157412
rect 257396 157400 257402 157412
rect 306742 157400 306748 157412
rect 257396 157372 306748 157400
rect 257396 157360 257402 157372
rect 306742 157360 306748 157372
rect 306800 157360 306806 157412
rect 169018 157292 169024 157344
rect 169076 157332 169082 157344
rect 213914 157332 213920 157344
rect 169076 157304 213920 157332
rect 169076 157292 169082 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 252462 157292 252468 157344
rect 252520 157332 252526 157344
rect 270678 157332 270684 157344
rect 252520 157304 270684 157332
rect 252520 157292 252526 157304
rect 270678 157292 270684 157304
rect 270736 157292 270742 157344
rect 496906 157292 496912 157344
rect 496964 157332 496970 157344
rect 582374 157332 582380 157344
rect 496964 157304 582380 157332
rect 496964 157292 496970 157304
rect 582374 157292 582380 157304
rect 582432 157292 582438 157344
rect 173158 157224 173164 157276
rect 173216 157264 173222 157276
rect 214006 157264 214012 157276
rect 173216 157236 214012 157264
rect 173216 157224 173222 157236
rect 214006 157224 214012 157236
rect 214064 157224 214070 157276
rect 253198 156612 253204 156664
rect 253256 156652 253262 156664
rect 267826 156652 267832 156664
rect 253256 156624 267832 156652
rect 253256 156612 253262 156624
rect 267826 156612 267832 156624
rect 267884 156612 267890 156664
rect 324314 156408 324320 156460
rect 324372 156448 324378 156460
rect 327258 156448 327264 156460
rect 324372 156420 327264 156448
rect 324372 156408 324378 156420
rect 327258 156408 327264 156420
rect 327316 156408 327322 156460
rect 281074 156068 281080 156120
rect 281132 156108 281138 156120
rect 307662 156108 307668 156120
rect 281132 156080 307668 156108
rect 281132 156068 281138 156080
rect 307662 156068 307668 156080
rect 307720 156068 307726 156120
rect 266998 156000 267004 156052
rect 267056 156040 267062 156052
rect 307570 156040 307576 156052
rect 267056 156012 307576 156040
rect 267056 156000 267062 156012
rect 307570 156000 307576 156012
rect 307628 156000 307634 156052
rect 260282 155932 260288 155984
rect 260340 155972 260346 155984
rect 306558 155972 306564 155984
rect 260340 155944 306564 155972
rect 260340 155932 260346 155944
rect 306558 155932 306564 155944
rect 306616 155932 306622 155984
rect 335998 155932 336004 155984
rect 336056 155972 336062 155984
rect 416774 155972 416780 155984
rect 336056 155944 416780 155972
rect 336056 155932 336062 155944
rect 416774 155932 416780 155944
rect 416832 155932 416838 155984
rect 170398 155864 170404 155916
rect 170456 155904 170462 155916
rect 213914 155904 213920 155916
rect 170456 155876 213920 155904
rect 170456 155864 170462 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 252462 155864 252468 155916
rect 252520 155904 252526 155916
rect 265066 155904 265072 155916
rect 252520 155876 265072 155904
rect 252520 155864 252526 155876
rect 265066 155864 265072 155876
rect 265124 155864 265130 155916
rect 496906 155864 496912 155916
rect 496964 155904 496970 155916
rect 519538 155904 519544 155916
rect 496964 155876 519544 155904
rect 496964 155864 496970 155876
rect 519538 155864 519544 155876
rect 519596 155864 519602 155916
rect 177390 155796 177396 155848
rect 177448 155836 177454 155848
rect 214006 155836 214012 155848
rect 177448 155808 214012 155836
rect 177448 155796 177454 155808
rect 214006 155796 214012 155808
rect 214064 155796 214070 155848
rect 252370 155796 252376 155848
rect 252428 155836 252434 155848
rect 255406 155836 255412 155848
rect 252428 155808 255412 155836
rect 252428 155796 252434 155808
rect 255406 155796 255412 155808
rect 255464 155796 255470 155848
rect 327718 155184 327724 155236
rect 327776 155224 327782 155236
rect 333974 155224 333980 155236
rect 327776 155196 333980 155224
rect 327776 155184 327782 155196
rect 333974 155184 333980 155196
rect 334032 155184 334038 155236
rect 304350 154708 304356 154760
rect 304408 154748 304414 154760
rect 307662 154748 307668 154760
rect 304408 154720 307668 154748
rect 304408 154708 304414 154720
rect 307662 154708 307668 154720
rect 307720 154708 307726 154760
rect 271230 154640 271236 154692
rect 271288 154680 271294 154692
rect 306558 154680 306564 154692
rect 271288 154652 306564 154680
rect 271288 154640 271294 154652
rect 306558 154640 306564 154652
rect 306616 154640 306622 154692
rect 261754 154572 261760 154624
rect 261812 154612 261818 154624
rect 307294 154612 307300 154624
rect 261812 154584 307300 154612
rect 261812 154572 261818 154584
rect 307294 154572 307300 154584
rect 307352 154572 307358 154624
rect 332042 154572 332048 154624
rect 332100 154612 332106 154624
rect 416774 154612 416780 154624
rect 332100 154584 416780 154612
rect 332100 154572 332106 154584
rect 416774 154572 416780 154584
rect 416832 154572 416838 154624
rect 252462 154504 252468 154556
rect 252520 154544 252526 154556
rect 274726 154544 274732 154556
rect 252520 154516 274732 154544
rect 252520 154504 252526 154516
rect 274726 154504 274732 154516
rect 274784 154504 274790 154556
rect 324406 154504 324412 154556
rect 324464 154544 324470 154556
rect 332778 154544 332784 154556
rect 324464 154516 332784 154544
rect 324464 154504 324470 154516
rect 332778 154504 332784 154516
rect 332836 154504 332842 154556
rect 496998 154504 497004 154556
rect 497056 154544 497062 154556
rect 505278 154544 505284 154556
rect 497056 154516 505284 154544
rect 497056 154504 497062 154516
rect 505278 154504 505284 154516
rect 505336 154504 505342 154556
rect 251450 154436 251456 154488
rect 251508 154476 251514 154488
rect 254210 154476 254216 154488
rect 251508 154448 254216 154476
rect 251508 154436 251514 154448
rect 254210 154436 254216 154448
rect 254268 154436 254274 154488
rect 324314 154436 324320 154488
rect 324372 154476 324378 154488
rect 328730 154476 328736 154488
rect 324372 154448 328736 154476
rect 324372 154436 324378 154448
rect 328730 154436 328736 154448
rect 328788 154436 328794 154488
rect 496906 154436 496912 154488
rect 496964 154476 496970 154488
rect 502610 154476 502616 154488
rect 496964 154448 502616 154476
rect 496964 154436 496970 154448
rect 502610 154436 502616 154448
rect 502668 154436 502674 154488
rect 167638 153824 167644 153876
rect 167696 153864 167702 153876
rect 208394 153864 208400 153876
rect 167696 153836 208400 153864
rect 167696 153824 167702 153836
rect 208394 153824 208400 153836
rect 208452 153824 208458 153876
rect 275370 153348 275376 153400
rect 275428 153388 275434 153400
rect 307570 153388 307576 153400
rect 275428 153360 307576 153388
rect 275428 153348 275434 153360
rect 307570 153348 307576 153360
rect 307628 153348 307634 153400
rect 258810 153280 258816 153332
rect 258868 153320 258874 153332
rect 307662 153320 307668 153332
rect 258868 153292 307668 153320
rect 258868 153280 258874 153292
rect 307662 153280 307668 153292
rect 307720 153280 307726 153332
rect 173158 153212 173164 153264
rect 173216 153252 173222 153264
rect 213914 153252 213920 153264
rect 173216 153224 213920 153252
rect 173216 153212 173222 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 258902 153212 258908 153264
rect 258960 153252 258966 153264
rect 307294 153252 307300 153264
rect 258960 153224 307300 153252
rect 258960 153212 258966 153224
rect 307294 153212 307300 153224
rect 307352 153212 307358 153264
rect 356790 153212 356796 153264
rect 356848 153252 356854 153264
rect 416774 153252 416780 153264
rect 356848 153224 416780 153252
rect 356848 153212 356854 153224
rect 416774 153212 416780 153224
rect 416832 153212 416838 153264
rect 252278 153144 252284 153196
rect 252336 153184 252342 153196
rect 271966 153184 271972 153196
rect 252336 153156 271972 153184
rect 252336 153144 252342 153156
rect 271966 153144 271972 153156
rect 272024 153144 272030 153196
rect 324314 153144 324320 153196
rect 324372 153184 324378 153196
rect 330018 153184 330024 153196
rect 324372 153156 330024 153184
rect 324372 153144 324378 153156
rect 330018 153144 330024 153156
rect 330076 153144 330082 153196
rect 496906 153144 496912 153196
rect 496964 153184 496970 153196
rect 507946 153184 507952 153196
rect 496964 153156 507952 153184
rect 496964 153144 496970 153156
rect 507946 153144 507952 153156
rect 508004 153144 508010 153196
rect 252462 153076 252468 153128
rect 252520 153116 252526 153128
rect 269206 153116 269212 153128
rect 252520 153088 269212 153116
rect 252520 153076 252526 153088
rect 269206 153076 269212 153088
rect 269264 153076 269270 153128
rect 252370 153008 252376 153060
rect 252428 153048 252434 153060
rect 267918 153048 267924 153060
rect 252428 153020 267924 153048
rect 252428 153008 252434 153020
rect 267918 153008 267924 153020
rect 267976 153008 267982 153060
rect 296070 151920 296076 151972
rect 296128 151960 296134 151972
rect 307662 151960 307668 151972
rect 296128 151932 307668 151960
rect 296128 151920 296134 151932
rect 307662 151920 307668 151932
rect 307720 151920 307726 151972
rect 206370 151852 206376 151904
rect 206428 151892 206434 151904
rect 213914 151892 213920 151904
rect 206428 151864 213920 151892
rect 206428 151852 206434 151864
rect 213914 151852 213920 151864
rect 213972 151852 213978 151904
rect 268470 151852 268476 151904
rect 268528 151892 268534 151904
rect 307570 151892 307576 151904
rect 268528 151864 307576 151892
rect 268528 151852 268534 151864
rect 307570 151852 307576 151864
rect 307628 151852 307634 151904
rect 199378 151784 199384 151836
rect 199436 151824 199442 151836
rect 214006 151824 214012 151836
rect 199436 151796 214012 151824
rect 199436 151784 199442 151796
rect 214006 151784 214012 151796
rect 214064 151784 214070 151836
rect 254578 151784 254584 151836
rect 254636 151824 254642 151836
rect 307478 151824 307484 151836
rect 254636 151796 307484 151824
rect 254636 151784 254642 151796
rect 307478 151784 307484 151796
rect 307536 151784 307542 151836
rect 324406 151716 324412 151768
rect 324464 151756 324470 151768
rect 347866 151756 347872 151768
rect 324464 151728 347872 151756
rect 324464 151716 324470 151728
rect 347866 151716 347872 151728
rect 347924 151716 347930 151768
rect 324314 151648 324320 151700
rect 324372 151688 324378 151700
rect 330110 151688 330116 151700
rect 324372 151660 330116 151688
rect 324372 151648 324378 151660
rect 330110 151648 330116 151660
rect 330168 151648 330174 151700
rect 252462 151444 252468 151496
rect 252520 151484 252526 151496
rect 255590 151484 255596 151496
rect 252520 151456 255596 151484
rect 252520 151444 252526 151456
rect 255590 151444 255596 151456
rect 255648 151444 255654 151496
rect 251450 151308 251456 151360
rect 251508 151348 251514 151360
rect 254118 151348 254124 151360
rect 251508 151320 254124 151348
rect 251508 151308 251514 151320
rect 254118 151308 254124 151320
rect 254176 151308 254182 151360
rect 251818 151104 251824 151156
rect 251876 151144 251882 151156
rect 283558 151144 283564 151156
rect 251876 151116 283564 151144
rect 251876 151104 251882 151116
rect 283558 151104 283564 151116
rect 283616 151104 283622 151156
rect 255958 151036 255964 151088
rect 256016 151076 256022 151088
rect 306650 151076 306656 151088
rect 256016 151048 306656 151076
rect 256016 151036 256022 151048
rect 306650 151036 306656 151048
rect 306708 151036 306714 151088
rect 279510 150560 279516 150612
rect 279568 150600 279574 150612
rect 307570 150600 307576 150612
rect 279568 150572 307576 150600
rect 279568 150560 279574 150572
rect 307570 150560 307576 150572
rect 307628 150560 307634 150612
rect 208486 150492 208492 150544
rect 208544 150532 208550 150544
rect 214006 150532 214012 150544
rect 208544 150504 214012 150532
rect 208544 150492 208550 150504
rect 214006 150492 214012 150504
rect 214064 150492 214070 150544
rect 298922 150492 298928 150544
rect 298980 150532 298986 150544
rect 307662 150532 307668 150544
rect 298980 150504 307668 150532
rect 298980 150492 298986 150504
rect 307662 150492 307668 150504
rect 307720 150492 307726 150544
rect 205082 150424 205088 150476
rect 205140 150464 205146 150476
rect 213914 150464 213920 150476
rect 205140 150436 213920 150464
rect 205140 150424 205146 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 360838 150424 360844 150476
rect 360896 150464 360902 150476
rect 416774 150464 416780 150476
rect 360896 150436 416780 150464
rect 360896 150424 360902 150436
rect 416774 150424 416780 150436
rect 416832 150424 416838 150476
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 25498 150396 25504 150408
rect 3476 150368 25504 150396
rect 3476 150356 3482 150368
rect 25498 150356 25504 150368
rect 25556 150356 25562 150408
rect 170490 150356 170496 150408
rect 170548 150396 170554 150408
rect 214006 150396 214012 150408
rect 170548 150368 214012 150396
rect 170548 150356 170554 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 252462 150356 252468 150408
rect 252520 150396 252526 150408
rect 278774 150396 278780 150408
rect 252520 150368 278780 150396
rect 252520 150356 252526 150368
rect 278774 150356 278780 150368
rect 278832 150356 278838 150408
rect 324314 150356 324320 150408
rect 324372 150396 324378 150408
rect 345290 150396 345296 150408
rect 324372 150368 345296 150396
rect 324372 150356 324378 150368
rect 345290 150356 345296 150368
rect 345348 150356 345354 150408
rect 496814 150356 496820 150408
rect 496872 150396 496878 150408
rect 503898 150396 503904 150408
rect 496872 150368 503904 150396
rect 496872 150356 496878 150368
rect 503898 150356 503904 150368
rect 503956 150356 503962 150408
rect 208394 150288 208400 150340
rect 208452 150328 208458 150340
rect 213914 150328 213920 150340
rect 208452 150300 213920 150328
rect 208452 150288 208458 150300
rect 213914 150288 213920 150300
rect 213972 150288 213978 150340
rect 251358 150288 251364 150340
rect 251416 150328 251422 150340
rect 254026 150328 254032 150340
rect 251416 150300 254032 150328
rect 251416 150288 251422 150300
rect 254026 150288 254032 150300
rect 254084 150288 254090 150340
rect 324406 150288 324412 150340
rect 324464 150328 324470 150340
rect 331398 150328 331404 150340
rect 324464 150300 331404 150328
rect 324464 150288 324470 150300
rect 331398 150288 331404 150300
rect 331456 150288 331462 150340
rect 324590 149676 324596 149728
rect 324648 149716 324654 149728
rect 343818 149716 343824 149728
rect 324648 149688 343824 149716
rect 324648 149676 324654 149688
rect 343818 149676 343824 149688
rect 343876 149676 343882 149728
rect 304258 149200 304264 149252
rect 304316 149240 304322 149252
rect 307662 149240 307668 149252
rect 304316 149212 307668 149240
rect 304316 149200 304322 149212
rect 307662 149200 307668 149212
rect 307720 149200 307726 149252
rect 283650 149132 283656 149184
rect 283708 149172 283714 149184
rect 306742 149172 306748 149184
rect 283708 149144 306748 149172
rect 283708 149132 283714 149144
rect 306742 149132 306748 149144
rect 306800 149132 306806 149184
rect 254854 149064 254860 149116
rect 254912 149104 254918 149116
rect 307570 149104 307576 149116
rect 254912 149076 307576 149104
rect 254912 149064 254918 149076
rect 307570 149064 307576 149076
rect 307628 149064 307634 149116
rect 363598 149064 363604 149116
rect 363656 149104 363662 149116
rect 416774 149104 416780 149116
rect 363656 149076 416780 149104
rect 363656 149064 363662 149076
rect 416774 149064 416780 149076
rect 416832 149064 416838 149116
rect 252462 148996 252468 149048
rect 252520 149036 252526 149048
rect 272058 149036 272064 149048
rect 252520 149008 272064 149036
rect 252520 148996 252526 149008
rect 272058 148996 272064 149008
rect 272116 148996 272122 149048
rect 324406 148996 324412 149048
rect 324464 149036 324470 149048
rect 335538 149036 335544 149048
rect 324464 149008 335544 149036
rect 324464 148996 324470 149008
rect 335538 148996 335544 149008
rect 335596 148996 335602 149048
rect 252370 148928 252376 148980
rect 252428 148968 252434 148980
rect 256970 148968 256976 148980
rect 252428 148940 256976 148968
rect 252428 148928 252434 148940
rect 256970 148928 256976 148940
rect 257028 148928 257034 148980
rect 324314 148928 324320 148980
rect 324372 148968 324378 148980
rect 328638 148968 328644 148980
rect 324372 148940 328644 148968
rect 324372 148928 324378 148940
rect 328638 148928 328644 148940
rect 328696 148928 328702 148980
rect 289262 147772 289268 147824
rect 289320 147812 289326 147824
rect 306926 147812 306932 147824
rect 289320 147784 306932 147812
rect 289320 147772 289326 147784
rect 306926 147772 306932 147784
rect 306984 147772 306990 147824
rect 265618 147704 265624 147756
rect 265676 147744 265682 147756
rect 307570 147744 307576 147756
rect 265676 147716 307576 147744
rect 265676 147704 265682 147716
rect 307570 147704 307576 147716
rect 307628 147704 307634 147756
rect 254762 147636 254768 147688
rect 254820 147676 254826 147688
rect 307662 147676 307668 147688
rect 254820 147648 307668 147676
rect 254820 147636 254826 147648
rect 307662 147636 307668 147648
rect 307720 147636 307726 147688
rect 332502 147636 332508 147688
rect 332560 147676 332566 147688
rect 416774 147676 416780 147688
rect 332560 147648 416780 147676
rect 332560 147636 332566 147648
rect 416774 147636 416780 147648
rect 416832 147636 416838 147688
rect 252462 147568 252468 147620
rect 252520 147608 252526 147620
rect 270586 147608 270592 147620
rect 252520 147580 270592 147608
rect 252520 147568 252526 147580
rect 270586 147568 270592 147580
rect 270644 147568 270650 147620
rect 324314 147568 324320 147620
rect 324372 147608 324378 147620
rect 340874 147608 340880 147620
rect 324372 147580 340880 147608
rect 324372 147568 324378 147580
rect 340874 147568 340880 147580
rect 340932 147568 340938 147620
rect 496814 147568 496820 147620
rect 496872 147608 496878 147620
rect 505186 147608 505192 147620
rect 496872 147580 505192 147608
rect 496872 147568 496878 147580
rect 505186 147568 505192 147580
rect 505244 147568 505250 147620
rect 251358 147500 251364 147552
rect 251416 147540 251422 147552
rect 253934 147540 253940 147552
rect 251416 147512 253940 147540
rect 251416 147500 251422 147512
rect 253934 147500 253940 147512
rect 253992 147500 253998 147552
rect 252094 147432 252100 147484
rect 252152 147472 252158 147484
rect 255498 147472 255504 147484
rect 252152 147444 255504 147472
rect 252152 147432 252158 147444
rect 255498 147432 255504 147444
rect 255556 147432 255562 147484
rect 285122 146412 285128 146464
rect 285180 146452 285186 146464
rect 307570 146452 307576 146464
rect 285180 146424 307576 146452
rect 285180 146412 285186 146424
rect 307570 146412 307576 146424
rect 307628 146412 307634 146464
rect 200850 146344 200856 146396
rect 200908 146384 200914 146396
rect 213914 146384 213920 146396
rect 200908 146356 213920 146384
rect 200908 146344 200914 146356
rect 213914 146344 213920 146356
rect 213972 146344 213978 146396
rect 272610 146344 272616 146396
rect 272668 146384 272674 146396
rect 307662 146384 307668 146396
rect 272668 146356 307668 146384
rect 272668 146344 272674 146356
rect 307662 146344 307668 146356
rect 307720 146344 307726 146396
rect 171778 146276 171784 146328
rect 171836 146316 171842 146328
rect 214006 146316 214012 146328
rect 171836 146288 214012 146316
rect 171836 146276 171842 146288
rect 214006 146276 214012 146288
rect 214064 146276 214070 146328
rect 257522 146276 257528 146328
rect 257580 146316 257586 146328
rect 306742 146316 306748 146328
rect 257580 146288 306748 146316
rect 257580 146276 257586 146288
rect 306742 146276 306748 146288
rect 306800 146276 306806 146328
rect 345658 146276 345664 146328
rect 345716 146316 345722 146328
rect 416774 146316 416780 146328
rect 345716 146288 416780 146316
rect 345716 146276 345722 146288
rect 416774 146276 416780 146288
rect 416832 146276 416838 146328
rect 252370 146208 252376 146260
rect 252428 146248 252434 146260
rect 267734 146248 267740 146260
rect 252428 146220 267740 146248
rect 252428 146208 252434 146220
rect 267734 146208 267740 146220
rect 267792 146208 267798 146260
rect 324314 146208 324320 146260
rect 324372 146248 324378 146260
rect 356054 146248 356060 146260
rect 324372 146220 356060 146248
rect 324372 146208 324378 146220
rect 356054 146208 356060 146220
rect 356112 146208 356118 146260
rect 496814 146208 496820 146260
rect 496872 146248 496878 146260
rect 510798 146248 510804 146260
rect 496872 146220 510804 146248
rect 496872 146208 496878 146220
rect 510798 146208 510804 146220
rect 510856 146208 510862 146260
rect 252462 146140 252468 146192
rect 252520 146180 252526 146192
rect 260834 146180 260840 146192
rect 252520 146152 260840 146180
rect 252520 146140 252526 146152
rect 260834 146140 260840 146152
rect 260892 146140 260898 146192
rect 180242 145528 180248 145580
rect 180300 145568 180306 145580
rect 215018 145568 215024 145580
rect 180300 145540 215024 145568
rect 180300 145528 180306 145540
rect 215018 145528 215024 145540
rect 215076 145528 215082 145580
rect 277026 145528 277032 145580
rect 277084 145568 277090 145580
rect 307110 145568 307116 145580
rect 277084 145540 307116 145568
rect 277084 145528 277090 145540
rect 307110 145528 307116 145540
rect 307168 145528 307174 145580
rect 324406 145528 324412 145580
rect 324464 145568 324470 145580
rect 338298 145568 338304 145580
rect 324464 145540 338304 145568
rect 324464 145528 324470 145540
rect 338298 145528 338304 145540
rect 338356 145528 338362 145580
rect 166258 144916 166264 144968
rect 166316 144956 166322 144968
rect 213914 144956 213920 144968
rect 166316 144928 213920 144956
rect 166316 144916 166322 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 256142 144916 256148 144968
rect 256200 144956 256206 144968
rect 307662 144956 307668 144968
rect 256200 144928 307668 144956
rect 256200 144916 256206 144928
rect 307662 144916 307668 144928
rect 307720 144916 307726 144968
rect 252370 144848 252376 144900
rect 252428 144888 252434 144900
rect 269114 144888 269120 144900
rect 252428 144860 269120 144888
rect 252428 144848 252434 144860
rect 269114 144848 269120 144860
rect 269172 144848 269178 144900
rect 324314 144848 324320 144900
rect 324372 144888 324378 144900
rect 345198 144888 345204 144900
rect 324372 144860 345204 144888
rect 324372 144848 324378 144860
rect 345198 144848 345204 144860
rect 345256 144848 345262 144900
rect 252462 144780 252468 144832
rect 252520 144820 252526 144832
rect 262214 144820 262220 144832
rect 252520 144792 262220 144820
rect 252520 144780 252526 144792
rect 262214 144780 262220 144792
rect 262272 144780 262278 144832
rect 506566 144440 506572 144492
rect 506624 144480 506630 144492
rect 507118 144480 507124 144492
rect 506624 144452 507124 144480
rect 506624 144440 506630 144452
rect 507118 144440 507124 144452
rect 507176 144440 507182 144492
rect 167730 144168 167736 144220
rect 167788 144208 167794 144220
rect 208486 144208 208492 144220
rect 167788 144180 208492 144208
rect 167788 144168 167794 144180
rect 208486 144168 208492 144180
rect 208544 144168 208550 144220
rect 276934 144168 276940 144220
rect 276992 144208 276998 144220
rect 307570 144208 307576 144220
rect 276992 144180 307576 144208
rect 276992 144168 276998 144180
rect 307570 144168 307576 144180
rect 307628 144168 307634 144220
rect 496814 144168 496820 144220
rect 496872 144208 496878 144220
rect 506566 144208 506572 144220
rect 496872 144180 506572 144208
rect 496872 144168 496878 144180
rect 506566 144168 506572 144180
rect 506624 144168 506630 144220
rect 206462 143624 206468 143676
rect 206520 143664 206526 143676
rect 213914 143664 213920 143676
rect 206520 143636 213920 143664
rect 206520 143624 206526 143636
rect 213914 143624 213920 143636
rect 213972 143624 213978 143676
rect 251910 143624 251916 143676
rect 251968 143664 251974 143676
rect 260098 143664 260104 143676
rect 251968 143636 260104 143664
rect 251968 143624 251974 143636
rect 260098 143624 260104 143636
rect 260156 143624 260162 143676
rect 260190 143624 260196 143676
rect 260248 143664 260254 143676
rect 307662 143664 307668 143676
rect 260248 143636 307668 143664
rect 260248 143624 260254 143636
rect 307662 143624 307668 143636
rect 307720 143624 307726 143676
rect 198090 143556 198096 143608
rect 198148 143596 198154 143608
rect 214006 143596 214012 143608
rect 198148 143568 214012 143596
rect 198148 143556 198154 143568
rect 214006 143556 214012 143568
rect 214064 143556 214070 143608
rect 256050 143556 256056 143608
rect 256108 143596 256114 143608
rect 306926 143596 306932 143608
rect 256108 143568 306932 143596
rect 256108 143556 256114 143568
rect 306926 143556 306932 143568
rect 306984 143556 306990 143608
rect 352650 143556 352656 143608
rect 352708 143596 352714 143608
rect 416774 143596 416780 143608
rect 352708 143568 416780 143596
rect 352708 143556 352714 143568
rect 416774 143556 416780 143568
rect 416832 143556 416838 143608
rect 252462 143488 252468 143540
rect 252520 143528 252526 143540
rect 266354 143528 266360 143540
rect 252520 143500 266360 143528
rect 252520 143488 252526 143500
rect 266354 143488 266360 143500
rect 266412 143488 266418 143540
rect 324314 143488 324320 143540
rect 324372 143528 324378 143540
rect 328546 143528 328552 143540
rect 324372 143500 328552 143528
rect 324372 143488 324378 143500
rect 328546 143488 328552 143500
rect 328604 143488 328610 143540
rect 496814 143488 496820 143540
rect 496872 143528 496878 143540
rect 510706 143528 510712 143540
rect 496872 143500 510712 143528
rect 496872 143488 496878 143500
rect 510706 143488 510712 143500
rect 510764 143528 510770 143540
rect 512638 143528 512644 143540
rect 510764 143500 512644 143528
rect 510764 143488 510770 143500
rect 512638 143488 512644 143500
rect 512696 143488 512702 143540
rect 252370 143420 252376 143472
rect 252428 143460 252434 143472
rect 266446 143460 266452 143472
rect 252428 143432 266452 143460
rect 252428 143420 252434 143432
rect 266446 143420 266452 143432
rect 266504 143420 266510 143472
rect 253290 142808 253296 142860
rect 253348 142848 253354 142860
rect 307570 142848 307576 142860
rect 253348 142820 307576 142848
rect 253348 142808 253354 142820
rect 307570 142808 307576 142820
rect 307628 142808 307634 142860
rect 209222 142196 209228 142248
rect 209280 142236 209286 142248
rect 213914 142236 213920 142248
rect 209280 142208 213920 142236
rect 209280 142196 209286 142208
rect 213914 142196 213920 142208
rect 213972 142196 213978 142248
rect 269758 142196 269764 142248
rect 269816 142236 269822 142248
rect 307662 142236 307668 142248
rect 269816 142208 307668 142236
rect 269816 142196 269822 142208
rect 307662 142196 307668 142208
rect 307720 142196 307726 142248
rect 167638 142128 167644 142180
rect 167696 142168 167702 142180
rect 214006 142168 214012 142180
rect 167696 142140 214012 142168
rect 167696 142128 167702 142140
rect 214006 142128 214012 142140
rect 214064 142128 214070 142180
rect 256234 142128 256240 142180
rect 256292 142168 256298 142180
rect 306558 142168 306564 142180
rect 256292 142140 306564 142168
rect 256292 142128 256298 142140
rect 306558 142128 306564 142140
rect 306616 142128 306622 142180
rect 333238 142128 333244 142180
rect 333296 142168 333302 142180
rect 416866 142168 416872 142180
rect 333296 142140 416872 142168
rect 333296 142128 333302 142140
rect 416866 142128 416872 142140
rect 416924 142128 416930 142180
rect 324406 142060 324412 142112
rect 324464 142100 324470 142112
rect 343634 142100 343640 142112
rect 324464 142072 343640 142100
rect 324464 142060 324470 142072
rect 343634 142060 343640 142072
rect 343692 142060 343698 142112
rect 353294 142060 353300 142112
rect 353352 142100 353358 142112
rect 416774 142100 416780 142112
rect 353352 142072 416780 142100
rect 353352 142060 353358 142072
rect 416774 142060 416780 142072
rect 416832 142060 416838 142112
rect 324314 141992 324320 142044
rect 324372 142032 324378 142044
rect 329834 142032 329840 142044
rect 324372 142004 329840 142032
rect 324372 141992 324378 142004
rect 329834 141992 329840 142004
rect 329892 141992 329898 142044
rect 252186 141448 252192 141500
rect 252244 141488 252250 141500
rect 265802 141488 265808 141500
rect 252244 141460 265808 141488
rect 252244 141448 252250 141460
rect 265802 141448 265808 141460
rect 265860 141448 265866 141500
rect 253566 141380 253572 141432
rect 253624 141420 253630 141432
rect 307018 141420 307024 141432
rect 253624 141392 307024 141420
rect 253624 141380 253630 141392
rect 307018 141380 307024 141392
rect 307076 141380 307082 141432
rect 334618 141380 334624 141432
rect 334676 141420 334682 141432
rect 353294 141420 353300 141432
rect 334676 141392 353300 141420
rect 334676 141380 334682 141392
rect 353294 141380 353300 141392
rect 353352 141380 353358 141432
rect 304350 140904 304356 140956
rect 304408 140944 304414 140956
rect 307478 140944 307484 140956
rect 304408 140916 307484 140944
rect 304408 140904 304414 140916
rect 307478 140904 307484 140916
rect 307536 140904 307542 140956
rect 204990 140836 204996 140888
rect 205048 140876 205054 140888
rect 214006 140876 214012 140888
rect 205048 140848 214012 140876
rect 205048 140836 205054 140848
rect 214006 140836 214012 140848
rect 214064 140836 214070 140888
rect 286502 140836 286508 140888
rect 286560 140876 286566 140888
rect 306558 140876 306564 140888
rect 286560 140848 306564 140876
rect 286560 140836 286566 140848
rect 306558 140836 306564 140848
rect 306616 140836 306622 140888
rect 496814 140836 496820 140888
rect 496872 140876 496878 140888
rect 520182 140876 520188 140888
rect 496872 140848 520188 140876
rect 496872 140836 496878 140848
rect 520182 140836 520188 140848
rect 520240 140876 520246 140888
rect 521654 140876 521660 140888
rect 520240 140848 521660 140876
rect 520240 140836 520246 140848
rect 521654 140836 521660 140848
rect 521712 140836 521718 140888
rect 178770 140768 178776 140820
rect 178828 140808 178834 140820
rect 213914 140808 213920 140820
rect 178828 140780 213920 140808
rect 178828 140768 178834 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 267090 140768 267096 140820
rect 267148 140808 267154 140820
rect 307662 140808 307668 140820
rect 267148 140780 307668 140808
rect 267148 140768 267154 140780
rect 307662 140768 307668 140780
rect 307720 140768 307726 140820
rect 495342 140768 495348 140820
rect 495400 140808 495406 140820
rect 502794 140808 502800 140820
rect 495400 140780 502800 140808
rect 495400 140768 495406 140780
rect 502794 140768 502800 140780
rect 502852 140768 502858 140820
rect 252462 140700 252468 140752
rect 252520 140740 252526 140752
rect 273254 140740 273260 140752
rect 252520 140712 273260 140740
rect 252520 140700 252526 140712
rect 273254 140700 273260 140712
rect 273312 140700 273318 140752
rect 496814 140700 496820 140752
rect 496872 140740 496878 140752
rect 502518 140740 502524 140752
rect 496872 140712 502524 140740
rect 496872 140700 496878 140712
rect 502518 140700 502524 140712
rect 502576 140700 502582 140752
rect 174630 140020 174636 140072
rect 174688 140060 174694 140072
rect 214742 140060 214748 140072
rect 174688 140032 214748 140060
rect 174688 140020 174694 140032
rect 214742 140020 214748 140032
rect 214800 140020 214806 140072
rect 502794 140020 502800 140072
rect 502852 140060 502858 140072
rect 580166 140060 580172 140072
rect 502852 140032 580172 140060
rect 502852 140020 502858 140032
rect 580166 140020 580172 140032
rect 580224 140020 580230 140072
rect 264238 139544 264244 139596
rect 264296 139584 264302 139596
rect 307662 139584 307668 139596
rect 264296 139556 307668 139584
rect 264296 139544 264302 139556
rect 307662 139544 307668 139556
rect 307720 139544 307726 139596
rect 211890 139476 211896 139528
rect 211948 139516 211954 139528
rect 214650 139516 214656 139528
rect 211948 139488 214656 139516
rect 211948 139476 211954 139488
rect 214650 139476 214656 139488
rect 214708 139476 214714 139528
rect 262950 139476 262956 139528
rect 263008 139516 263014 139528
rect 307570 139516 307576 139528
rect 263008 139488 307576 139516
rect 263008 139476 263014 139488
rect 307570 139476 307576 139488
rect 307628 139476 307634 139528
rect 166350 139408 166356 139460
rect 166408 139448 166414 139460
rect 213914 139448 213920 139460
rect 166408 139420 213920 139448
rect 166408 139408 166414 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 250622 139408 250628 139460
rect 250680 139448 250686 139460
rect 307294 139448 307300 139460
rect 250680 139420 307300 139448
rect 250680 139408 250686 139420
rect 307294 139408 307300 139420
rect 307352 139408 307358 139460
rect 367830 139408 367836 139460
rect 367888 139448 367894 139460
rect 416774 139448 416780 139460
rect 367888 139420 416780 139448
rect 367888 139408 367894 139420
rect 416774 139408 416780 139420
rect 416832 139408 416838 139460
rect 252462 139340 252468 139392
rect 252520 139380 252526 139392
rect 280154 139380 280160 139392
rect 252520 139352 280160 139380
rect 252520 139340 252526 139352
rect 280154 139340 280160 139352
rect 280212 139340 280218 139392
rect 324314 139340 324320 139392
rect 324372 139380 324378 139392
rect 346578 139380 346584 139392
rect 324372 139352 346584 139380
rect 324372 139340 324378 139352
rect 346578 139340 346584 139352
rect 346636 139340 346642 139392
rect 496814 139340 496820 139392
rect 496872 139380 496878 139392
rect 520918 139380 520924 139392
rect 496872 139352 520924 139380
rect 496872 139340 496878 139352
rect 520918 139340 520924 139352
rect 520976 139340 520982 139392
rect 287790 138116 287796 138168
rect 287848 138156 287854 138168
rect 307294 138156 307300 138168
rect 287848 138128 307300 138156
rect 287848 138116 287854 138128
rect 307294 138116 307300 138128
rect 307352 138116 307358 138168
rect 253198 138048 253204 138100
rect 253256 138088 253262 138100
rect 306558 138088 306564 138100
rect 253256 138060 306564 138088
rect 253256 138048 253262 138060
rect 306558 138048 306564 138060
rect 306616 138048 306622 138100
rect 170398 137980 170404 138032
rect 170456 138020 170462 138032
rect 213914 138020 213920 138032
rect 170456 137992 213920 138020
rect 170456 137980 170462 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 250530 137980 250536 138032
rect 250588 138020 250594 138032
rect 307662 138020 307668 138032
rect 250588 137992 307668 138020
rect 250588 137980 250594 137992
rect 307662 137980 307668 137992
rect 307720 137980 307726 138032
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 15838 137952 15844 137964
rect 3292 137924 15844 137952
rect 3292 137912 3298 137924
rect 15838 137912 15844 137924
rect 15896 137912 15902 137964
rect 252462 137912 252468 137964
rect 252520 137952 252526 137964
rect 274634 137952 274640 137964
rect 252520 137924 274640 137952
rect 252520 137912 252526 137924
rect 274634 137912 274640 137924
rect 274692 137912 274698 137964
rect 324406 137912 324412 137964
rect 324464 137952 324470 137964
rect 339586 137952 339592 137964
rect 324464 137924 339592 137952
rect 324464 137912 324470 137924
rect 339586 137912 339592 137924
rect 339644 137912 339650 137964
rect 358814 137912 358820 137964
rect 358872 137952 358878 137964
rect 416774 137952 416780 137964
rect 358872 137924 416780 137952
rect 358872 137912 358878 137924
rect 416774 137912 416780 137924
rect 416832 137912 416838 137964
rect 496814 137912 496820 137964
rect 496872 137952 496878 137964
rect 548518 137952 548524 137964
rect 496872 137924 548524 137952
rect 496872 137912 496878 137924
rect 548518 137912 548524 137924
rect 548576 137912 548582 137964
rect 324314 137844 324320 137896
rect 324372 137884 324378 137896
rect 336918 137884 336924 137896
rect 324372 137856 336924 137884
rect 324372 137844 324378 137856
rect 336918 137844 336924 137856
rect 336976 137844 336982 137896
rect 290458 137232 290464 137284
rect 290516 137272 290522 137284
rect 307202 137272 307208 137284
rect 290516 137244 307208 137272
rect 290516 137232 290522 137244
rect 307202 137232 307208 137244
rect 307260 137232 307266 137284
rect 354030 137232 354036 137284
rect 354088 137272 354094 137284
rect 358814 137272 358820 137284
rect 354088 137244 358820 137272
rect 354088 137232 354094 137244
rect 358814 137232 358820 137244
rect 358872 137232 358878 137284
rect 202414 136688 202420 136740
rect 202472 136728 202478 136740
rect 213914 136728 213920 136740
rect 202472 136700 213920 136728
rect 202472 136688 202478 136700
rect 213914 136688 213920 136700
rect 213972 136688 213978 136740
rect 181530 136620 181536 136672
rect 181588 136660 181594 136672
rect 214006 136660 214012 136672
rect 181588 136632 214012 136660
rect 181588 136620 181594 136632
rect 214006 136620 214012 136632
rect 214064 136620 214070 136672
rect 250438 136620 250444 136672
rect 250496 136660 250502 136672
rect 307662 136660 307668 136672
rect 250496 136632 307668 136660
rect 250496 136620 250502 136632
rect 307662 136620 307668 136632
rect 307720 136620 307726 136672
rect 252278 136552 252284 136604
rect 252336 136592 252342 136604
rect 284938 136592 284944 136604
rect 252336 136564 284944 136592
rect 252336 136552 252342 136564
rect 284938 136552 284944 136564
rect 284996 136552 285002 136604
rect 324406 136552 324412 136604
rect 324464 136592 324470 136604
rect 351914 136592 351920 136604
rect 324464 136564 351920 136592
rect 324464 136552 324470 136564
rect 351914 136552 351920 136564
rect 351972 136552 351978 136604
rect 496906 136552 496912 136604
rect 496964 136592 496970 136604
rect 508498 136592 508504 136604
rect 496964 136564 508504 136592
rect 496964 136552 496970 136564
rect 508498 136552 508504 136564
rect 508556 136552 508562 136604
rect 252462 136484 252468 136536
rect 252520 136524 252526 136536
rect 271874 136524 271880 136536
rect 252520 136496 271880 136524
rect 252520 136484 252526 136496
rect 271874 136484 271880 136496
rect 271932 136484 271938 136536
rect 324314 136484 324320 136536
rect 324372 136524 324378 136536
rect 338206 136524 338212 136536
rect 324372 136496 338212 136524
rect 324372 136484 324378 136496
rect 338206 136484 338212 136496
rect 338264 136484 338270 136536
rect 252370 136416 252376 136468
rect 252428 136456 252434 136468
rect 263042 136456 263048 136468
rect 252428 136428 263048 136456
rect 252428 136416 252434 136428
rect 263042 136416 263048 136428
rect 263100 136416 263106 136468
rect 496814 136348 496820 136400
rect 496872 136388 496878 136400
rect 501230 136388 501236 136400
rect 496872 136360 501236 136388
rect 496872 136348 496878 136360
rect 501230 136348 501236 136360
rect 501288 136348 501294 136400
rect 300118 135464 300124 135516
rect 300176 135504 300182 135516
rect 307662 135504 307668 135516
rect 300176 135476 307668 135504
rect 300176 135464 300182 135476
rect 307662 135464 307668 135476
rect 307720 135464 307726 135516
rect 289170 135396 289176 135448
rect 289228 135436 289234 135448
rect 307294 135436 307300 135448
rect 289228 135408 307300 135436
rect 289228 135396 289234 135408
rect 307294 135396 307300 135408
rect 307352 135396 307358 135448
rect 280982 135328 280988 135380
rect 281040 135368 281046 135380
rect 307570 135368 307576 135380
rect 281040 135340 307576 135368
rect 281040 135328 281046 135340
rect 307570 135328 307576 135340
rect 307628 135328 307634 135380
rect 196710 135260 196716 135312
rect 196768 135300 196774 135312
rect 213914 135300 213920 135312
rect 196768 135272 213920 135300
rect 196768 135260 196774 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 254670 135260 254676 135312
rect 254728 135300 254734 135312
rect 306558 135300 306564 135312
rect 254728 135272 306564 135300
rect 254728 135260 254734 135272
rect 306558 135260 306564 135272
rect 306616 135260 306622 135312
rect 370498 135260 370504 135312
rect 370556 135300 370562 135312
rect 416774 135300 416780 135312
rect 370556 135272 416780 135300
rect 370556 135260 370562 135272
rect 416774 135260 416780 135272
rect 416832 135260 416838 135312
rect 252370 135192 252376 135244
rect 252428 135232 252434 135244
rect 302878 135232 302884 135244
rect 252428 135204 302884 135232
rect 252428 135192 252434 135204
rect 302878 135192 302884 135204
rect 302936 135192 302942 135244
rect 334710 135192 334716 135244
rect 334768 135232 334774 135244
rect 417326 135232 417332 135244
rect 334768 135204 417332 135232
rect 334768 135192 334774 135204
rect 417326 135192 417332 135204
rect 417384 135192 417390 135244
rect 252462 135124 252468 135176
rect 252520 135164 252526 135176
rect 276750 135164 276756 135176
rect 252520 135136 276756 135164
rect 252520 135124 252526 135136
rect 276750 135124 276756 135136
rect 276808 135124 276814 135176
rect 265802 134512 265808 134564
rect 265860 134552 265866 134564
rect 307386 134552 307392 134564
rect 265860 134524 307392 134552
rect 265860 134512 265866 134524
rect 307386 134512 307392 134524
rect 307444 134512 307450 134564
rect 198274 133968 198280 134020
rect 198332 134008 198338 134020
rect 214006 134008 214012 134020
rect 198332 133980 214012 134008
rect 198332 133968 198338 133980
rect 214006 133968 214012 133980
rect 214064 133968 214070 134020
rect 177390 133900 177396 133952
rect 177448 133940 177454 133952
rect 213914 133940 213920 133952
rect 177448 133912 213920 133940
rect 177448 133900 177454 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 286410 133900 286416 133952
rect 286468 133940 286474 133952
rect 306558 133940 306564 133952
rect 286468 133912 306564 133940
rect 286468 133900 286474 133912
rect 306558 133900 306564 133912
rect 306616 133900 306622 133952
rect 252462 133832 252468 133884
rect 252520 133872 252526 133884
rect 298738 133872 298744 133884
rect 252520 133844 298744 133872
rect 252520 133832 252526 133844
rect 298738 133832 298744 133844
rect 298796 133832 298802 133884
rect 374638 133832 374644 133884
rect 374696 133872 374702 133884
rect 419442 133872 419448 133884
rect 374696 133844 419448 133872
rect 374696 133832 374702 133844
rect 419442 133832 419448 133844
rect 419500 133832 419506 133884
rect 496814 133832 496820 133884
rect 496872 133872 496878 133884
rect 511994 133872 512000 133884
rect 496872 133844 512000 133872
rect 496872 133832 496878 133844
rect 511994 133832 512000 133844
rect 512052 133832 512058 133884
rect 252278 133764 252284 133816
rect 252336 133804 252342 133816
rect 295978 133804 295984 133816
rect 252336 133776 295984 133804
rect 252336 133764 252342 133776
rect 295978 133764 295984 133776
rect 296036 133764 296042 133816
rect 252370 133696 252376 133748
rect 252428 133736 252434 133748
rect 265710 133736 265716 133748
rect 252428 133708 265716 133736
rect 252428 133696 252434 133708
rect 265710 133696 265716 133708
rect 265768 133696 265774 133748
rect 404262 133152 404268 133204
rect 404320 133192 404326 133204
rect 419626 133192 419632 133204
rect 404320 133164 419632 133192
rect 404320 133152 404326 133164
rect 419626 133152 419632 133164
rect 419684 133152 419690 133204
rect 210510 132880 210516 132932
rect 210568 132920 210574 132932
rect 213914 132920 213920 132932
rect 210568 132892 213920 132920
rect 210568 132880 210574 132892
rect 213914 132880 213920 132892
rect 213972 132880 213978 132932
rect 300210 132608 300216 132660
rect 300268 132648 300274 132660
rect 306926 132648 306932 132660
rect 300268 132620 306932 132648
rect 300268 132608 300274 132620
rect 306926 132608 306932 132620
rect 306984 132608 306990 132660
rect 297358 132540 297364 132592
rect 297416 132580 297422 132592
rect 307294 132580 307300 132592
rect 297416 132552 307300 132580
rect 297416 132540 297422 132552
rect 307294 132540 307300 132552
rect 307352 132540 307358 132592
rect 171962 132472 171968 132524
rect 172020 132512 172026 132524
rect 213914 132512 213920 132524
rect 172020 132484 213920 132512
rect 172020 132472 172026 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 292022 132472 292028 132524
rect 292080 132512 292086 132524
rect 306558 132512 306564 132524
rect 292080 132484 306564 132512
rect 292080 132472 292086 132484
rect 306558 132472 306564 132484
rect 306616 132472 306622 132524
rect 252278 132404 252284 132456
rect 252336 132444 252342 132456
rect 297450 132444 297456 132456
rect 252336 132416 297456 132444
rect 252336 132404 252342 132416
rect 297450 132404 297456 132416
rect 297508 132404 297514 132456
rect 367738 132404 367744 132456
rect 367796 132444 367802 132456
rect 417510 132444 417516 132456
rect 367796 132416 417516 132444
rect 367796 132404 367802 132416
rect 417510 132404 417516 132416
rect 417568 132404 417574 132456
rect 252462 132336 252468 132388
rect 252520 132376 252526 132388
rect 278222 132376 278228 132388
rect 252520 132348 278228 132376
rect 252520 132336 252526 132348
rect 278222 132336 278228 132348
rect 278280 132336 278286 132388
rect 252370 132268 252376 132320
rect 252428 132308 252434 132320
rect 264330 132308 264336 132320
rect 252428 132280 264336 132308
rect 252428 132268 252434 132280
rect 264330 132268 264336 132280
rect 264388 132268 264394 132320
rect 294598 131248 294604 131300
rect 294656 131288 294662 131300
rect 307478 131288 307484 131300
rect 294656 131260 307484 131288
rect 294656 131248 294662 131260
rect 307478 131248 307484 131260
rect 307536 131248 307542 131300
rect 290550 131180 290556 131232
rect 290608 131220 290614 131232
rect 307570 131220 307576 131232
rect 290608 131192 307576 131220
rect 290608 131180 290614 131192
rect 307570 131180 307576 131192
rect 307628 131180 307634 131232
rect 202322 131112 202328 131164
rect 202380 131152 202386 131164
rect 213914 131152 213920 131164
rect 202380 131124 213920 131152
rect 202380 131112 202386 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 278130 131112 278136 131164
rect 278188 131152 278194 131164
rect 307662 131152 307668 131164
rect 278188 131124 307668 131152
rect 278188 131112 278194 131124
rect 307662 131112 307668 131124
rect 307720 131112 307726 131164
rect 497458 131112 497464 131164
rect 497516 131152 497522 131164
rect 498286 131152 498292 131164
rect 497516 131124 498292 131152
rect 497516 131112 497522 131124
rect 498286 131112 498292 131124
rect 498344 131112 498350 131164
rect 252462 131044 252468 131096
rect 252520 131084 252526 131096
rect 267182 131084 267188 131096
rect 252520 131056 267188 131084
rect 252520 131044 252526 131056
rect 267182 131044 267188 131056
rect 267240 131044 267246 131096
rect 324406 131044 324412 131096
rect 324464 131084 324470 131096
rect 346486 131084 346492 131096
rect 324464 131056 346492 131084
rect 324464 131044 324470 131056
rect 346486 131044 346492 131056
rect 346544 131044 346550 131096
rect 252370 130976 252376 131028
rect 252428 131016 252434 131028
rect 261662 131016 261668 131028
rect 252428 130988 261668 131016
rect 252428 130976 252434 130988
rect 261662 130976 261668 130988
rect 261720 130976 261726 131028
rect 324314 130976 324320 131028
rect 324372 131016 324378 131028
rect 331306 131016 331312 131028
rect 324372 130988 331312 131016
rect 324372 130976 324378 130988
rect 331306 130976 331312 130988
rect 331364 130976 331370 131028
rect 252462 130160 252468 130212
rect 252520 130200 252526 130212
rect 258994 130200 259000 130212
rect 252520 130172 259000 130200
rect 252520 130160 252526 130172
rect 258994 130160 259000 130172
rect 259052 130160 259058 130212
rect 301498 129888 301504 129940
rect 301556 129928 301562 129940
rect 307478 129928 307484 129940
rect 301556 129900 307484 129928
rect 301556 129888 301562 129900
rect 307478 129888 307484 129900
rect 307536 129888 307542 129940
rect 176010 129820 176016 129872
rect 176068 129860 176074 129872
rect 213914 129860 213920 129872
rect 176068 129832 213920 129860
rect 176068 129820 176074 129832
rect 213914 129820 213920 129832
rect 213972 129820 213978 129872
rect 304442 129820 304448 129872
rect 304500 129860 304506 129872
rect 306926 129860 306932 129872
rect 304500 129832 306932 129860
rect 304500 129820 304506 129832
rect 306926 129820 306932 129832
rect 306984 129820 306990 129872
rect 173342 129752 173348 129804
rect 173400 129792 173406 129804
rect 214006 129792 214012 129804
rect 173400 129764 214012 129792
rect 173400 129752 173406 129764
rect 214006 129752 214012 129764
rect 214064 129752 214070 129804
rect 261570 129752 261576 129804
rect 261628 129792 261634 129804
rect 306558 129792 306564 129804
rect 261628 129764 306564 129792
rect 261628 129752 261634 129764
rect 306558 129752 306564 129764
rect 306616 129752 306622 129804
rect 252278 129684 252284 129736
rect 252336 129724 252342 129736
rect 300302 129724 300308 129736
rect 252336 129696 300308 129724
rect 252336 129684 252342 129696
rect 300302 129684 300308 129696
rect 300360 129684 300366 129736
rect 324314 129684 324320 129736
rect 324372 129724 324378 129736
rect 349338 129724 349344 129736
rect 324372 129696 349344 129724
rect 324372 129684 324378 129696
rect 349338 129684 349344 129696
rect 349396 129684 349402 129736
rect 496814 129684 496820 129736
rect 496872 129724 496878 129736
rect 509234 129724 509240 129736
rect 496872 129696 509240 129724
rect 496872 129684 496878 129696
rect 509234 129684 509240 129696
rect 509292 129684 509298 129736
rect 252462 129616 252468 129668
rect 252520 129656 252526 129668
rect 291930 129656 291936 129668
rect 252520 129628 291936 129656
rect 252520 129616 252526 129628
rect 291930 129616 291936 129628
rect 291988 129616 291994 129668
rect 252370 129548 252376 129600
rect 252428 129588 252434 129600
rect 264422 129588 264428 129600
rect 252428 129560 264428 129588
rect 252428 129548 252434 129560
rect 264422 129548 264428 129560
rect 264480 129548 264486 129600
rect 298830 128460 298836 128512
rect 298888 128500 298894 128512
rect 307662 128500 307668 128512
rect 298888 128472 307668 128500
rect 298888 128460 298894 128472
rect 307662 128460 307668 128472
rect 307720 128460 307726 128512
rect 284938 128392 284944 128444
rect 284996 128432 285002 128444
rect 306926 128432 306932 128444
rect 284996 128404 306932 128432
rect 284996 128392 285002 128404
rect 306926 128392 306932 128404
rect 306984 128392 306990 128444
rect 177482 128324 177488 128376
rect 177540 128364 177546 128376
rect 213914 128364 213920 128376
rect 177540 128336 213920 128364
rect 177540 128324 177546 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 264330 128324 264336 128376
rect 264388 128364 264394 128376
rect 307570 128364 307576 128376
rect 264388 128336 307576 128364
rect 264388 128324 264394 128336
rect 307570 128324 307576 128336
rect 307628 128324 307634 128376
rect 252370 128256 252376 128308
rect 252428 128296 252434 128308
rect 271138 128296 271144 128308
rect 252428 128268 271144 128296
rect 252428 128256 252434 128268
rect 271138 128256 271144 128268
rect 271196 128256 271202 128308
rect 324314 128256 324320 128308
rect 324372 128296 324378 128308
rect 350626 128296 350632 128308
rect 324372 128268 350632 128296
rect 324372 128256 324378 128268
rect 350626 128256 350632 128268
rect 350684 128256 350690 128308
rect 382918 128256 382924 128308
rect 382976 128296 382982 128308
rect 418706 128296 418712 128308
rect 382976 128268 418712 128296
rect 382976 128256 382982 128268
rect 418706 128256 418712 128268
rect 418764 128256 418770 128308
rect 496814 128256 496820 128308
rect 496872 128296 496878 128308
rect 507854 128296 507860 128308
rect 496872 128268 507860 128296
rect 496872 128256 496878 128268
rect 507854 128256 507860 128268
rect 507912 128256 507918 128308
rect 252462 128188 252468 128240
rect 252520 128228 252526 128240
rect 268378 128228 268384 128240
rect 252520 128200 268384 128228
rect 252520 128188 252526 128200
rect 268378 128188 268384 128200
rect 268436 128188 268442 128240
rect 324406 128188 324412 128240
rect 324464 128228 324470 128240
rect 329926 128228 329932 128240
rect 324464 128200 329932 128228
rect 324464 128188 324470 128200
rect 329926 128188 329932 128200
rect 329984 128188 329990 128240
rect 252278 128120 252284 128172
rect 252336 128160 252342 128172
rect 257614 128160 257620 128172
rect 252336 128132 257620 128160
rect 252336 128120 252342 128132
rect 257614 128120 257620 128132
rect 257672 128120 257678 128172
rect 268562 127644 268568 127696
rect 268620 127684 268626 127696
rect 307386 127684 307392 127696
rect 268620 127656 307392 127684
rect 268620 127644 268626 127656
rect 307386 127644 307392 127656
rect 307444 127644 307450 127696
rect 252186 127576 252192 127628
rect 252244 127616 252250 127628
rect 305638 127616 305644 127628
rect 252244 127588 305644 127616
rect 252244 127576 252250 127588
rect 305638 127576 305644 127588
rect 305696 127576 305702 127628
rect 530578 127576 530584 127628
rect 530636 127616 530642 127628
rect 580166 127616 580172 127628
rect 530636 127588 580172 127616
rect 530636 127576 530642 127588
rect 580166 127576 580172 127588
rect 580224 127576 580230 127628
rect 496906 127236 496912 127288
rect 496964 127276 496970 127288
rect 499850 127276 499856 127288
rect 496964 127248 499856 127276
rect 496964 127236 496970 127248
rect 499850 127236 499856 127248
rect 499908 127236 499914 127288
rect 184382 127032 184388 127084
rect 184440 127072 184446 127084
rect 214006 127072 214012 127084
rect 184440 127044 214012 127072
rect 184440 127032 184446 127044
rect 214006 127032 214012 127044
rect 214064 127032 214070 127084
rect 295978 127032 295984 127084
rect 296036 127072 296042 127084
rect 307570 127072 307576 127084
rect 296036 127044 307576 127072
rect 296036 127032 296042 127044
rect 307570 127032 307576 127044
rect 307628 127032 307634 127084
rect 57790 126964 57796 127016
rect 57848 127004 57854 127016
rect 65518 127004 65524 127016
rect 57848 126976 65524 127004
rect 57848 126964 57854 126976
rect 65518 126964 65524 126976
rect 65576 126964 65582 127016
rect 173250 126964 173256 127016
rect 173308 127004 173314 127016
rect 213914 127004 213920 127016
rect 173308 126976 213920 127004
rect 173308 126964 173314 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 293218 126964 293224 127016
rect 293276 127004 293282 127016
rect 307662 127004 307668 127016
rect 293276 126976 307668 127004
rect 293276 126964 293282 126976
rect 307662 126964 307668 126976
rect 307720 126964 307726 127016
rect 252462 126896 252468 126948
rect 252520 126936 252526 126948
rect 272518 126936 272524 126948
rect 252520 126908 272524 126936
rect 252520 126896 252526 126908
rect 272518 126896 272524 126908
rect 272576 126896 272582 126948
rect 496814 126896 496820 126948
rect 496872 126936 496878 126948
rect 514754 126936 514760 126948
rect 496872 126908 514760 126936
rect 496872 126896 496878 126908
rect 514754 126896 514760 126908
rect 514812 126896 514818 126948
rect 251174 126828 251180 126880
rect 251232 126868 251238 126880
rect 253382 126868 253388 126880
rect 251232 126840 253388 126868
rect 251232 126828 251238 126840
rect 253382 126828 253388 126840
rect 253440 126828 253446 126880
rect 252462 126420 252468 126472
rect 252520 126460 252526 126472
rect 258718 126460 258724 126472
rect 252520 126432 258724 126460
rect 252520 126420 252526 126432
rect 258718 126420 258724 126432
rect 258776 126420 258782 126472
rect 252278 126216 252284 126268
rect 252336 126256 252342 126268
rect 293310 126256 293316 126268
rect 252336 126228 293316 126256
rect 252336 126216 252342 126228
rect 293310 126216 293316 126228
rect 293368 126216 293374 126268
rect 296162 125740 296168 125792
rect 296220 125780 296226 125792
rect 307662 125780 307668 125792
rect 296220 125752 307668 125780
rect 296220 125740 296226 125752
rect 307662 125740 307668 125752
rect 307720 125740 307726 125792
rect 192478 125672 192484 125724
rect 192536 125712 192542 125724
rect 214006 125712 214012 125724
rect 192536 125684 214012 125712
rect 192536 125672 192542 125684
rect 214006 125672 214012 125684
rect 214064 125672 214070 125724
rect 283558 125672 283564 125724
rect 283616 125712 283622 125724
rect 307478 125712 307484 125724
rect 283616 125684 307484 125712
rect 283616 125672 283622 125684
rect 307478 125672 307484 125684
rect 307536 125672 307542 125724
rect 169110 125604 169116 125656
rect 169168 125644 169174 125656
rect 213914 125644 213920 125656
rect 169168 125616 213920 125644
rect 169168 125604 169174 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 275278 125604 275284 125656
rect 275336 125644 275342 125656
rect 307570 125644 307576 125656
rect 275336 125616 307576 125644
rect 275336 125604 275342 125616
rect 307570 125604 307576 125616
rect 307628 125604 307634 125656
rect 252094 125536 252100 125588
rect 252152 125576 252158 125588
rect 253566 125576 253572 125588
rect 252152 125548 253572 125576
rect 252152 125536 252158 125548
rect 253566 125536 253572 125548
rect 253624 125536 253630 125588
rect 324406 125536 324412 125588
rect 324464 125576 324470 125588
rect 346394 125576 346400 125588
rect 324464 125548 346400 125576
rect 324464 125536 324470 125548
rect 346394 125536 346400 125548
rect 346452 125536 346458 125588
rect 496814 125536 496820 125588
rect 496872 125576 496878 125588
rect 513374 125576 513380 125588
rect 496872 125548 513380 125576
rect 496872 125536 496878 125548
rect 513374 125536 513380 125548
rect 513432 125536 513438 125588
rect 252462 125468 252468 125520
rect 252520 125508 252526 125520
rect 269850 125508 269856 125520
rect 252520 125480 269856 125508
rect 252520 125468 252526 125480
rect 269850 125468 269856 125480
rect 269908 125468 269914 125520
rect 324314 125468 324320 125520
rect 324372 125508 324378 125520
rect 327718 125508 327724 125520
rect 324372 125480 327724 125508
rect 324372 125468 324378 125480
rect 327718 125468 327724 125480
rect 327776 125468 327782 125520
rect 252370 125400 252376 125452
rect 252428 125440 252434 125452
rect 301590 125440 301596 125452
rect 252428 125412 301596 125440
rect 252428 125400 252434 125412
rect 301590 125400 301596 125412
rect 301648 125400 301654 125452
rect 301682 124312 301688 124364
rect 301740 124352 301746 124364
rect 307662 124352 307668 124364
rect 301740 124324 307668 124352
rect 301740 124312 301746 124324
rect 307662 124312 307668 124324
rect 307720 124312 307726 124364
rect 180334 124244 180340 124296
rect 180392 124284 180398 124296
rect 213914 124284 213920 124296
rect 180392 124256 213920 124284
rect 180392 124244 180398 124256
rect 213914 124244 213920 124256
rect 213972 124244 213978 124296
rect 285030 124244 285036 124296
rect 285088 124284 285094 124296
rect 307570 124284 307576 124296
rect 285088 124256 307576 124284
rect 285088 124244 285094 124256
rect 307570 124244 307576 124256
rect 307628 124244 307634 124296
rect 171870 124176 171876 124228
rect 171928 124216 171934 124228
rect 214006 124216 214012 124228
rect 171928 124188 214012 124216
rect 171928 124176 171934 124188
rect 214006 124176 214012 124188
rect 214064 124176 214070 124228
rect 272518 124176 272524 124228
rect 272576 124216 272582 124228
rect 307478 124216 307484 124228
rect 272576 124188 307484 124216
rect 272576 124176 272582 124188
rect 307478 124176 307484 124188
rect 307536 124176 307542 124228
rect 252462 124108 252468 124160
rect 252520 124148 252526 124160
rect 302970 124148 302976 124160
rect 252520 124120 302976 124148
rect 252520 124108 252526 124120
rect 302970 124108 302976 124120
rect 303028 124108 303034 124160
rect 324406 124108 324412 124160
rect 324464 124148 324470 124160
rect 349246 124148 349252 124160
rect 324464 124120 349252 124148
rect 324464 124108 324470 124120
rect 349246 124108 349252 124120
rect 349304 124108 349310 124160
rect 324314 124040 324320 124092
rect 324372 124080 324378 124092
rect 347774 124080 347780 124092
rect 324372 124052 347780 124080
rect 324372 124040 324378 124052
rect 347774 124040 347780 124052
rect 347832 124040 347838 124092
rect 496814 124040 496820 124092
rect 496872 124080 496878 124092
rect 499574 124080 499580 124092
rect 496872 124052 499580 124080
rect 496872 124040 496878 124052
rect 499574 124040 499580 124052
rect 499632 124040 499638 124092
rect 251726 123428 251732 123480
rect 251784 123468 251790 123480
rect 264514 123468 264520 123480
rect 251784 123440 264520 123468
rect 251784 123428 251790 123440
rect 264514 123428 264520 123440
rect 264572 123428 264578 123480
rect 293310 122952 293316 123004
rect 293368 122992 293374 123004
rect 307570 122992 307576 123004
rect 293368 122964 307576 122992
rect 293368 122952 293374 122964
rect 307570 122952 307576 122964
rect 307628 122952 307634 123004
rect 196802 122884 196808 122936
rect 196860 122924 196866 122936
rect 213914 122924 213920 122936
rect 196860 122896 213920 122924
rect 196860 122884 196866 122896
rect 213914 122884 213920 122896
rect 213972 122884 213978 122936
rect 56502 122816 56508 122868
rect 56560 122856 56566 122868
rect 66070 122856 66076 122868
rect 56560 122828 66076 122856
rect 56560 122816 56566 122828
rect 66070 122816 66076 122828
rect 66128 122816 66134 122868
rect 170490 122816 170496 122868
rect 170548 122856 170554 122868
rect 214006 122856 214012 122868
rect 170548 122828 214012 122856
rect 170548 122816 170554 122828
rect 214006 122816 214012 122828
rect 214064 122816 214070 122868
rect 303062 122816 303068 122868
rect 303120 122856 303126 122868
rect 307662 122856 307668 122868
rect 303120 122828 307668 122856
rect 303120 122816 303126 122828
rect 307662 122816 307668 122828
rect 307720 122816 307726 122868
rect 252462 122748 252468 122800
rect 252520 122788 252526 122800
rect 299014 122788 299020 122800
rect 252520 122760 299020 122788
rect 252520 122748 252526 122760
rect 299014 122748 299020 122760
rect 299072 122748 299078 122800
rect 324314 122748 324320 122800
rect 324372 122788 324378 122800
rect 347958 122788 347964 122800
rect 324372 122760 347964 122788
rect 324372 122748 324378 122760
rect 347958 122748 347964 122760
rect 348016 122748 348022 122800
rect 376662 122748 376668 122800
rect 376720 122788 376726 122800
rect 416774 122788 416780 122800
rect 376720 122760 416780 122788
rect 376720 122748 376726 122760
rect 416774 122748 416780 122760
rect 416832 122748 416838 122800
rect 496814 122748 496820 122800
rect 496872 122788 496878 122800
rect 505094 122788 505100 122800
rect 496872 122760 505100 122788
rect 496872 122748 496878 122760
rect 505094 122748 505100 122760
rect 505152 122748 505158 122800
rect 252370 122680 252376 122732
rect 252428 122720 252434 122732
rect 269942 122720 269948 122732
rect 252428 122692 269948 122720
rect 252428 122680 252434 122692
rect 269942 122680 269948 122692
rect 270000 122680 270006 122732
rect 324406 122680 324412 122732
rect 324464 122720 324470 122732
rect 342254 122720 342260 122732
rect 324464 122692 342260 122720
rect 324464 122680 324470 122692
rect 342254 122680 342260 122692
rect 342312 122680 342318 122732
rect 252278 122612 252284 122664
rect 252336 122652 252342 122664
rect 262858 122652 262864 122664
rect 252336 122624 262864 122652
rect 252336 122612 252342 122624
rect 262858 122612 262864 122624
rect 262916 122612 262922 122664
rect 279418 122068 279424 122120
rect 279476 122108 279482 122120
rect 308490 122108 308496 122120
rect 279476 122080 308496 122108
rect 279476 122068 279482 122080
rect 308490 122068 308496 122080
rect 308548 122068 308554 122120
rect 298738 121592 298744 121644
rect 298796 121632 298802 121644
rect 307662 121632 307668 121644
rect 298796 121604 307668 121632
rect 298796 121592 298802 121604
rect 307662 121592 307668 121604
rect 307720 121592 307726 121644
rect 203518 121524 203524 121576
rect 203576 121564 203582 121576
rect 214006 121564 214012 121576
rect 203576 121536 214012 121564
rect 203576 121524 203582 121536
rect 214006 121524 214012 121536
rect 214064 121524 214070 121576
rect 297450 121524 297456 121576
rect 297508 121564 297514 121576
rect 307478 121564 307484 121576
rect 297508 121536 307484 121564
rect 297508 121524 297514 121536
rect 307478 121524 307484 121536
rect 307536 121524 307542 121576
rect 166442 121456 166448 121508
rect 166500 121496 166506 121508
rect 213914 121496 213920 121508
rect 166500 121468 213920 121496
rect 166500 121456 166506 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 269850 121456 269856 121508
rect 269908 121496 269914 121508
rect 307570 121496 307576 121508
rect 269908 121468 307576 121496
rect 269908 121456 269914 121468
rect 307570 121456 307576 121468
rect 307628 121456 307634 121508
rect 252462 121388 252468 121440
rect 252520 121428 252526 121440
rect 287974 121428 287980 121440
rect 252520 121400 287980 121428
rect 252520 121388 252526 121400
rect 287974 121388 287980 121400
rect 288032 121388 288038 121440
rect 324314 121388 324320 121440
rect 324372 121428 324378 121440
rect 335354 121428 335360 121440
rect 324372 121400 335360 121428
rect 324372 121388 324378 121400
rect 335354 121388 335360 121400
rect 335412 121388 335418 121440
rect 407758 121388 407764 121440
rect 407816 121428 407822 121440
rect 416774 121428 416780 121440
rect 407816 121400 416780 121428
rect 407816 121388 407822 121400
rect 416774 121388 416780 121400
rect 416832 121388 416838 121440
rect 252462 120300 252468 120352
rect 252520 120340 252526 120352
rect 260466 120340 260472 120352
rect 252520 120312 260472 120340
rect 252520 120300 252526 120312
rect 260466 120300 260472 120312
rect 260524 120300 260530 120352
rect 287882 120232 287888 120284
rect 287940 120272 287946 120284
rect 307662 120272 307668 120284
rect 287940 120244 307668 120272
rect 287940 120232 287946 120244
rect 307662 120232 307668 120244
rect 307720 120232 307726 120284
rect 183002 120164 183008 120216
rect 183060 120204 183066 120216
rect 214006 120204 214012 120216
rect 183060 120176 214012 120204
rect 183060 120164 183066 120176
rect 214006 120164 214012 120176
rect 214064 120164 214070 120216
rect 268378 120164 268384 120216
rect 268436 120204 268442 120216
rect 307478 120204 307484 120216
rect 268436 120176 307484 120204
rect 268436 120164 268442 120176
rect 307478 120164 307484 120176
rect 307536 120164 307542 120216
rect 57882 120096 57888 120148
rect 57940 120136 57946 120148
rect 65150 120136 65156 120148
rect 57940 120108 65156 120136
rect 57940 120096 57946 120108
rect 65150 120096 65156 120108
rect 65208 120096 65214 120148
rect 169018 120096 169024 120148
rect 169076 120136 169082 120148
rect 213914 120136 213920 120148
rect 169076 120108 213920 120136
rect 169076 120096 169082 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 260098 120096 260104 120148
rect 260156 120136 260162 120148
rect 307570 120136 307576 120148
rect 260156 120108 307576 120136
rect 260156 120096 260162 120108
rect 307570 120096 307576 120108
rect 307628 120096 307634 120148
rect 252462 120028 252468 120080
rect 252520 120068 252526 120080
rect 273898 120068 273904 120080
rect 252520 120040 273904 120068
rect 252520 120028 252526 120040
rect 273898 120028 273904 120040
rect 273956 120028 273962 120080
rect 324314 119960 324320 120012
rect 324372 120000 324378 120012
rect 325970 120000 325976 120012
rect 324372 119972 325976 120000
rect 324372 119960 324378 119972
rect 325970 119960 325976 119972
rect 326028 119960 326034 120012
rect 496906 119552 496912 119604
rect 496964 119592 496970 119604
rect 500954 119592 500960 119604
rect 496964 119564 500960 119592
rect 496964 119552 496970 119564
rect 500954 119552 500960 119564
rect 501012 119552 501018 119604
rect 263042 119416 263048 119468
rect 263100 119456 263106 119468
rect 307110 119456 307116 119468
rect 263100 119428 307116 119456
rect 263100 119416 263106 119428
rect 307110 119416 307116 119428
rect 307168 119416 307174 119468
rect 251910 119348 251916 119400
rect 251968 119388 251974 119400
rect 304350 119388 304356 119400
rect 251968 119360 304356 119388
rect 251968 119348 251974 119360
rect 304350 119348 304356 119360
rect 304408 119348 304414 119400
rect 252462 118940 252468 118992
rect 252520 118980 252526 118992
rect 260374 118980 260380 118992
rect 252520 118952 260380 118980
rect 252520 118940 252526 118952
rect 260374 118940 260380 118952
rect 260432 118940 260438 118992
rect 170582 118804 170588 118856
rect 170640 118844 170646 118856
rect 214006 118844 214012 118856
rect 170640 118816 214012 118844
rect 170640 118804 170646 118816
rect 214006 118804 214012 118816
rect 214064 118804 214070 118856
rect 278314 118804 278320 118856
rect 278372 118844 278378 118856
rect 307662 118844 307668 118856
rect 278372 118816 307668 118844
rect 278372 118804 278378 118816
rect 307662 118804 307668 118816
rect 307720 118804 307726 118856
rect 178862 118736 178868 118788
rect 178920 118776 178926 118788
rect 213914 118776 213920 118788
rect 178920 118748 213920 118776
rect 178920 118736 178926 118748
rect 213914 118736 213920 118748
rect 213972 118736 213978 118788
rect 300302 118668 300308 118720
rect 300360 118708 300366 118720
rect 307478 118708 307484 118720
rect 300360 118680 307484 118708
rect 300360 118668 300366 118680
rect 307478 118668 307484 118680
rect 307536 118668 307542 118720
rect 252462 118600 252468 118652
rect 252520 118640 252526 118652
rect 290458 118640 290464 118652
rect 252520 118612 290464 118640
rect 252520 118600 252526 118612
rect 290458 118600 290464 118612
rect 290516 118600 290522 118652
rect 324406 118600 324412 118652
rect 324464 118640 324470 118652
rect 345106 118640 345112 118652
rect 324464 118612 345112 118640
rect 324464 118600 324470 118612
rect 345106 118600 345112 118612
rect 345164 118600 345170 118652
rect 371878 118600 371884 118652
rect 371936 118640 371942 118652
rect 416774 118640 416780 118652
rect 371936 118612 416780 118640
rect 371936 118600 371942 118612
rect 416774 118600 416780 118612
rect 416832 118600 416838 118652
rect 496814 118600 496820 118652
rect 496872 118640 496878 118652
rect 517514 118640 517520 118652
rect 496872 118612 517520 118640
rect 496872 118600 496878 118612
rect 517514 118600 517520 118612
rect 517572 118600 517578 118652
rect 252370 118532 252376 118584
rect 252428 118572 252434 118584
rect 257338 118572 257344 118584
rect 252428 118544 257344 118572
rect 252428 118532 252434 118544
rect 257338 118532 257344 118544
rect 257396 118532 257402 118584
rect 324314 118532 324320 118584
rect 324372 118572 324378 118584
rect 342346 118572 342352 118584
rect 324372 118544 342352 118572
rect 324372 118532 324378 118544
rect 342346 118532 342352 118544
rect 342404 118532 342410 118584
rect 252094 117920 252100 117972
rect 252152 117960 252158 117972
rect 275370 117960 275376 117972
rect 252152 117932 275376 117960
rect 252152 117920 252158 117932
rect 275370 117920 275376 117932
rect 275428 117920 275434 117972
rect 304534 117444 304540 117496
rect 304592 117484 304598 117496
rect 307570 117484 307576 117496
rect 304592 117456 307576 117484
rect 304592 117444 304598 117456
rect 307570 117444 307576 117456
rect 307628 117444 307634 117496
rect 203610 117376 203616 117428
rect 203668 117416 203674 117428
rect 213914 117416 213920 117428
rect 203668 117388 213920 117416
rect 203668 117376 203674 117388
rect 213914 117376 213920 117388
rect 213972 117376 213978 117428
rect 282362 117376 282368 117428
rect 282420 117416 282426 117428
rect 306558 117416 306564 117428
rect 282420 117388 306564 117416
rect 282420 117376 282426 117388
rect 306558 117376 306564 117388
rect 306616 117376 306622 117428
rect 173434 117308 173440 117360
rect 173492 117348 173498 117360
rect 214006 117348 214012 117360
rect 173492 117320 214012 117348
rect 173492 117308 173498 117320
rect 214006 117308 214012 117320
rect 214064 117308 214070 117360
rect 261662 117308 261668 117360
rect 261720 117348 261726 117360
rect 307662 117348 307668 117360
rect 261720 117320 307668 117348
rect 261720 117308 261726 117320
rect 307662 117308 307668 117320
rect 307720 117308 307726 117360
rect 252370 117240 252376 117292
rect 252428 117280 252434 117292
rect 277026 117280 277032 117292
rect 252428 117252 277032 117280
rect 252428 117240 252434 117252
rect 277026 117240 277032 117252
rect 277084 117240 277090 117292
rect 340230 117240 340236 117292
rect 340288 117280 340294 117292
rect 416774 117280 416780 117292
rect 340288 117252 416780 117280
rect 340288 117240 340294 117252
rect 416774 117240 416780 117252
rect 416832 117240 416838 117292
rect 496814 117240 496820 117292
rect 496872 117280 496878 117292
rect 503806 117280 503812 117292
rect 496872 117252 503812 117280
rect 496872 117240 496878 117252
rect 503806 117240 503812 117252
rect 503864 117240 503870 117292
rect 252278 117172 252284 117224
rect 252336 117212 252342 117224
rect 266998 117212 267004 117224
rect 252336 117184 267004 117212
rect 252336 117172 252342 117184
rect 266998 117172 267004 117184
rect 267056 117172 267062 117224
rect 324406 117172 324412 117224
rect 324464 117212 324470 117224
rect 338114 117212 338120 117224
rect 324464 117184 338120 117212
rect 324464 117172 324470 117184
rect 338114 117172 338120 117184
rect 338172 117172 338178 117224
rect 324314 117104 324320 117156
rect 324372 117144 324378 117156
rect 340966 117144 340972 117156
rect 324372 117116 340972 117144
rect 324372 117104 324378 117116
rect 340966 117104 340972 117116
rect 341024 117104 341030 117156
rect 252462 116832 252468 116884
rect 252520 116872 252526 116884
rect 260282 116872 260288 116884
rect 252520 116844 260288 116872
rect 252520 116832 252526 116844
rect 260282 116832 260288 116844
rect 260340 116832 260346 116884
rect 276842 116084 276848 116136
rect 276900 116124 276906 116136
rect 306742 116124 306748 116136
rect 276900 116096 306748 116124
rect 276900 116084 276906 116096
rect 306742 116084 306748 116096
rect 306800 116084 306806 116136
rect 207842 116016 207848 116068
rect 207900 116056 207906 116068
rect 213914 116056 213920 116068
rect 207900 116028 213920 116056
rect 207900 116016 207906 116028
rect 213914 116016 213920 116028
rect 213972 116016 213978 116068
rect 273898 116016 273904 116068
rect 273956 116056 273962 116068
rect 307662 116056 307668 116068
rect 273956 116028 307668 116056
rect 273956 116016 273962 116028
rect 307662 116016 307668 116028
rect 307720 116016 307726 116068
rect 181622 115948 181628 116000
rect 181680 115988 181686 116000
rect 214006 115988 214012 116000
rect 181680 115960 214012 115988
rect 181680 115948 181686 115960
rect 214006 115948 214012 115960
rect 214064 115948 214070 116000
rect 258718 115948 258724 116000
rect 258776 115988 258782 116000
rect 307570 115988 307576 116000
rect 258776 115960 307576 115988
rect 258776 115948 258782 115960
rect 307570 115948 307576 115960
rect 307628 115948 307634 116000
rect 252462 115880 252468 115932
rect 252520 115920 252526 115932
rect 281074 115920 281080 115932
rect 252520 115892 281080 115920
rect 252520 115880 252526 115892
rect 281074 115880 281080 115892
rect 281132 115880 281138 115932
rect 324406 115880 324412 115932
rect 324464 115920 324470 115932
rect 343726 115920 343732 115932
rect 324464 115892 343732 115920
rect 324464 115880 324470 115892
rect 343726 115880 343732 115892
rect 343784 115880 343790 115932
rect 252370 115812 252376 115864
rect 252428 115852 252434 115864
rect 271230 115852 271236 115864
rect 252428 115824 271236 115852
rect 252428 115812 252434 115824
rect 271230 115812 271236 115824
rect 271288 115812 271294 115864
rect 324314 115812 324320 115864
rect 324372 115852 324378 115864
rect 332686 115852 332692 115864
rect 324372 115824 332692 115852
rect 324372 115812 324378 115824
rect 332686 115812 332692 115824
rect 332744 115812 332750 115864
rect 290458 114656 290464 114708
rect 290516 114696 290522 114708
rect 307662 114696 307668 114708
rect 290516 114668 307668 114696
rect 290516 114656 290522 114668
rect 307662 114656 307668 114668
rect 307720 114656 307726 114708
rect 280890 114588 280896 114640
rect 280948 114628 280954 114640
rect 307570 114628 307576 114640
rect 280948 114600 307576 114628
rect 280948 114588 280954 114600
rect 307570 114588 307576 114600
rect 307628 114588 307634 114640
rect 195514 114520 195520 114572
rect 195572 114560 195578 114572
rect 213914 114560 213920 114572
rect 195572 114532 213920 114560
rect 195572 114520 195578 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 252370 114520 252376 114572
rect 252428 114560 252434 114572
rect 258902 114560 258908 114572
rect 252428 114532 258908 114560
rect 252428 114520 252434 114532
rect 258902 114520 258908 114532
rect 258960 114520 258966 114572
rect 271138 114520 271144 114572
rect 271196 114560 271202 114572
rect 307478 114560 307484 114572
rect 271196 114532 307484 114560
rect 271196 114520 271202 114532
rect 307478 114520 307484 114532
rect 307536 114520 307542 114572
rect 252462 114452 252468 114504
rect 252520 114492 252526 114504
rect 261754 114492 261760 114504
rect 252520 114464 261760 114492
rect 252520 114452 252526 114464
rect 261754 114452 261760 114464
rect 261812 114452 261818 114504
rect 324406 114452 324412 114504
rect 324464 114492 324470 114504
rect 345014 114492 345020 114504
rect 324464 114464 345020 114492
rect 324464 114452 324470 114464
rect 345014 114452 345020 114464
rect 345072 114452 345078 114504
rect 385678 114452 385684 114504
rect 385736 114492 385742 114504
rect 416774 114492 416780 114504
rect 385736 114464 416780 114492
rect 385736 114452 385742 114464
rect 416774 114452 416780 114464
rect 416832 114452 416838 114504
rect 324314 114384 324320 114436
rect 324372 114424 324378 114436
rect 341150 114424 341156 114436
rect 324372 114396 341156 114424
rect 324372 114384 324378 114396
rect 341150 114384 341156 114396
rect 341208 114384 341214 114436
rect 496814 114180 496820 114232
rect 496872 114220 496878 114232
rect 499666 114220 499672 114232
rect 496872 114192 499672 114220
rect 496872 114180 496878 114192
rect 499666 114180 499672 114192
rect 499724 114180 499730 114232
rect 252462 113772 252468 113824
rect 252520 113812 252526 113824
rect 268470 113812 268476 113824
rect 252520 113784 268476 113812
rect 252520 113772 252526 113784
rect 268470 113772 268476 113784
rect 268528 113772 268534 113824
rect 291930 113296 291936 113348
rect 291988 113336 291994 113348
rect 307662 113336 307668 113348
rect 291988 113308 307668 113336
rect 291988 113296 291994 113308
rect 307662 113296 307668 113308
rect 307720 113296 307726 113348
rect 200942 113228 200948 113280
rect 201000 113268 201006 113280
rect 214006 113268 214012 113280
rect 201000 113240 214012 113268
rect 201000 113228 201006 113240
rect 214006 113228 214012 113240
rect 214064 113228 214070 113280
rect 265710 113228 265716 113280
rect 265768 113268 265774 113280
rect 307570 113268 307576 113280
rect 265768 113240 307576 113268
rect 265768 113228 265774 113240
rect 307570 113228 307576 113240
rect 307628 113228 307634 113280
rect 196894 113160 196900 113212
rect 196952 113200 196958 113212
rect 213914 113200 213920 113212
rect 196952 113172 213920 113200
rect 196952 113160 196958 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 249058 113160 249064 113212
rect 249116 113200 249122 113212
rect 307662 113200 307668 113212
rect 249116 113172 307668 113200
rect 249116 113160 249122 113172
rect 307662 113160 307668 113172
rect 307720 113160 307726 113212
rect 324314 113092 324320 113144
rect 324372 113132 324378 113144
rect 349154 113132 349160 113144
rect 324372 113104 349160 113132
rect 324372 113092 324378 113104
rect 349154 113092 349160 113104
rect 349212 113092 349218 113144
rect 252462 112888 252468 112940
rect 252520 112928 252526 112940
rect 255958 112928 255964 112940
rect 252520 112900 255964 112928
rect 252520 112888 252526 112900
rect 255958 112888 255964 112900
rect 256016 112888 256022 112940
rect 413278 112888 413284 112940
rect 413336 112928 413342 112940
rect 416774 112928 416780 112940
rect 413336 112900 416780 112928
rect 413336 112888 413342 112900
rect 416774 112888 416780 112900
rect 416832 112888 416838 112940
rect 252094 112480 252100 112532
rect 252152 112520 252158 112532
rect 289262 112520 289268 112532
rect 252152 112492 289268 112520
rect 252152 112480 252158 112492
rect 289262 112480 289268 112492
rect 289320 112480 289326 112532
rect 252186 112412 252192 112464
rect 252244 112452 252250 112464
rect 304258 112452 304264 112464
rect 252244 112424 304264 112452
rect 252244 112412 252250 112424
rect 304258 112412 304264 112424
rect 304316 112412 304322 112464
rect 205174 111868 205180 111920
rect 205232 111908 205238 111920
rect 213914 111908 213920 111920
rect 205232 111880 213920 111908
rect 205232 111868 205238 111880
rect 213914 111868 213920 111880
rect 213972 111868 213978 111920
rect 252462 111868 252468 111920
rect 252520 111908 252526 111920
rect 258810 111908 258816 111920
rect 252520 111880 258816 111908
rect 252520 111868 252526 111880
rect 258810 111868 258816 111880
rect 258868 111868 258874 111920
rect 304350 111868 304356 111920
rect 304408 111908 304414 111920
rect 307662 111908 307668 111920
rect 304408 111880 307668 111908
rect 304408 111868 304414 111880
rect 307662 111868 307668 111880
rect 307720 111868 307726 111920
rect 174722 111800 174728 111852
rect 174780 111840 174786 111852
rect 214006 111840 214012 111852
rect 174780 111812 214012 111840
rect 174780 111800 174786 111812
rect 214006 111800 214012 111812
rect 214064 111800 214070 111852
rect 266998 111800 267004 111852
rect 267056 111840 267062 111852
rect 306926 111840 306932 111852
rect 267056 111812 306932 111840
rect 267056 111800 267062 111812
rect 306926 111800 306932 111812
rect 306984 111800 306990 111852
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 11698 111772 11704 111784
rect 3476 111744 11704 111772
rect 3476 111732 3482 111744
rect 11698 111732 11704 111744
rect 11756 111732 11762 111784
rect 167914 111732 167920 111784
rect 167972 111772 167978 111784
rect 205082 111772 205088 111784
rect 167972 111744 205088 111772
rect 167972 111732 167978 111744
rect 205082 111732 205088 111744
rect 205140 111732 205146 111784
rect 252462 111732 252468 111784
rect 252520 111772 252526 111784
rect 296070 111772 296076 111784
rect 252520 111744 296076 111772
rect 252520 111732 252526 111744
rect 296070 111732 296076 111744
rect 296128 111732 296134 111784
rect 324314 111732 324320 111784
rect 324372 111772 324378 111784
rect 336826 111772 336832 111784
rect 324372 111744 336832 111772
rect 324372 111732 324378 111744
rect 336826 111732 336832 111744
rect 336884 111732 336890 111784
rect 388438 111732 388444 111784
rect 388496 111772 388502 111784
rect 416774 111772 416780 111784
rect 388496 111744 416780 111772
rect 388496 111732 388502 111744
rect 416774 111732 416780 111744
rect 416832 111732 416838 111784
rect 496814 111732 496820 111784
rect 496872 111772 496878 111784
rect 506474 111772 506480 111784
rect 496872 111744 506480 111772
rect 496872 111732 496878 111744
rect 506474 111732 506480 111744
rect 506532 111732 506538 111784
rect 252278 111664 252284 111716
rect 252336 111704 252342 111716
rect 254578 111704 254584 111716
rect 252336 111676 254584 111704
rect 252336 111664 252342 111676
rect 254578 111664 254584 111676
rect 254636 111664 254642 111716
rect 324406 111664 324412 111716
rect 324464 111704 324470 111716
rect 336734 111704 336740 111716
rect 324464 111676 336740 111704
rect 324464 111664 324470 111676
rect 336734 111664 336740 111676
rect 336792 111664 336798 111716
rect 496814 111596 496820 111648
rect 496872 111636 496878 111648
rect 501138 111636 501144 111648
rect 496872 111608 501144 111636
rect 496872 111596 496878 111608
rect 501138 111596 501144 111608
rect 501196 111596 501202 111648
rect 294782 110576 294788 110628
rect 294840 110616 294846 110628
rect 307478 110616 307484 110628
rect 294840 110588 307484 110616
rect 294840 110576 294846 110588
rect 307478 110576 307484 110588
rect 307536 110576 307542 110628
rect 176194 110508 176200 110560
rect 176252 110548 176258 110560
rect 213914 110548 213920 110560
rect 176252 110520 213920 110548
rect 176252 110508 176258 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 273990 110508 273996 110560
rect 274048 110548 274054 110560
rect 307570 110548 307576 110560
rect 274048 110520 307576 110548
rect 274048 110508 274054 110520
rect 307570 110508 307576 110520
rect 307628 110508 307634 110560
rect 166534 110440 166540 110492
rect 166592 110480 166598 110492
rect 214006 110480 214012 110492
rect 166592 110452 214012 110480
rect 166592 110440 166598 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 253382 110440 253388 110492
rect 253440 110480 253446 110492
rect 307662 110480 307668 110492
rect 253440 110452 307668 110480
rect 253440 110440 253446 110452
rect 307662 110440 307668 110452
rect 307720 110440 307726 110492
rect 252278 110372 252284 110424
rect 252336 110412 252342 110424
rect 305822 110412 305828 110424
rect 252336 110384 305828 110412
rect 252336 110372 252342 110384
rect 305822 110372 305828 110384
rect 305880 110372 305886 110424
rect 324314 110372 324320 110424
rect 324372 110412 324378 110424
rect 341058 110412 341064 110424
rect 324372 110384 341064 110412
rect 324372 110372 324378 110384
rect 341058 110372 341064 110384
rect 341116 110372 341122 110424
rect 377398 110372 377404 110424
rect 377456 110412 377462 110424
rect 416774 110412 416780 110424
rect 377456 110384 416780 110412
rect 377456 110372 377462 110384
rect 416774 110372 416780 110384
rect 416832 110372 416838 110424
rect 496814 110372 496820 110424
rect 496872 110412 496878 110424
rect 510614 110412 510620 110424
rect 496872 110384 510620 110412
rect 496872 110372 496878 110384
rect 510614 110372 510620 110384
rect 510672 110372 510678 110424
rect 252370 110304 252376 110356
rect 252428 110344 252434 110356
rect 298922 110344 298928 110356
rect 252428 110316 298928 110344
rect 252428 110304 252434 110316
rect 298922 110304 298928 110316
rect 298980 110304 298986 110356
rect 252462 110236 252468 110288
rect 252520 110276 252526 110288
rect 279510 110276 279516 110288
rect 252520 110248 279516 110276
rect 252520 110236 252526 110248
rect 279510 110236 279516 110248
rect 279568 110236 279574 110288
rect 324406 109692 324412 109744
rect 324464 109732 324470 109744
rect 328454 109732 328460 109744
rect 324464 109704 328460 109732
rect 324464 109692 324470 109704
rect 328454 109692 328460 109704
rect 328512 109692 328518 109744
rect 174814 109080 174820 109132
rect 174872 109120 174878 109132
rect 213914 109120 213920 109132
rect 174872 109092 213920 109120
rect 174872 109080 174878 109092
rect 213914 109080 213920 109092
rect 213972 109080 213978 109132
rect 302878 109080 302884 109132
rect 302936 109120 302942 109132
rect 306926 109120 306932 109132
rect 302936 109092 306932 109120
rect 302936 109080 302942 109092
rect 306926 109080 306932 109092
rect 306984 109080 306990 109132
rect 167822 109012 167828 109064
rect 167880 109052 167886 109064
rect 214006 109052 214012 109064
rect 167880 109024 214012 109052
rect 167880 109012 167886 109024
rect 214006 109012 214012 109024
rect 214064 109012 214070 109064
rect 289262 109012 289268 109064
rect 289320 109052 289326 109064
rect 307662 109052 307668 109064
rect 289320 109024 307668 109052
rect 289320 109012 289326 109024
rect 307662 109012 307668 109024
rect 307720 109012 307726 109064
rect 168098 108944 168104 108996
rect 168156 108984 168162 108996
rect 180242 108984 180248 108996
rect 168156 108956 180248 108984
rect 168156 108944 168162 108956
rect 180242 108944 180248 108956
rect 180300 108944 180306 108996
rect 252462 108944 252468 108996
rect 252520 108984 252526 108996
rect 283650 108984 283656 108996
rect 252520 108956 283656 108984
rect 252520 108944 252526 108956
rect 283650 108944 283656 108956
rect 283708 108944 283714 108996
rect 251726 108876 251732 108928
rect 251784 108916 251790 108928
rect 254854 108916 254860 108928
rect 251784 108888 254860 108916
rect 251784 108876 251790 108888
rect 254854 108876 254860 108888
rect 254912 108876 254918 108928
rect 251818 108332 251824 108384
rect 251876 108372 251882 108384
rect 256234 108372 256240 108384
rect 251876 108344 256240 108372
rect 251876 108332 251882 108344
rect 256234 108332 256240 108344
rect 256292 108332 256298 108384
rect 324314 108196 324320 108248
rect 324372 108236 324378 108248
rect 327166 108236 327172 108248
rect 324372 108208 327172 108236
rect 324372 108196 324378 108208
rect 327166 108196 327172 108208
rect 327224 108196 327230 108248
rect 255958 107856 255964 107908
rect 256016 107896 256022 107908
rect 307662 107896 307668 107908
rect 256016 107868 307668 107896
rect 256016 107856 256022 107868
rect 307662 107856 307668 107868
rect 307720 107856 307726 107908
rect 180426 107720 180432 107772
rect 180484 107760 180490 107772
rect 214006 107760 214012 107772
rect 180484 107732 214012 107760
rect 180484 107720 180490 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 279418 107720 279424 107772
rect 279476 107760 279482 107772
rect 307662 107760 307668 107772
rect 279476 107732 307668 107760
rect 279476 107720 279482 107732
rect 307662 107720 307668 107732
rect 307720 107720 307726 107772
rect 169202 107652 169208 107704
rect 169260 107692 169266 107704
rect 213914 107692 213920 107704
rect 169260 107664 213920 107692
rect 169260 107652 169266 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 302970 107652 302976 107704
rect 303028 107692 303034 107704
rect 307570 107692 307576 107704
rect 303028 107664 307576 107692
rect 303028 107652 303034 107664
rect 307570 107652 307576 107664
rect 307628 107652 307634 107704
rect 252462 107584 252468 107636
rect 252520 107624 252526 107636
rect 265618 107624 265624 107636
rect 252520 107596 265624 107624
rect 252520 107584 252526 107596
rect 265618 107584 265624 107596
rect 265676 107584 265682 107636
rect 324314 107584 324320 107636
rect 324372 107624 324378 107636
rect 354674 107624 354680 107636
rect 324372 107596 354680 107624
rect 324372 107584 324378 107596
rect 354674 107584 354680 107596
rect 354732 107584 354738 107636
rect 389818 107584 389824 107636
rect 389876 107624 389882 107636
rect 416774 107624 416780 107636
rect 389876 107596 416780 107624
rect 389876 107584 389882 107596
rect 416774 107584 416780 107596
rect 416832 107584 416838 107636
rect 496814 107584 496820 107636
rect 496872 107624 496878 107636
rect 502334 107624 502340 107636
rect 496872 107596 502340 107624
rect 496872 107584 496878 107596
rect 502334 107584 502340 107596
rect 502392 107584 502398 107636
rect 251726 107516 251732 107568
rect 251784 107556 251790 107568
rect 254762 107556 254768 107568
rect 251784 107528 254768 107556
rect 251784 107516 251790 107528
rect 254762 107516 254768 107528
rect 254820 107516 254826 107568
rect 304258 106428 304264 106480
rect 304316 106468 304322 106480
rect 307570 106468 307576 106480
rect 304316 106440 307576 106468
rect 304316 106428 304322 106440
rect 307570 106428 307576 106440
rect 307628 106428 307634 106480
rect 176102 106360 176108 106412
rect 176160 106400 176166 106412
rect 214006 106400 214012 106412
rect 176160 106372 214012 106400
rect 176160 106360 176166 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 254578 106360 254584 106412
rect 254636 106400 254642 106412
rect 307478 106400 307484 106412
rect 254636 106372 307484 106400
rect 254636 106360 254642 106372
rect 307478 106360 307484 106372
rect 307536 106360 307542 106412
rect 170674 106292 170680 106344
rect 170732 106332 170738 106344
rect 213914 106332 213920 106344
rect 170732 106304 213920 106332
rect 170732 106292 170738 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 250714 106292 250720 106344
rect 250772 106332 250778 106344
rect 307662 106332 307668 106344
rect 250772 106304 307668 106332
rect 250772 106292 250778 106304
rect 307662 106292 307668 106304
rect 307720 106292 307726 106344
rect 252370 106224 252376 106276
rect 252428 106264 252434 106276
rect 285122 106264 285128 106276
rect 252428 106236 285128 106264
rect 252428 106224 252434 106236
rect 285122 106224 285128 106236
rect 285180 106224 285186 106276
rect 342898 106224 342904 106276
rect 342956 106264 342962 106276
rect 416774 106264 416780 106276
rect 342956 106236 416780 106264
rect 342956 106224 342962 106236
rect 416774 106224 416780 106236
rect 416832 106224 416838 106276
rect 252462 106156 252468 106208
rect 252520 106196 252526 106208
rect 265802 106196 265808 106208
rect 252520 106168 265808 106196
rect 252520 106156 252526 106168
rect 265802 106156 265808 106168
rect 265860 106156 265866 106208
rect 252278 106088 252284 106140
rect 252336 106128 252342 106140
rect 257522 106128 257528 106140
rect 252336 106100 257528 106128
rect 252336 106088 252342 106100
rect 257522 106088 257528 106100
rect 257580 106088 257586 106140
rect 283650 105000 283656 105052
rect 283708 105040 283714 105052
rect 307478 105040 307484 105052
rect 283708 105012 307484 105040
rect 283708 105000 283714 105012
rect 307478 105000 307484 105012
rect 307536 105000 307542 105052
rect 192570 104932 192576 104984
rect 192628 104972 192634 104984
rect 213914 104972 213920 104984
rect 192628 104944 213920 104972
rect 192628 104932 192634 104944
rect 213914 104932 213920 104944
rect 213972 104932 213978 104984
rect 265618 104932 265624 104984
rect 265676 104972 265682 104984
rect 307662 104972 307668 104984
rect 265676 104944 307668 104972
rect 265676 104932 265682 104944
rect 307662 104932 307668 104944
rect 307720 104932 307726 104984
rect 172054 104864 172060 104916
rect 172112 104904 172118 104916
rect 214006 104904 214012 104916
rect 172112 104876 214012 104904
rect 172112 104864 172118 104876
rect 214006 104864 214012 104876
rect 214064 104864 214070 104916
rect 257338 104864 257344 104916
rect 257396 104904 257402 104916
rect 306926 104904 306932 104916
rect 257396 104876 306932 104904
rect 257396 104864 257402 104876
rect 306926 104864 306932 104876
rect 306984 104864 306990 104916
rect 252370 104796 252376 104848
rect 252428 104836 252434 104848
rect 276934 104836 276940 104848
rect 252428 104808 276940 104836
rect 252428 104796 252434 104808
rect 276934 104796 276940 104808
rect 276992 104796 276998 104848
rect 356698 104796 356704 104848
rect 356756 104836 356762 104848
rect 416774 104836 416780 104848
rect 356756 104808 416780 104836
rect 356756 104796 356762 104808
rect 416774 104796 416780 104808
rect 416832 104796 416838 104848
rect 252462 104728 252468 104780
rect 252520 104768 252526 104780
rect 272610 104768 272616 104780
rect 252520 104740 272616 104768
rect 252520 104728 252526 104740
rect 272610 104728 272616 104740
rect 272668 104728 272674 104780
rect 252278 104660 252284 104712
rect 252336 104700 252342 104712
rect 256142 104700 256148 104712
rect 252336 104672 256148 104700
rect 252336 104660 252342 104672
rect 256142 104660 256148 104672
rect 256200 104660 256206 104712
rect 325694 104116 325700 104168
rect 325752 104156 325758 104168
rect 354030 104156 354036 104168
rect 325752 104128 354036 104156
rect 325752 104116 325758 104128
rect 354030 104116 354036 104128
rect 354088 104116 354094 104168
rect 276750 103640 276756 103692
rect 276808 103680 276814 103692
rect 306926 103680 306932 103692
rect 276808 103652 306932 103680
rect 276808 103640 276814 103652
rect 306926 103640 306932 103652
rect 306984 103640 306990 103692
rect 275370 103572 275376 103624
rect 275428 103612 275434 103624
rect 307662 103612 307668 103624
rect 275428 103584 307668 103612
rect 275428 103572 275434 103584
rect 307662 103572 307668 103584
rect 307720 103572 307726 103624
rect 199470 103504 199476 103556
rect 199528 103544 199534 103556
rect 213914 103544 213920 103556
rect 199528 103516 213920 103544
rect 199528 103504 199534 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 267182 103504 267188 103556
rect 267240 103544 267246 103556
rect 307570 103544 307576 103556
rect 267240 103516 307576 103544
rect 267240 103504 267246 103516
rect 307570 103504 307576 103516
rect 307628 103504 307634 103556
rect 252462 103436 252468 103488
rect 252520 103476 252526 103488
rect 303154 103476 303160 103488
rect 252520 103448 303160 103476
rect 252520 103436 252526 103448
rect 303154 103436 303160 103448
rect 303212 103436 303218 103488
rect 393958 103436 393964 103488
rect 394016 103476 394022 103488
rect 416774 103476 416780 103488
rect 394016 103448 416780 103476
rect 394016 103436 394022 103448
rect 416774 103436 416780 103448
rect 416832 103436 416838 103488
rect 252370 103028 252376 103080
rect 252428 103068 252434 103080
rect 256050 103068 256056 103080
rect 252428 103040 256056 103068
rect 252428 103028 252434 103040
rect 256050 103028 256056 103040
rect 256108 103028 256114 103080
rect 252462 102892 252468 102944
rect 252520 102932 252526 102944
rect 260190 102932 260196 102944
rect 252520 102904 260196 102932
rect 252520 102892 252526 102904
rect 260190 102892 260196 102904
rect 260248 102892 260254 102944
rect 323578 102756 323584 102808
rect 323636 102796 323642 102808
rect 367830 102796 367836 102808
rect 323636 102768 367836 102796
rect 323636 102756 323642 102768
rect 367830 102756 367836 102768
rect 367888 102756 367894 102808
rect 297542 102212 297548 102264
rect 297600 102252 297606 102264
rect 307662 102252 307668 102264
rect 297600 102224 307668 102252
rect 297600 102212 297606 102224
rect 307662 102212 307668 102224
rect 307720 102212 307726 102264
rect 211982 102144 211988 102196
rect 212040 102184 212046 102196
rect 213914 102184 213920 102196
rect 212040 102156 213920 102184
rect 212040 102144 212046 102156
rect 213914 102144 213920 102156
rect 213972 102144 213978 102196
rect 258902 102144 258908 102196
rect 258960 102184 258966 102196
rect 307570 102184 307576 102196
rect 258960 102156 307576 102184
rect 258960 102144 258966 102156
rect 307570 102144 307576 102156
rect 307628 102144 307634 102196
rect 252462 102076 252468 102128
rect 252520 102116 252526 102128
rect 269758 102116 269764 102128
rect 252520 102088 269764 102116
rect 252520 102076 252526 102088
rect 269758 102076 269764 102088
rect 269816 102076 269822 102128
rect 324314 102076 324320 102128
rect 324372 102116 324378 102128
rect 332962 102116 332968 102128
rect 324372 102088 332968 102116
rect 324372 102076 324378 102088
rect 332962 102076 332968 102088
rect 333020 102076 333026 102128
rect 396718 102076 396724 102128
rect 396776 102116 396782 102128
rect 416774 102116 416780 102128
rect 396776 102088 416780 102116
rect 396776 102076 396782 102088
rect 416774 102076 416780 102088
rect 416832 102076 416838 102128
rect 251358 102008 251364 102060
rect 251416 102048 251422 102060
rect 253290 102048 253296 102060
rect 251416 102020 253296 102048
rect 251416 102008 251422 102020
rect 253290 102008 253296 102020
rect 253348 102008 253354 102060
rect 252186 101396 252192 101448
rect 252244 101436 252250 101448
rect 267090 101436 267096 101448
rect 252244 101408 267096 101436
rect 252244 101396 252250 101408
rect 267090 101396 267096 101408
rect 267148 101396 267154 101448
rect 301590 100920 301596 100972
rect 301648 100960 301654 100972
rect 306558 100960 306564 100972
rect 301648 100932 306564 100960
rect 301648 100920 301654 100932
rect 306558 100920 306564 100932
rect 306616 100920 306622 100972
rect 285122 100852 285128 100904
rect 285180 100892 285186 100904
rect 307662 100892 307668 100904
rect 285180 100864 307668 100892
rect 285180 100852 285186 100864
rect 307662 100852 307668 100864
rect 307720 100852 307726 100904
rect 207750 100784 207756 100836
rect 207808 100824 207814 100836
rect 214006 100824 214012 100836
rect 207808 100796 214012 100824
rect 207808 100784 207814 100796
rect 214006 100784 214012 100796
rect 214064 100784 214070 100836
rect 269942 100784 269948 100836
rect 270000 100824 270006 100836
rect 307570 100824 307576 100836
rect 270000 100796 307576 100824
rect 270000 100784 270006 100796
rect 307570 100784 307576 100796
rect 307628 100784 307634 100836
rect 66162 100716 66168 100768
rect 66220 100756 66226 100768
rect 68278 100756 68284 100768
rect 66220 100728 68284 100756
rect 66220 100716 66226 100728
rect 68278 100716 68284 100728
rect 68336 100716 68342 100768
rect 205082 100716 205088 100768
rect 205140 100756 205146 100768
rect 213914 100756 213920 100768
rect 205140 100728 213920 100756
rect 205140 100716 205146 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 264422 100716 264428 100768
rect 264480 100756 264486 100768
rect 306926 100756 306932 100768
rect 264480 100728 306932 100756
rect 264480 100716 264486 100728
rect 306926 100716 306932 100728
rect 306984 100716 306990 100768
rect 252370 100648 252376 100700
rect 252428 100688 252434 100700
rect 286502 100688 286508 100700
rect 252428 100660 286508 100688
rect 252428 100648 252434 100660
rect 286502 100648 286508 100660
rect 286560 100648 286566 100700
rect 378778 100648 378784 100700
rect 378836 100688 378842 100700
rect 493962 100688 493968 100700
rect 378836 100660 493968 100688
rect 378836 100648 378842 100660
rect 493962 100648 493968 100660
rect 494020 100648 494026 100700
rect 520182 100648 520188 100700
rect 520240 100688 520246 100700
rect 580166 100688 580172 100700
rect 520240 100660 580172 100688
rect 520240 100648 520246 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 252278 100580 252284 100632
rect 252336 100620 252342 100632
rect 268562 100620 268568 100632
rect 252336 100592 268568 100620
rect 252336 100580 252342 100592
rect 268562 100580 268568 100592
rect 268620 100580 268626 100632
rect 395338 100580 395344 100632
rect 395396 100620 395402 100632
rect 494238 100620 494244 100632
rect 395396 100592 494244 100620
rect 395396 100580 395402 100592
rect 494238 100580 494244 100592
rect 494296 100580 494302 100632
rect 252462 100512 252468 100564
rect 252520 100552 252526 100564
rect 263042 100552 263048 100564
rect 252520 100524 263048 100552
rect 252520 100512 252526 100524
rect 263042 100512 263048 100524
rect 263100 100512 263106 100564
rect 330478 99968 330484 100020
rect 330536 100008 330542 100020
rect 370498 100008 370504 100020
rect 330536 99980 370504 100008
rect 330536 99968 330542 99980
rect 370498 99968 370504 99980
rect 370556 99968 370562 100020
rect 296070 99492 296076 99544
rect 296128 99532 296134 99544
rect 306558 99532 306564 99544
rect 296128 99504 306564 99532
rect 296128 99492 296134 99504
rect 306558 99492 306564 99504
rect 306616 99492 306622 99544
rect 272610 99424 272616 99476
rect 272668 99464 272674 99476
rect 307662 99464 307668 99476
rect 272668 99436 307668 99464
rect 272668 99424 272674 99436
rect 307662 99424 307668 99436
rect 307720 99424 307726 99476
rect 167730 99356 167736 99408
rect 167788 99396 167794 99408
rect 213914 99396 213920 99408
rect 167788 99368 213920 99396
rect 167788 99356 167794 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 262858 99356 262864 99408
rect 262916 99396 262922 99408
rect 307570 99396 307576 99408
rect 262916 99368 307576 99396
rect 262916 99356 262922 99368
rect 307570 99356 307576 99368
rect 307628 99356 307634 99408
rect 252462 99288 252468 99340
rect 252520 99328 252526 99340
rect 261478 99328 261484 99340
rect 252520 99300 261484 99328
rect 252520 99288 252526 99300
rect 261478 99288 261484 99300
rect 261536 99288 261542 99340
rect 324314 99288 324320 99340
rect 324372 99328 324378 99340
rect 339494 99328 339500 99340
rect 324372 99300 339500 99328
rect 324372 99288 324378 99300
rect 339494 99288 339500 99300
rect 339552 99288 339558 99340
rect 419626 99288 419632 99340
rect 419684 99328 419690 99340
rect 580258 99328 580264 99340
rect 419684 99300 580264 99328
rect 419684 99288 419690 99300
rect 580258 99288 580264 99300
rect 580316 99288 580322 99340
rect 399478 99220 399484 99272
rect 399536 99260 399542 99272
rect 496906 99260 496912 99272
rect 399536 99232 496912 99260
rect 399536 99220 399542 99232
rect 496906 99220 496912 99232
rect 496964 99220 496970 99272
rect 324406 98744 324412 98796
rect 324464 98784 324470 98796
rect 324682 98784 324688 98796
rect 324464 98756 324688 98784
rect 324464 98744 324470 98756
rect 324682 98744 324688 98756
rect 324740 98744 324746 98796
rect 169294 98608 169300 98660
rect 169352 98648 169358 98660
rect 214006 98648 214012 98660
rect 169352 98620 214012 98648
rect 169352 98608 169358 98620
rect 214006 98608 214012 98620
rect 214064 98608 214070 98660
rect 252462 98608 252468 98660
rect 252520 98648 252526 98660
rect 262950 98648 262956 98660
rect 252520 98620 262956 98648
rect 252520 98608 252526 98620
rect 262950 98608 262956 98620
rect 263008 98608 263014 98660
rect 324406 98608 324412 98660
rect 324464 98648 324470 98660
rect 331214 98648 331220 98660
rect 324464 98620 331220 98648
rect 324464 98608 324470 98620
rect 331214 98608 331220 98620
rect 331272 98608 331278 98660
rect 298922 98132 298928 98184
rect 298980 98172 298986 98184
rect 306926 98172 306932 98184
rect 298980 98144 306932 98172
rect 298980 98132 298986 98144
rect 306926 98132 306932 98144
rect 306984 98132 306990 98184
rect 264514 98064 264520 98116
rect 264572 98104 264578 98116
rect 307570 98104 307576 98116
rect 264572 98076 307576 98104
rect 264572 98064 264578 98076
rect 307570 98064 307576 98076
rect 307628 98064 307634 98116
rect 165246 97996 165252 98048
rect 165304 98036 165310 98048
rect 213914 98036 213920 98048
rect 165304 98008 213920 98036
rect 165304 97996 165310 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 256050 97996 256056 98048
rect 256108 98036 256114 98048
rect 307662 98036 307668 98048
rect 256108 98008 307668 98036
rect 256108 97996 256114 98008
rect 307662 97996 307668 98008
rect 307720 97996 307726 98048
rect 256694 97928 256700 97980
rect 256752 97968 256758 97980
rect 257430 97968 257436 97980
rect 256752 97940 257436 97968
rect 256752 97928 256758 97940
rect 257430 97928 257436 97940
rect 257488 97928 257494 97980
rect 324314 97928 324320 97980
rect 324372 97968 324378 97980
rect 350534 97968 350540 97980
rect 324372 97940 350540 97968
rect 324372 97928 324378 97940
rect 350534 97928 350540 97940
rect 350592 97928 350598 97980
rect 392578 97928 392584 97980
rect 392636 97968 392642 97980
rect 495434 97968 495440 97980
rect 392636 97940 495440 97968
rect 392636 97928 392642 97940
rect 495434 97928 495440 97940
rect 495492 97928 495498 97980
rect 410518 97860 410524 97912
rect 410576 97900 410582 97912
rect 496998 97900 497004 97912
rect 410576 97872 497004 97900
rect 410576 97860 410582 97872
rect 496998 97860 497004 97872
rect 497056 97860 497062 97912
rect 2774 97724 2780 97776
rect 2832 97764 2838 97776
rect 4798 97764 4804 97776
rect 2832 97736 4804 97764
rect 2832 97724 2838 97736
rect 4798 97724 4804 97736
rect 4856 97724 4862 97776
rect 420178 97316 420184 97368
rect 420236 97356 420242 97368
rect 427722 97356 427728 97368
rect 420236 97328 427728 97356
rect 420236 97316 420242 97328
rect 427722 97316 427728 97328
rect 427780 97316 427786 97368
rect 421558 97248 421564 97300
rect 421616 97288 421622 97300
rect 458910 97288 458916 97300
rect 421616 97260 458916 97288
rect 421616 97248 421622 97260
rect 458910 97248 458916 97260
rect 458968 97248 458974 97300
rect 467098 97248 467104 97300
rect 467156 97288 467162 97300
rect 492490 97288 492496 97300
rect 467156 97260 492496 97288
rect 467156 97248 467162 97260
rect 492490 97248 492496 97260
rect 492548 97248 492554 97300
rect 439498 96908 439504 96960
rect 439556 96948 439562 96960
rect 440878 96948 440884 96960
rect 439556 96920 440884 96948
rect 439556 96908 439562 96920
rect 440878 96908 440884 96920
rect 440936 96908 440942 96960
rect 454034 96908 454040 96960
rect 454092 96948 454098 96960
rect 455046 96948 455052 96960
rect 454092 96920 455052 96948
rect 454092 96908 454098 96920
rect 455046 96908 455052 96920
rect 455104 96908 455110 96960
rect 461578 96908 461584 96960
rect 461636 96948 461642 96960
rect 464890 96948 464896 96960
rect 461636 96920 464896 96948
rect 461636 96908 461642 96920
rect 464890 96908 464896 96920
rect 464948 96908 464954 96960
rect 465718 96908 465724 96960
rect 465776 96948 465782 96960
rect 467282 96948 467288 96960
rect 465776 96920 467288 96948
rect 465776 96908 465782 96920
rect 467282 96908 467288 96920
rect 467340 96908 467346 96960
rect 472618 96908 472624 96960
rect 472676 96948 472682 96960
rect 474550 96948 474556 96960
rect 472676 96920 474556 96948
rect 472676 96908 472682 96920
rect 474550 96908 474556 96920
rect 474608 96908 474614 96960
rect 481634 96908 481640 96960
rect 481692 96948 481698 96960
rect 482646 96948 482652 96960
rect 481692 96920 482652 96948
rect 481692 96908 481698 96920
rect 482646 96908 482652 96920
rect 482704 96908 482710 96960
rect 486418 96908 486424 96960
rect 486476 96948 486482 96960
rect 487706 96948 487712 96960
rect 486476 96920 487712 96948
rect 486476 96908 486482 96920
rect 487706 96908 487712 96920
rect 487764 96908 487770 96960
rect 417418 96772 417424 96824
rect 417476 96812 417482 96824
rect 420546 96812 420552 96824
rect 417476 96784 420552 96812
rect 417476 96772 417482 96784
rect 420546 96772 420552 96784
rect 420604 96772 420610 96824
rect 252462 96704 252468 96756
rect 252520 96744 252526 96756
rect 256694 96744 256700 96756
rect 252520 96716 256700 96744
rect 252520 96704 252526 96716
rect 256694 96704 256700 96716
rect 256752 96704 256758 96756
rect 269758 96704 269764 96756
rect 269816 96744 269822 96756
rect 307662 96744 307668 96756
rect 269816 96716 307668 96744
rect 269816 96704 269822 96716
rect 307662 96704 307668 96716
rect 307720 96704 307726 96756
rect 251818 96636 251824 96688
rect 251876 96676 251882 96688
rect 307478 96676 307484 96688
rect 251876 96648 307484 96676
rect 251876 96636 251882 96648
rect 307478 96636 307484 96648
rect 307536 96636 307542 96688
rect 282270 96568 282276 96620
rect 282328 96608 282334 96620
rect 321554 96608 321560 96620
rect 282328 96580 321560 96608
rect 282328 96568 282334 96580
rect 321554 96568 321560 96580
rect 321612 96568 321618 96620
rect 406378 96568 406384 96620
rect 406436 96608 406442 96620
rect 496814 96608 496820 96620
rect 406436 96580 496820 96608
rect 406436 96568 406442 96580
rect 496814 96568 496820 96580
rect 496872 96568 496878 96620
rect 309778 96500 309784 96552
rect 309836 96540 309842 96552
rect 322934 96540 322940 96552
rect 309836 96512 322940 96540
rect 309836 96500 309842 96512
rect 322934 96500 322940 96512
rect 322992 96500 322998 96552
rect 308398 96432 308404 96484
rect 308456 96472 308462 96484
rect 321646 96472 321652 96484
rect 308456 96444 321652 96472
rect 308456 96432 308462 96444
rect 321646 96432 321652 96444
rect 321704 96432 321710 96484
rect 184290 95956 184296 96008
rect 184348 95996 184354 96008
rect 222838 95996 222844 96008
rect 184348 95968 222844 95996
rect 184348 95956 184354 95968
rect 222838 95956 222844 95968
rect 222896 95956 222902 96008
rect 168282 95888 168288 95940
rect 168340 95928 168346 95940
rect 214558 95928 214564 95940
rect 168340 95900 214564 95928
rect 168340 95888 168346 95900
rect 214558 95888 214564 95900
rect 214616 95888 214622 95940
rect 343634 95888 343640 95940
rect 343692 95928 343698 95940
rect 498470 95928 498476 95940
rect 343692 95900 498476 95928
rect 343692 95888 343698 95900
rect 498470 95888 498476 95900
rect 498528 95888 498534 95940
rect 249242 95208 249248 95260
rect 249300 95248 249306 95260
rect 307662 95248 307668 95260
rect 249300 95220 307668 95248
rect 249300 95208 249306 95220
rect 307662 95208 307668 95220
rect 307720 95208 307726 95260
rect 198182 95140 198188 95192
rect 198240 95180 198246 95192
rect 321462 95180 321468 95192
rect 198240 95152 321468 95180
rect 198240 95140 198246 95152
rect 321462 95140 321468 95152
rect 321520 95140 321526 95192
rect 202230 95072 202236 95124
rect 202288 95112 202294 95124
rect 321830 95112 321836 95124
rect 202288 95084 321836 95112
rect 202288 95072 202294 95084
rect 321830 95072 321836 95084
rect 321888 95072 321894 95124
rect 204898 95004 204904 95056
rect 204956 95044 204962 95056
rect 321738 95044 321744 95056
rect 204956 95016 321744 95044
rect 204956 95004 204962 95016
rect 321738 95004 321744 95016
rect 321796 95004 321802 95056
rect 294690 94936 294696 94988
rect 294748 94976 294754 94988
rect 324682 94976 324688 94988
rect 294748 94948 324688 94976
rect 294748 94936 294754 94948
rect 324682 94936 324688 94948
rect 324740 94936 324746 94988
rect 308490 94868 308496 94920
rect 308548 94908 308554 94920
rect 324498 94908 324504 94920
rect 308548 94880 324504 94908
rect 308548 94868 308554 94880
rect 324498 94868 324504 94880
rect 324556 94868 324562 94920
rect 161474 94528 161480 94580
rect 161532 94568 161538 94580
rect 207842 94568 207848 94580
rect 161532 94540 207848 94568
rect 161532 94528 161538 94540
rect 207842 94528 207848 94540
rect 207900 94528 207906 94580
rect 130378 94460 130384 94512
rect 130436 94500 130442 94512
rect 214006 94500 214012 94512
rect 130436 94472 214012 94500
rect 130436 94460 130442 94472
rect 214006 94460 214012 94472
rect 214064 94460 214070 94512
rect 289078 94460 289084 94512
rect 289136 94500 289142 94512
rect 324314 94500 324320 94512
rect 289136 94472 324320 94500
rect 289136 94460 289142 94472
rect 324314 94460 324320 94472
rect 324372 94500 324378 94512
rect 426526 94500 426532 94512
rect 324372 94472 426532 94500
rect 324372 94460 324378 94472
rect 426526 94460 426532 94472
rect 426584 94460 426590 94512
rect 125410 93984 125416 94036
rect 125468 94024 125474 94036
rect 169110 94024 169116 94036
rect 125468 93996 169116 94024
rect 125468 93984 125474 93996
rect 169110 93984 169116 93996
rect 169168 93984 169174 94036
rect 112346 93916 112352 93968
rect 112404 93956 112410 93968
rect 178862 93956 178868 93968
rect 112404 93928 178868 93956
rect 112404 93916 112410 93928
rect 178862 93916 178868 93928
rect 178920 93916 178926 93968
rect 85574 93848 85580 93900
rect 85632 93888 85638 93900
rect 165246 93888 165252 93900
rect 85632 93860 165252 93888
rect 85632 93848 85638 93860
rect 165246 93848 165252 93860
rect 165304 93848 165310 93900
rect 67358 93780 67364 93832
rect 67416 93820 67422 93832
rect 214834 93820 214840 93832
rect 67416 93792 214840 93820
rect 67416 93780 67422 93792
rect 214834 93780 214840 93792
rect 214892 93780 214898 93832
rect 278038 93780 278044 93832
rect 278096 93820 278102 93832
rect 323578 93820 323584 93832
rect 278096 93792 323584 93820
rect 278096 93780 278102 93792
rect 323578 93780 323584 93792
rect 323636 93780 323642 93832
rect 198918 93712 198924 93764
rect 198976 93752 198982 93764
rect 324590 93752 324596 93764
rect 198976 93724 324596 93752
rect 198976 93712 198982 93724
rect 324590 93712 324596 93724
rect 324648 93712 324654 93764
rect 151722 93372 151728 93424
rect 151780 93412 151786 93424
rect 173158 93412 173164 93424
rect 151780 93384 173164 93412
rect 151780 93372 151786 93384
rect 173158 93372 173164 93384
rect 173216 93372 173222 93424
rect 118234 93304 118240 93356
rect 118292 93344 118298 93356
rect 166442 93344 166448 93356
rect 118292 93316 166448 93344
rect 118292 93304 118298 93316
rect 166442 93304 166448 93316
rect 166500 93304 166506 93356
rect 133138 93236 133144 93288
rect 133196 93276 133202 93288
rect 200850 93276 200856 93288
rect 133196 93248 200856 93276
rect 133196 93236 133202 93248
rect 200850 93236 200856 93248
rect 200908 93236 200914 93288
rect 129458 93168 129464 93220
rect 129516 93208 129522 93220
rect 198090 93208 198096 93220
rect 129516 93180 198096 93208
rect 129516 93168 129522 93180
rect 198090 93168 198096 93180
rect 198148 93168 198154 93220
rect 320818 93168 320824 93220
rect 320876 93208 320882 93220
rect 420178 93208 420184 93220
rect 320876 93180 420184 93208
rect 320876 93168 320882 93180
rect 420178 93168 420184 93180
rect 420236 93168 420242 93220
rect 98546 93100 98552 93152
rect 98604 93140 98610 93152
rect 176194 93140 176200 93152
rect 98604 93112 176200 93140
rect 98604 93100 98610 93112
rect 176194 93100 176200 93112
rect 176252 93100 176258 93152
rect 182910 93100 182916 93152
rect 182968 93140 182974 93152
rect 262950 93140 262956 93152
rect 182968 93112 262956 93140
rect 182968 93100 182974 93112
rect 262950 93100 262956 93112
rect 263008 93100 263014 93152
rect 419258 93100 419264 93152
rect 419316 93140 419322 93152
rect 580258 93140 580264 93152
rect 419316 93112 580264 93140
rect 419316 93100 419322 93112
rect 580258 93100 580264 93112
rect 580316 93100 580322 93152
rect 322934 93032 322940 93084
rect 322992 93072 322998 93084
rect 323578 93072 323584 93084
rect 322992 93044 323584 93072
rect 322992 93032 322998 93044
rect 323578 93032 323584 93044
rect 323636 93032 323642 93084
rect 110138 92420 110144 92472
rect 110196 92460 110202 92472
rect 203610 92460 203616 92472
rect 110196 92432 203616 92460
rect 110196 92420 110202 92432
rect 203610 92420 203616 92432
rect 203668 92420 203674 92472
rect 216122 92420 216128 92472
rect 216180 92460 216186 92472
rect 497090 92460 497096 92472
rect 216180 92432 497096 92460
rect 216180 92420 216186 92432
rect 497090 92420 497096 92432
rect 497148 92420 497154 92472
rect 120350 92352 120356 92404
rect 120408 92392 120414 92404
rect 211890 92392 211896 92404
rect 120408 92364 211896 92392
rect 120408 92352 120414 92364
rect 211890 92352 211896 92364
rect 211948 92352 211954 92404
rect 115474 92284 115480 92336
rect 115532 92324 115538 92336
rect 202414 92324 202420 92336
rect 115532 92296 202420 92324
rect 115532 92284 115538 92296
rect 202414 92284 202420 92296
rect 202472 92284 202478 92336
rect 88978 92216 88984 92268
rect 89036 92256 89042 92268
rect 169294 92256 169300 92268
rect 89036 92228 169300 92256
rect 89036 92216 89042 92228
rect 169294 92216 169300 92228
rect 169352 92216 169358 92268
rect 86770 92148 86776 92200
rect 86828 92188 86834 92200
rect 130378 92188 130384 92200
rect 86828 92160 130384 92188
rect 86828 92148 86834 92160
rect 130378 92148 130384 92160
rect 130436 92148 130442 92200
rect 130746 92148 130752 92200
rect 130804 92188 130810 92200
rect 174630 92188 174636 92200
rect 130804 92160 174636 92188
rect 130804 92148 130810 92160
rect 174630 92148 174636 92160
rect 174688 92148 174694 92200
rect 136082 92080 136088 92132
rect 136140 92120 136146 92132
rect 168282 92120 168288 92132
rect 136140 92092 168288 92120
rect 136140 92080 136146 92092
rect 168282 92080 168288 92092
rect 168340 92080 168346 92132
rect 85114 91060 85120 91112
rect 85172 91100 85178 91112
rect 120718 91100 120724 91112
rect 85172 91072 120724 91100
rect 85172 91060 85178 91072
rect 120718 91060 120724 91072
rect 120776 91060 120782 91112
rect 56502 90992 56508 91044
rect 56560 91032 56566 91044
rect 211982 91032 211988 91044
rect 56560 91004 211988 91032
rect 56560 90992 56566 91004
rect 211982 90992 211988 91004
rect 212040 90992 212046 91044
rect 114370 90924 114376 90976
rect 114428 90964 114434 90976
rect 196710 90964 196716 90976
rect 114428 90936 196716 90964
rect 114428 90924 114434 90936
rect 196710 90924 196716 90936
rect 196768 90924 196774 90976
rect 107746 90856 107752 90908
rect 107804 90896 107810 90908
rect 161474 90896 161480 90908
rect 107804 90868 161480 90896
rect 107804 90856 107810 90868
rect 161474 90856 161480 90868
rect 161532 90856 161538 90908
rect 122098 90788 122104 90840
rect 122156 90828 122162 90840
rect 170490 90828 170496 90840
rect 122156 90800 170496 90828
rect 122156 90788 122162 90800
rect 170490 90788 170496 90800
rect 170548 90788 170554 90840
rect 151630 90720 151636 90772
rect 151688 90760 151694 90772
rect 199378 90760 199384 90772
rect 151688 90732 199384 90760
rect 151688 90720 151694 90732
rect 199378 90720 199384 90732
rect 199436 90720 199442 90772
rect 135162 90652 135168 90704
rect 135220 90692 135226 90704
rect 171778 90692 171784 90704
rect 135220 90664 171784 90692
rect 135220 90652 135226 90664
rect 171778 90652 171784 90664
rect 171836 90652 171842 90704
rect 189810 90312 189816 90364
rect 189868 90352 189874 90364
rect 321554 90352 321560 90364
rect 189868 90324 321560 90352
rect 189868 90312 189874 90324
rect 321554 90312 321560 90324
rect 321612 90352 321618 90364
rect 465074 90352 465080 90364
rect 321612 90324 465080 90352
rect 321612 90312 321618 90324
rect 465074 90312 465080 90324
rect 465132 90312 465138 90364
rect 90542 89632 90548 89684
rect 90600 89672 90606 89684
rect 172054 89672 172060 89684
rect 90600 89644 172060 89672
rect 90600 89632 90606 89644
rect 172054 89632 172060 89644
rect 172112 89632 172118 89684
rect 249150 89632 249156 89684
rect 249208 89672 249214 89684
rect 256694 89672 256700 89684
rect 249208 89644 256700 89672
rect 249208 89632 249214 89644
rect 256694 89632 256700 89644
rect 256752 89672 256758 89684
rect 420914 89672 420920 89684
rect 256752 89644 420920 89672
rect 256752 89632 256758 89644
rect 420914 89632 420920 89644
rect 420972 89632 420978 89684
rect 95050 89564 95056 89616
rect 95108 89604 95114 89616
rect 169202 89604 169208 89616
rect 95108 89576 169208 89604
rect 95108 89564 95114 89576
rect 169202 89564 169208 89576
rect 169260 89564 169266 89616
rect 103330 89496 103336 89548
rect 103388 89536 103394 89548
rect 173342 89536 173348 89548
rect 103388 89508 173348 89536
rect 103388 89496 103394 89508
rect 173342 89496 173348 89508
rect 173400 89496 173406 89548
rect 126514 89428 126520 89480
rect 126572 89468 126578 89480
rect 192478 89468 192484 89480
rect 126572 89440 192484 89468
rect 126572 89428 126578 89440
rect 192478 89428 192484 89440
rect 192536 89428 192542 89480
rect 122834 89360 122840 89412
rect 122892 89400 122898 89412
rect 180334 89400 180340 89412
rect 122892 89372 180340 89400
rect 122892 89360 122898 89372
rect 180334 89360 180340 89372
rect 180392 89360 180398 89412
rect 153010 89292 153016 89344
rect 153068 89332 153074 89344
rect 206370 89332 206376 89344
rect 153068 89304 206376 89332
rect 153068 89292 153074 89304
rect 206370 89292 206376 89304
rect 206428 89292 206434 89344
rect 280798 89020 280804 89072
rect 280856 89060 280862 89072
rect 311894 89060 311900 89072
rect 280856 89032 311900 89060
rect 280856 89020 280862 89032
rect 311894 89020 311900 89032
rect 311952 89060 311958 89072
rect 352650 89060 352656 89072
rect 311952 89032 352656 89060
rect 311952 89020 311958 89032
rect 352650 89020 352656 89032
rect 352708 89020 352714 89072
rect 171778 88952 171784 89004
rect 171836 88992 171842 89004
rect 307294 88992 307300 89004
rect 171836 88964 307300 88992
rect 171836 88952 171842 88964
rect 307294 88952 307300 88964
rect 307352 88952 307358 89004
rect 352558 88952 352564 89004
rect 352616 88992 352622 89004
rect 462314 88992 462320 89004
rect 352616 88964 462320 88992
rect 352616 88952 352622 88964
rect 462314 88952 462320 88964
rect 462372 88952 462378 89004
rect 100570 88272 100576 88324
rect 100628 88312 100634 88324
rect 205174 88312 205180 88324
rect 100628 88284 205180 88312
rect 100628 88272 100634 88284
rect 205174 88272 205180 88284
rect 205232 88272 205238 88324
rect 104434 88204 104440 88256
rect 104492 88244 104498 88256
rect 200942 88244 200948 88256
rect 104492 88216 200948 88244
rect 104492 88204 104498 88216
rect 200942 88204 200948 88216
rect 201000 88204 201006 88256
rect 124766 88136 124772 88188
rect 124824 88176 124830 88188
rect 204990 88176 204996 88188
rect 124824 88148 204996 88176
rect 124824 88136 124830 88148
rect 204990 88136 204996 88148
rect 205048 88136 205054 88188
rect 107286 88068 107292 88120
rect 107344 88108 107350 88120
rect 171962 88108 171968 88120
rect 107344 88080 171968 88108
rect 107344 88068 107350 88080
rect 171962 88068 171968 88080
rect 172020 88068 172026 88120
rect 151446 88000 151452 88052
rect 151504 88040 151510 88052
rect 213362 88040 213368 88052
rect 151504 88012 213368 88040
rect 151504 88000 151510 88012
rect 213362 88000 213368 88012
rect 213420 88000 213426 88052
rect 114922 87932 114928 87984
rect 114980 87972 114986 87984
rect 170582 87972 170588 87984
rect 114980 87944 170588 87972
rect 114980 87932 114986 87944
rect 170582 87932 170588 87944
rect 170640 87932 170646 87984
rect 175918 87660 175924 87712
rect 175976 87700 175982 87712
rect 257430 87700 257436 87712
rect 175976 87672 257436 87700
rect 175976 87660 175982 87672
rect 257430 87660 257436 87672
rect 257488 87660 257494 87712
rect 242158 87592 242164 87644
rect 242216 87632 242222 87644
rect 347038 87632 347044 87644
rect 242216 87604 347044 87632
rect 242216 87592 242222 87604
rect 347038 87592 347044 87604
rect 347096 87592 347102 87644
rect 354030 87592 354036 87644
rect 354088 87632 354094 87644
rect 456794 87632 456800 87644
rect 354088 87604 456800 87632
rect 354088 87592 354094 87604
rect 456794 87592 456800 87604
rect 456852 87592 456858 87644
rect 75362 86912 75368 86964
rect 75420 86952 75426 86964
rect 214742 86952 214748 86964
rect 75420 86924 214748 86952
rect 75420 86912 75426 86924
rect 214742 86912 214748 86924
rect 214800 86912 214806 86964
rect 358170 86912 358176 86964
rect 358228 86952 358234 86964
rect 421558 86952 421564 86964
rect 358228 86924 421564 86952
rect 358228 86912 358234 86924
rect 421558 86912 421564 86924
rect 421616 86912 421622 86964
rect 504358 86912 504364 86964
rect 504416 86952 504422 86964
rect 580166 86952 580172 86964
rect 504416 86924 580172 86952
rect 504416 86912 504422 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 105538 86844 105544 86896
rect 105596 86884 105602 86896
rect 216674 86884 216680 86896
rect 105596 86856 216680 86884
rect 105596 86844 105602 86856
rect 216674 86844 216680 86856
rect 216732 86844 216738 86896
rect 106090 86776 106096 86828
rect 106148 86816 106154 86828
rect 202322 86816 202328 86828
rect 106148 86788 202328 86816
rect 106148 86776 106154 86788
rect 202322 86776 202328 86788
rect 202380 86776 202386 86828
rect 100202 86708 100208 86760
rect 100260 86748 100266 86760
rect 166534 86748 166540 86760
rect 100260 86720 166540 86748
rect 100260 86708 100266 86720
rect 166534 86708 166540 86720
rect 166592 86708 166598 86760
rect 123294 86640 123300 86692
rect 123352 86680 123358 86692
rect 178770 86680 178776 86692
rect 123352 86652 178776 86680
rect 123352 86640 123358 86652
rect 178770 86640 178776 86652
rect 178828 86640 178834 86692
rect 115842 86572 115848 86624
rect 115900 86612 115906 86624
rect 169018 86612 169024 86624
rect 115900 86584 169024 86612
rect 115900 86572 115906 86584
rect 169018 86572 169024 86584
rect 169076 86572 169082 86624
rect 342254 86368 342260 86420
rect 342312 86408 342318 86420
rect 357526 86408 357532 86420
rect 342312 86380 357532 86408
rect 342312 86368 342318 86380
rect 357526 86368 357532 86380
rect 357584 86408 357590 86420
rect 358170 86408 358176 86420
rect 357584 86380 358176 86408
rect 357584 86368 357590 86380
rect 358170 86368 358176 86380
rect 358228 86368 358234 86420
rect 177298 86300 177304 86352
rect 177356 86340 177362 86352
rect 253290 86340 253296 86352
rect 177356 86312 253296 86340
rect 177356 86300 177362 86312
rect 253290 86300 253296 86312
rect 253348 86300 253354 86352
rect 308398 86300 308404 86352
rect 308456 86340 308462 86352
rect 345658 86340 345664 86352
rect 308456 86312 345664 86340
rect 308456 86300 308462 86312
rect 345658 86300 345664 86312
rect 345716 86300 345722 86352
rect 209130 86232 209136 86284
rect 209188 86272 209194 86284
rect 244274 86272 244280 86284
rect 209188 86244 244280 86272
rect 209188 86232 209194 86244
rect 244274 86232 244280 86244
rect 244332 86272 244338 86284
rect 342990 86272 342996 86284
rect 244332 86244 342996 86272
rect 244332 86232 244338 86244
rect 342990 86232 342996 86244
rect 343048 86232 343054 86284
rect 377398 86232 377404 86284
rect 377456 86272 377462 86284
rect 455414 86272 455420 86284
rect 377456 86244 455420 86272
rect 377456 86232 377462 86244
rect 455414 86232 455420 86244
rect 455472 86232 455478 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 32398 85524 32404 85536
rect 3200 85496 32404 85524
rect 3200 85484 3206 85496
rect 32398 85484 32404 85496
rect 32456 85484 32462 85536
rect 88058 85484 88064 85536
rect 88116 85524 88122 85536
rect 167730 85524 167736 85536
rect 88116 85496 167736 85524
rect 88116 85484 88122 85496
rect 167730 85484 167736 85496
rect 167788 85484 167794 85536
rect 127618 85416 127624 85468
rect 127676 85456 127682 85468
rect 206462 85456 206468 85468
rect 127676 85428 206468 85456
rect 127676 85416 127682 85428
rect 206462 85416 206468 85428
rect 206520 85416 206526 85468
rect 120626 85348 120632 85400
rect 120684 85388 120690 85400
rect 196802 85388 196808 85400
rect 120684 85360 196808 85388
rect 120684 85348 120690 85360
rect 196802 85348 196808 85360
rect 196860 85348 196866 85400
rect 101858 85280 101864 85332
rect 101916 85320 101922 85332
rect 174722 85320 174728 85332
rect 101916 85292 174728 85320
rect 101916 85280 101922 85292
rect 174722 85280 174728 85292
rect 174780 85280 174786 85332
rect 111242 85212 111248 85264
rect 111300 85252 111306 85264
rect 173434 85252 173440 85264
rect 111300 85224 173440 85252
rect 111300 85212 111306 85224
rect 173434 85212 173440 85224
rect 173492 85212 173498 85264
rect 195330 84872 195336 84924
rect 195388 84912 195394 84924
rect 266354 84912 266360 84924
rect 195388 84884 266360 84912
rect 195388 84872 195394 84884
rect 266354 84872 266360 84884
rect 266412 84872 266418 84924
rect 195422 84804 195428 84856
rect 195480 84844 195486 84856
rect 307202 84844 307208 84856
rect 195480 84816 307208 84844
rect 195480 84804 195486 84816
rect 307202 84804 307208 84816
rect 307260 84804 307266 84856
rect 316034 84804 316040 84856
rect 316092 84844 316098 84856
rect 333238 84844 333244 84856
rect 316092 84816 333244 84844
rect 316092 84804 316098 84816
rect 333238 84804 333244 84816
rect 333296 84804 333302 84856
rect 336090 84804 336096 84856
rect 336148 84844 336154 84856
rect 460934 84844 460940 84856
rect 336148 84816 460940 84844
rect 336148 84804 336154 84816
rect 460934 84804 460940 84816
rect 460992 84804 460998 84856
rect 65978 84124 65984 84176
rect 66036 84164 66042 84176
rect 214650 84164 214656 84176
rect 66036 84136 214656 84164
rect 66036 84124 66042 84136
rect 214650 84124 214656 84136
rect 214708 84124 214714 84176
rect 291838 84124 291844 84176
rect 291896 84164 291902 84176
rect 332042 84164 332048 84176
rect 291896 84136 332048 84164
rect 291896 84124 291902 84136
rect 332042 84124 332048 84136
rect 332100 84124 332106 84176
rect 103422 84056 103428 84108
rect 103480 84096 103486 84108
rect 196894 84096 196900 84108
rect 103480 84068 196900 84096
rect 103480 84056 103486 84068
rect 196894 84056 196900 84068
rect 196952 84056 196958 84108
rect 96522 83988 96528 84040
rect 96580 84028 96586 84040
rect 174814 84028 174820 84040
rect 96580 84000 174820 84028
rect 96580 83988 96586 84000
rect 174814 83988 174820 84000
rect 174872 83988 174878 84040
rect 92382 83920 92388 83972
rect 92440 83960 92446 83972
rect 170674 83960 170680 83972
rect 92440 83932 170680 83960
rect 92440 83920 92446 83932
rect 170674 83920 170680 83932
rect 170732 83920 170738 83972
rect 117130 83852 117136 83904
rect 117188 83892 117194 83904
rect 181530 83892 181536 83904
rect 117188 83864 181536 83892
rect 117188 83852 117194 83864
rect 181530 83852 181536 83864
rect 181588 83852 181594 83904
rect 132402 83784 132408 83836
rect 132460 83824 132466 83836
rect 166258 83824 166264 83836
rect 132460 83796 166264 83824
rect 132460 83784 132466 83796
rect 166258 83784 166264 83796
rect 166316 83784 166322 83836
rect 185670 83444 185676 83496
rect 185728 83484 185734 83496
rect 254762 83484 254768 83496
rect 185728 83456 254768 83484
rect 185728 83444 185734 83456
rect 254762 83444 254768 83456
rect 254820 83444 254826 83496
rect 331950 83444 331956 83496
rect 332008 83484 332014 83496
rect 463694 83484 463700 83496
rect 332008 83456 463700 83484
rect 332008 83444 332014 83456
rect 463694 83444 463700 83456
rect 463752 83444 463758 83496
rect 291194 82832 291200 82884
rect 291252 82872 291258 82884
rect 291838 82872 291844 82884
rect 291252 82844 291844 82872
rect 291252 82832 291258 82844
rect 291838 82832 291844 82844
rect 291896 82832 291902 82884
rect 108942 82764 108948 82816
rect 109000 82804 109006 82816
rect 210510 82804 210516 82816
rect 109000 82776 210516 82804
rect 109000 82764 109006 82776
rect 210510 82764 210516 82776
rect 210568 82764 210574 82816
rect 107562 82696 107568 82748
rect 107620 82736 107626 82748
rect 195514 82736 195520 82748
rect 107620 82708 195520 82736
rect 107620 82696 107626 82708
rect 195514 82696 195520 82708
rect 195572 82696 195578 82748
rect 101950 82628 101956 82680
rect 102008 82668 102014 82680
rect 176010 82668 176016 82680
rect 102008 82640 176016 82668
rect 102008 82628 102014 82640
rect 176010 82628 176016 82640
rect 176068 82628 176074 82680
rect 117222 82560 117228 82612
rect 117280 82600 117286 82612
rect 183002 82600 183008 82612
rect 117280 82572 183008 82600
rect 117280 82560 117286 82572
rect 183002 82560 183008 82572
rect 183060 82560 183066 82612
rect 119890 82492 119896 82544
rect 119948 82532 119954 82544
rect 170398 82532 170404 82544
rect 119948 82504 170404 82532
rect 119948 82492 119954 82504
rect 170398 82492 170404 82504
rect 170456 82492 170462 82544
rect 122742 82424 122748 82476
rect 122800 82464 122806 82476
rect 166350 82464 166356 82476
rect 122800 82436 166356 82464
rect 122800 82424 122806 82436
rect 166350 82424 166356 82436
rect 166408 82424 166414 82476
rect 238018 82084 238024 82136
rect 238076 82124 238082 82136
rect 251174 82124 251180 82136
rect 238076 82096 251180 82124
rect 238076 82084 238082 82096
rect 251174 82084 251180 82096
rect 251232 82084 251238 82136
rect 324958 82084 324964 82136
rect 325016 82124 325022 82136
rect 461578 82124 461584 82136
rect 325016 82096 461584 82124
rect 325016 82084 325022 82096
rect 461578 82084 461584 82096
rect 461636 82084 461642 82136
rect 99190 81336 99196 81388
rect 99248 81376 99254 81388
rect 184382 81376 184388 81388
rect 99248 81348 184388 81376
rect 99248 81336 99254 81348
rect 184382 81336 184388 81348
rect 184440 81336 184446 81388
rect 345750 81336 345756 81388
rect 345808 81376 345814 81388
rect 465718 81376 465724 81388
rect 345808 81348 465724 81376
rect 345808 81336 345814 81348
rect 465718 81336 465724 81348
rect 465776 81336 465782 81388
rect 119982 81268 119988 81320
rect 120040 81308 120046 81320
rect 203518 81308 203524 81320
rect 120040 81280 203524 81308
rect 120040 81268 120046 81280
rect 203518 81268 203524 81280
rect 203576 81268 203582 81320
rect 110230 81200 110236 81252
rect 110288 81240 110294 81252
rect 181622 81240 181628 81252
rect 110288 81212 181628 81240
rect 110288 81200 110294 81212
rect 181622 81200 181628 81212
rect 181680 81200 181686 81252
rect 97810 81132 97816 81184
rect 97868 81172 97874 81184
rect 167822 81172 167828 81184
rect 97868 81144 167828 81172
rect 97868 81132 97874 81144
rect 167822 81132 167828 81144
rect 167880 81132 167886 81184
rect 184198 80656 184204 80708
rect 184256 80696 184262 80708
rect 313918 80696 313924 80708
rect 184256 80668 313924 80696
rect 184256 80656 184262 80668
rect 313918 80656 313924 80668
rect 313976 80656 313982 80708
rect 317414 80044 317420 80096
rect 317472 80084 317478 80096
rect 345750 80084 345756 80096
rect 317472 80056 345756 80084
rect 317472 80044 317478 80056
rect 345750 80044 345756 80056
rect 345808 80044 345814 80096
rect 68278 79976 68284 80028
rect 68336 80016 68342 80028
rect 199470 80016 199476 80028
rect 68336 79988 199476 80016
rect 68336 79976 68342 79988
rect 199470 79976 199476 79988
rect 199528 79976 199534 80028
rect 93762 79908 93768 79960
rect 93820 79948 93826 79960
rect 176102 79948 176108 79960
rect 93820 79920 176108 79948
rect 93820 79908 93826 79920
rect 176102 79908 176108 79920
rect 176160 79908 176166 79960
rect 126882 79840 126888 79892
rect 126940 79880 126946 79892
rect 209222 79880 209228 79892
rect 126940 79852 209228 79880
rect 126940 79840 126946 79852
rect 209222 79840 209228 79852
rect 209280 79840 209286 79892
rect 102042 79772 102048 79824
rect 102100 79812 102106 79824
rect 177482 79812 177488 79824
rect 102100 79784 177488 79812
rect 102100 79772 102106 79784
rect 177482 79772 177488 79784
rect 177540 79772 177546 79824
rect 97902 79704 97908 79756
rect 97960 79744 97966 79756
rect 173250 79744 173256 79756
rect 97960 79716 173256 79744
rect 97960 79704 97966 79716
rect 173250 79704 173256 79716
rect 173308 79704 173314 79756
rect 195238 79364 195244 79416
rect 195296 79404 195302 79416
rect 232498 79404 232504 79416
rect 195296 79376 232504 79404
rect 195296 79364 195302 79376
rect 232498 79364 232504 79376
rect 232556 79364 232562 79416
rect 200758 79296 200764 79348
rect 200816 79336 200822 79348
rect 246298 79336 246304 79348
rect 200816 79308 246304 79336
rect 200816 79296 200822 79308
rect 246298 79296 246304 79308
rect 246356 79296 246362 79348
rect 309778 79296 309784 79348
rect 309836 79336 309842 79348
rect 470594 79336 470600 79348
rect 309836 79308 470600 79336
rect 309836 79296 309842 79308
rect 470594 79296 470600 79308
rect 470652 79296 470658 79348
rect 114462 78616 114468 78668
rect 114520 78656 114526 78668
rect 213454 78656 213460 78668
rect 114520 78628 213460 78656
rect 114520 78616 114526 78628
rect 213454 78616 213460 78628
rect 213512 78616 213518 78668
rect 266354 78616 266360 78668
rect 266412 78656 266418 78668
rect 338758 78656 338764 78668
rect 266412 78628 338764 78656
rect 266412 78616 266418 78628
rect 338758 78616 338764 78628
rect 338816 78616 338822 78668
rect 339126 78616 339132 78668
rect 339184 78656 339190 78668
rect 471974 78656 471980 78668
rect 339184 78628 471980 78656
rect 339184 78616 339190 78628
rect 471974 78616 471980 78628
rect 472032 78616 472038 78668
rect 95142 78548 95148 78600
rect 95200 78588 95206 78600
rect 180426 78588 180432 78600
rect 95200 78560 180432 78588
rect 95200 78548 95206 78560
rect 180426 78548 180432 78560
rect 180484 78548 180490 78600
rect 110322 78480 110328 78532
rect 110380 78520 110386 78532
rect 177390 78520 177396 78532
rect 110380 78492 177396 78520
rect 110380 78480 110386 78492
rect 177390 78480 177396 78492
rect 177448 78480 177454 78532
rect 188430 78004 188436 78056
rect 188488 78044 188494 78056
rect 286502 78044 286508 78056
rect 188488 78016 286508 78044
rect 188488 78004 188494 78016
rect 286502 78004 286508 78016
rect 286560 78004 286566 78056
rect 42702 77936 42708 77988
rect 42760 77976 42766 77988
rect 128354 77976 128360 77988
rect 42760 77948 128360 77976
rect 42760 77936 42766 77948
rect 128354 77936 128360 77948
rect 128412 77936 128418 77988
rect 180150 77936 180156 77988
rect 180208 77976 180214 77988
rect 278222 77976 278228 77988
rect 180208 77948 278228 77976
rect 180208 77936 180214 77948
rect 278222 77936 278228 77948
rect 278280 77936 278286 77988
rect 120718 77188 120724 77240
rect 120776 77228 120782 77240
rect 205082 77228 205088 77240
rect 120776 77200 205088 77228
rect 120776 77188 120782 77200
rect 205082 77188 205088 77200
rect 205140 77188 205146 77240
rect 123938 77120 123944 77172
rect 123996 77160 124002 77172
rect 171870 77160 171876 77172
rect 123996 77132 171876 77160
rect 123996 77120 124002 77132
rect 171870 77120 171876 77132
rect 171928 77120 171934 77172
rect 102134 76508 102140 76560
rect 102192 76548 102198 76560
rect 305914 76548 305920 76560
rect 102192 76520 305920 76548
rect 102192 76508 102198 76520
rect 305914 76508 305920 76520
rect 305972 76508 305978 76560
rect 307202 76508 307208 76560
rect 307260 76548 307266 76560
rect 473354 76548 473360 76560
rect 307260 76520 473360 76548
rect 307260 76508 307266 76520
rect 473354 76508 473360 76520
rect 473412 76508 473418 76560
rect 93854 75216 93860 75268
rect 93912 75256 93918 75268
rect 297450 75256 297456 75268
rect 93912 75228 297456 75256
rect 93912 75216 93918 75228
rect 297450 75216 297456 75228
rect 297508 75216 297514 75268
rect 53834 75148 53840 75200
rect 53892 75188 53898 75200
rect 267182 75188 267188 75200
rect 53892 75160 267188 75188
rect 53892 75148 53898 75160
rect 267182 75148 267188 75160
rect 267240 75148 267246 75200
rect 297634 75148 297640 75200
rect 297692 75188 297698 75200
rect 472618 75188 472624 75200
rect 297692 75160 472624 75188
rect 297692 75148 297698 75160
rect 472618 75148 472624 75160
rect 472676 75148 472682 75200
rect 57882 74468 57888 74520
rect 57940 74508 57946 74520
rect 207750 74508 207756 74520
rect 57940 74480 207756 74508
rect 57940 74468 57946 74480
rect 207750 74468 207756 74480
rect 207808 74468 207814 74520
rect 86954 73856 86960 73908
rect 87012 73896 87018 73908
rect 269850 73896 269856 73908
rect 87012 73868 269856 73896
rect 87012 73856 87018 73868
rect 269850 73856 269856 73868
rect 269908 73856 269914 73908
rect 121454 73788 121460 73840
rect 121512 73828 121518 73840
rect 309134 73828 309140 73840
rect 121512 73800 309140 73828
rect 121512 73788 121518 73800
rect 309134 73788 309140 73800
rect 309192 73788 309198 73840
rect 311158 73788 311164 73840
rect 311216 73828 311222 73840
rect 469214 73828 469220 73840
rect 311216 73800 469220 73828
rect 311216 73788 311222 73800
rect 469214 73788 469220 73800
rect 469272 73788 469278 73840
rect 64598 73108 64604 73160
rect 64656 73148 64662 73160
rect 320818 73148 320824 73160
rect 64656 73120 320824 73148
rect 64656 73108 64662 73120
rect 320818 73108 320824 73120
rect 320876 73108 320882 73160
rect 419442 73108 419448 73160
rect 419500 73148 419506 73160
rect 579982 73148 579988 73160
rect 419500 73120 579988 73148
rect 419500 73108 419506 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 262950 73040 262956 73092
rect 263008 73080 263014 73092
rect 414658 73080 414664 73092
rect 263008 73052 414664 73080
rect 263008 73040 263014 73052
rect 414658 73040 414664 73052
rect 414716 73040 414722 73092
rect 107654 72496 107660 72548
rect 107712 72536 107718 72548
rect 253382 72536 253388 72548
rect 107712 72508 253388 72536
rect 107712 72496 107718 72508
rect 253382 72496 253388 72508
rect 253440 72496 253446 72548
rect 60734 72428 60740 72480
rect 60792 72468 60798 72480
rect 290550 72468 290556 72480
rect 60792 72440 290556 72468
rect 60792 72428 60798 72440
rect 290550 72428 290556 72440
rect 290608 72428 290614 72480
rect 262214 71748 262220 71800
rect 262272 71788 262278 71800
rect 262950 71788 262956 71800
rect 262272 71760 262956 71788
rect 262272 71748 262278 71760
rect 262950 71748 262956 71760
rect 263008 71748 263014 71800
rect 320174 71748 320180 71800
rect 320232 71788 320238 71800
rect 320818 71788 320824 71800
rect 320232 71760 320824 71788
rect 320232 71748 320238 71760
rect 320818 71748 320824 71760
rect 320876 71748 320882 71800
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 41322 71720 41328 71732
rect 3476 71692 41328 71720
rect 3476 71680 3482 71692
rect 41322 71680 41328 71692
rect 41380 71720 41386 71732
rect 494146 71720 494152 71732
rect 41380 71692 494152 71720
rect 41380 71680 41386 71692
rect 494146 71680 494152 71692
rect 494204 71680 494210 71732
rect 80054 71068 80060 71120
rect 80112 71108 80118 71120
rect 287882 71108 287888 71120
rect 80112 71080 287888 71108
rect 80112 71068 80118 71080
rect 287882 71068 287888 71080
rect 287940 71068 287946 71120
rect 66254 71000 66260 71052
rect 66312 71040 66318 71052
rect 278314 71040 278320 71052
rect 66312 71012 278320 71040
rect 66312 71000 66318 71012
rect 278314 71000 278320 71012
rect 278372 71000 278378 71052
rect 362954 70320 362960 70372
rect 363012 70360 363018 70372
rect 459554 70360 459560 70372
rect 363012 70332 459560 70360
rect 363012 70320 363018 70332
rect 459554 70320 459560 70332
rect 459612 70320 459618 70372
rect 178678 69776 178684 69828
rect 178736 69816 178742 69828
rect 347038 69816 347044 69828
rect 178736 69788 347044 69816
rect 178736 69776 178742 69788
rect 347038 69776 347044 69788
rect 347096 69776 347102 69828
rect 54754 69708 54760 69760
rect 54812 69748 54818 69760
rect 226978 69748 226984 69760
rect 54812 69720 226984 69748
rect 54812 69708 54818 69720
rect 226978 69708 226984 69720
rect 227036 69708 227042 69760
rect 55214 69640 55220 69692
rect 55272 69680 55278 69692
rect 304534 69680 304540 69692
rect 55272 69652 304540 69680
rect 55272 69640 55278 69652
rect 304534 69640 304540 69652
rect 304592 69640 304598 69692
rect 339494 69640 339500 69692
rect 339552 69680 339558 69692
rect 362954 69680 362960 69692
rect 339552 69652 362960 69680
rect 339552 69640 339558 69652
rect 362954 69640 362960 69652
rect 363012 69640 363018 69692
rect 60642 68960 60648 69012
rect 60700 69000 60706 69012
rect 335354 69000 335360 69012
rect 60700 68972 335360 69000
rect 60700 68960 60706 68972
rect 335354 68960 335360 68972
rect 335412 69000 335418 69012
rect 336090 69000 336096 69012
rect 335412 68972 336096 69000
rect 335412 68960 335418 68972
rect 336090 68960 336096 68972
rect 336148 68960 336154 69012
rect 104894 68348 104900 68400
rect 104952 68388 104958 68400
rect 293310 68388 293316 68400
rect 104952 68360 293316 68388
rect 104952 68348 104958 68360
rect 293310 68348 293316 68360
rect 293368 68348 293374 68400
rect 52362 68280 52368 68332
rect 52420 68320 52426 68332
rect 246390 68320 246396 68332
rect 52420 68292 246396 68320
rect 52420 68280 52426 68292
rect 246390 68280 246396 68292
rect 246448 68280 246454 68332
rect 286318 68280 286324 68332
rect 286376 68320 286382 68332
rect 292574 68320 292580 68332
rect 286376 68292 292580 68320
rect 286376 68280 286382 68292
rect 292574 68280 292580 68292
rect 292632 68320 292638 68332
rect 474734 68320 474740 68332
rect 292632 68292 474740 68320
rect 292632 68280 292638 68292
rect 474734 68280 474740 68292
rect 474792 68280 474798 68332
rect 287698 67532 287704 67584
rect 287756 67572 287762 67584
rect 289814 67572 289820 67584
rect 287756 67544 289820 67572
rect 287756 67532 287762 67544
rect 289814 67532 289820 67544
rect 289872 67532 289878 67584
rect 114554 66988 114560 67040
rect 114612 67028 114618 67040
rect 294782 67028 294788 67040
rect 114612 67000 294788 67028
rect 114612 66988 114618 67000
rect 294782 66988 294788 67000
rect 294840 66988 294846 67040
rect 289814 66920 289820 66972
rect 289872 66960 289878 66972
rect 476114 66960 476120 66972
rect 289872 66932 476120 66960
rect 289872 66920 289878 66932
rect 476114 66920 476120 66932
rect 476172 66920 476178 66972
rect 35894 66852 35900 66904
rect 35952 66892 35958 66904
rect 298830 66892 298836 66904
rect 35952 66864 298836 66892
rect 35952 66852 35958 66864
rect 298830 66852 298836 66864
rect 298888 66852 298894 66904
rect 285674 66172 285680 66224
rect 285732 66212 285738 66224
rect 286502 66212 286508 66224
rect 285732 66184 286508 66212
rect 285732 66172 285738 66184
rect 286502 66172 286508 66184
rect 286560 66212 286566 66224
rect 477494 66212 477500 66224
rect 286560 66184 477500 66212
rect 286560 66172 286566 66184
rect 477494 66172 477500 66184
rect 477552 66172 477558 66224
rect 193858 65628 193864 65680
rect 193916 65668 193922 65680
rect 332042 65668 332048 65680
rect 193916 65640 332048 65668
rect 193916 65628 193922 65640
rect 332042 65628 332048 65640
rect 332100 65628 332106 65680
rect 61654 65560 61660 65612
rect 61712 65600 61718 65612
rect 269850 65600 269856 65612
rect 61712 65572 269856 65600
rect 61712 65560 61718 65572
rect 269850 65560 269856 65572
rect 269908 65560 269914 65612
rect 40034 65492 40040 65544
rect 40092 65532 40098 65544
rect 297542 65532 297548 65544
rect 40092 65504 297548 65532
rect 40092 65492 40098 65504
rect 297542 65492 297548 65504
rect 297600 65492 297606 65544
rect 188338 64268 188344 64320
rect 188396 64308 188402 64320
rect 333238 64308 333244 64320
rect 188396 64280 333244 64308
rect 188396 64268 188402 64280
rect 333238 64268 333244 64280
rect 333296 64268 333302 64320
rect 59170 64200 59176 64252
rect 59228 64240 59234 64252
rect 274082 64240 274088 64252
rect 59228 64212 274088 64240
rect 59228 64200 59234 64212
rect 274082 64200 274088 64212
rect 274140 64200 274146 64252
rect 276658 64200 276664 64252
rect 276716 64240 276722 64252
rect 278774 64240 278780 64252
rect 276716 64212 278780 64240
rect 276716 64200 276722 64212
rect 278774 64200 278780 64212
rect 278832 64240 278838 64252
rect 480254 64240 480260 64252
rect 278832 64212 480260 64240
rect 278832 64200 278838 64212
rect 480254 64200 480260 64212
rect 480312 64200 480318 64252
rect 73154 64132 73160 64184
rect 73212 64172 73218 64184
rect 300302 64172 300308 64184
rect 73212 64144 300308 64172
rect 73212 64132 73218 64144
rect 300302 64132 300308 64144
rect 300360 64132 300366 64184
rect 97994 62840 98000 62892
rect 98052 62880 98058 62892
rect 303062 62880 303068 62892
rect 98052 62852 303068 62880
rect 98052 62840 98058 62852
rect 303062 62840 303068 62852
rect 303120 62840 303126 62892
rect 33134 62772 33140 62824
rect 33192 62812 33198 62824
rect 269942 62812 269948 62824
rect 33192 62784 269948 62812
rect 33192 62772 33198 62784
rect 269942 62772 269948 62784
rect 270000 62772 270006 62824
rect 278038 62772 278044 62824
rect 278096 62812 278102 62824
rect 481726 62812 481732 62824
rect 278096 62784 481732 62812
rect 278096 62772 278102 62784
rect 481726 62772 481732 62784
rect 481784 62772 481790 62824
rect 118694 61412 118700 61464
rect 118752 61452 118758 61464
rect 272518 61452 272524 61464
rect 118752 61424 272524 61452
rect 118752 61412 118758 61424
rect 272518 61412 272524 61424
rect 272576 61412 272582 61464
rect 273162 61344 273168 61396
rect 273220 61384 273226 61396
rect 481634 61384 481640 61396
rect 273220 61356 481640 61384
rect 273220 61344 273226 61356
rect 481634 61344 481640 61356
rect 481692 61344 481698 61396
rect 512638 60664 512644 60716
rect 512696 60704 512702 60716
rect 580166 60704 580172 60716
rect 512696 60676 580172 60704
rect 512696 60664 512702 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 52454 60052 52460 60104
rect 52512 60092 52518 60104
rect 261570 60092 261576 60104
rect 52512 60064 261576 60092
rect 52512 60052 52518 60064
rect 261570 60052 261576 60064
rect 261628 60052 261634 60104
rect 268470 60052 268476 60104
rect 268528 60092 268534 60104
rect 483014 60092 483020 60104
rect 268528 60064 483020 60092
rect 268528 60052 268534 60064
rect 483014 60052 483020 60064
rect 483072 60052 483078 60104
rect 56594 59984 56600 60036
rect 56652 60024 56658 60036
rect 278130 60024 278136 60036
rect 56652 59996 278136 60024
rect 56652 59984 56658 59996
rect 278130 59984 278136 59996
rect 278188 59984 278194 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 17218 59344 17224 59356
rect 3108 59316 17224 59344
rect 3108 59304 3114 59316
rect 17218 59304 17224 59316
rect 17276 59304 17282 59356
rect 332594 59304 332600 59356
rect 332652 59344 332658 59356
rect 400858 59344 400864 59356
rect 332652 59316 400864 59344
rect 332652 59304 332658 59316
rect 400858 59304 400864 59316
rect 400916 59304 400922 59356
rect 246390 58828 246396 58880
rect 246448 58868 246454 58880
rect 264974 58868 264980 58880
rect 246448 58840 264980 58868
rect 246448 58828 246454 58840
rect 264974 58828 264980 58840
rect 265032 58828 265038 58880
rect 84194 58760 84200 58812
rect 84252 58800 84258 58812
rect 268378 58800 268384 58812
rect 84252 58772 268384 58800
rect 84252 58760 84258 58772
rect 268378 58760 268384 58772
rect 268436 58760 268442 58812
rect 49694 58692 49700 58744
rect 49752 58732 49758 58744
rect 304442 58732 304448 58744
rect 49752 58704 304448 58732
rect 49752 58692 49758 58704
rect 304442 58692 304448 58704
rect 304500 58692 304506 58744
rect 6914 58624 6920 58676
rect 6972 58664 6978 58676
rect 264514 58664 264520 58676
rect 6972 58636 264520 58664
rect 6972 58624 6978 58636
rect 264514 58624 264520 58636
rect 264572 58624 264578 58676
rect 264974 58624 264980 58676
rect 265032 58664 265038 58676
rect 484394 58664 484400 58676
rect 265032 58636 484400 58664
rect 265032 58624 265038 58636
rect 484394 58624 484400 58636
rect 484452 58624 484458 58676
rect 261478 57876 261484 57928
rect 261536 57916 261542 57928
rect 485774 57916 485780 57928
rect 261536 57888 485780 57916
rect 261536 57876 261542 57888
rect 485774 57876 485780 57888
rect 485832 57876 485838 57928
rect 260834 57400 260840 57452
rect 260892 57440 260898 57452
rect 261478 57440 261484 57452
rect 260892 57412 261484 57440
rect 260892 57400 260898 57412
rect 261478 57400 261484 57412
rect 261536 57400 261542 57452
rect 52546 57196 52552 57248
rect 52604 57236 52610 57248
rect 261662 57236 261668 57248
rect 52604 57208 261668 57236
rect 52604 57196 52610 57208
rect 261662 57196 261668 57208
rect 261720 57196 261726 57248
rect 122834 55972 122840 56024
rect 122892 56012 122898 56024
rect 296162 56012 296168 56024
rect 122892 55984 296168 56012
rect 122892 55972 122898 55984
rect 296162 55972 296168 55984
rect 296220 55972 296226 56024
rect 46934 55904 46940 55956
rect 46992 55944 46998 55956
rect 258902 55944 258908 55956
rect 46992 55916 258908 55944
rect 46992 55904 46998 55916
rect 258902 55904 258908 55916
rect 258960 55904 258966 55956
rect 19334 55836 19340 55888
rect 19392 55876 19398 55888
rect 256050 55876 256056 55888
rect 19392 55848 256056 55876
rect 19392 55836 19398 55848
rect 256050 55836 256056 55848
rect 256108 55836 256114 55888
rect 488534 55876 488540 55888
rect 258046 55848 488540 55876
rect 254762 55768 254768 55820
rect 254820 55808 254826 55820
rect 258046 55808 258074 55848
rect 488534 55836 488540 55848
rect 488592 55836 488598 55888
rect 254820 55780 258074 55808
rect 254820 55768 254826 55780
rect 51074 54612 51080 54664
rect 51132 54652 51138 54664
rect 275370 54652 275376 54664
rect 51132 54624 275376 54652
rect 51132 54612 51138 54624
rect 275370 54612 275376 54624
rect 275428 54612 275434 54664
rect 67634 54544 67640 54596
rect 67692 54584 67698 54596
rect 297358 54584 297364 54596
rect 67692 54556 297364 54584
rect 67692 54544 67698 54556
rect 297358 54544 297364 54556
rect 297416 54544 297422 54596
rect 124214 54476 124220 54528
rect 124272 54516 124278 54528
rect 250622 54516 250628 54528
rect 124272 54488 250628 54516
rect 124272 54476 124278 54488
rect 250622 54476 250628 54488
rect 250680 54476 250686 54528
rect 251910 54476 251916 54528
rect 251968 54516 251974 54528
rect 489914 54516 489920 54528
rect 251968 54488 489920 54516
rect 251968 54476 251974 54488
rect 489914 54476 489920 54488
rect 489972 54476 489978 54528
rect 74534 53184 74540 53236
rect 74592 53224 74598 53236
rect 292022 53224 292028 53236
rect 74592 53196 292028 53224
rect 74592 53184 74598 53196
rect 292022 53184 292028 53196
rect 292080 53184 292086 53236
rect 31754 53116 31760 53168
rect 31812 53156 31818 53168
rect 264330 53156 264336 53168
rect 31812 53128 264336 53156
rect 31812 53116 31818 53128
rect 264330 53116 264336 53128
rect 264388 53116 264394 53168
rect 37182 53048 37188 53100
rect 37240 53088 37246 53100
rect 232590 53088 232596 53100
rect 37240 53060 232596 53088
rect 37240 53048 37246 53060
rect 232590 53048 232596 53060
rect 232648 53048 232654 53100
rect 247954 53048 247960 53100
rect 248012 53088 248018 53100
rect 491294 53088 491300 53100
rect 248012 53060 491300 53088
rect 248012 53048 248018 53060
rect 491294 53048 491300 53060
rect 491352 53048 491358 53100
rect 243538 51824 243544 51876
rect 243596 51864 243602 51876
rect 467098 51864 467104 51876
rect 243596 51836 467104 51864
rect 243596 51824 243602 51836
rect 467098 51824 467104 51836
rect 467156 51824 467162 51876
rect 70394 51756 70400 51808
rect 70452 51796 70458 51808
rect 300210 51796 300216 51808
rect 70452 51768 300216 51796
rect 70452 51756 70458 51768
rect 300210 51756 300216 51768
rect 300268 51756 300274 51808
rect 4154 51688 4160 51740
rect 4212 51728 4218 51740
rect 249242 51728 249248 51740
rect 4212 51700 249248 51728
rect 4212 51688 4218 51700
rect 249242 51688 249248 51700
rect 249300 51688 249306 51740
rect 196618 51008 196624 51060
rect 196676 51048 196682 51060
rect 247034 51048 247040 51060
rect 196676 51020 247040 51048
rect 196676 51008 196682 51020
rect 247034 51008 247040 51020
rect 247092 51048 247098 51060
rect 247954 51048 247960 51060
rect 247092 51020 247960 51048
rect 247092 51008 247098 51020
rect 247954 51008 247960 51020
rect 248012 51008 248018 51060
rect 71774 50464 71780 50516
rect 71832 50504 71838 50516
rect 250714 50504 250720 50516
rect 71832 50476 250720 50504
rect 71832 50464 71838 50476
rect 250714 50464 250720 50476
rect 250772 50464 250778 50516
rect 240778 50396 240784 50448
rect 240836 50436 240842 50448
rect 492674 50436 492680 50448
rect 240836 50408 492680 50436
rect 240836 50396 240842 50408
rect 492674 50396 492680 50408
rect 492732 50396 492738 50448
rect 24854 50328 24860 50380
rect 24912 50368 24918 50380
rect 298922 50368 298928 50380
rect 24912 50340 298928 50368
rect 24912 50328 24918 50340
rect 298922 50328 298928 50340
rect 298980 50328 298986 50380
rect 64690 49648 64696 49700
rect 64748 49688 64754 49700
rect 310514 49688 310520 49700
rect 64748 49660 310520 49688
rect 64748 49648 64754 49660
rect 310514 49648 310520 49660
rect 310572 49688 310578 49700
rect 311158 49688 311164 49700
rect 310572 49660 311164 49688
rect 310572 49648 310578 49660
rect 311158 49648 311164 49660
rect 311216 49648 311222 49700
rect 349154 49648 349160 49700
rect 349212 49688 349218 49700
rect 352006 49688 352012 49700
rect 349212 49660 352012 49688
rect 349212 49648 349218 49660
rect 352006 49648 352012 49660
rect 352064 49688 352070 49700
rect 494054 49688 494060 49700
rect 352064 49660 494060 49688
rect 352064 49648 352070 49660
rect 494054 49648 494060 49660
rect 494112 49648 494118 49700
rect 269114 49580 269120 49632
rect 269172 49620 269178 49632
rect 269850 49620 269856 49632
rect 269172 49592 269856 49620
rect 269172 49580 269178 49592
rect 269850 49580 269856 49592
rect 269908 49620 269914 49632
rect 359458 49620 359464 49632
rect 269908 49592 359464 49620
rect 269908 49580 269914 49592
rect 359458 49580 359464 49592
rect 359516 49580 359522 49632
rect 88334 49036 88340 49088
rect 88392 49076 88398 49088
rect 289170 49076 289176 49088
rect 88392 49048 289176 49076
rect 88392 49036 88398 49048
rect 289170 49036 289176 49048
rect 289228 49036 289234 49088
rect 37274 48968 37280 49020
rect 37332 49008 37338 49020
rect 271138 49008 271144 49020
rect 37332 48980 271144 49008
rect 37332 48968 37338 48980
rect 271138 48968 271144 48980
rect 271196 48968 271202 49020
rect 274082 48220 274088 48272
rect 274140 48260 274146 48272
rect 340138 48260 340144 48272
rect 274140 48232 340144 48260
rect 274140 48220 274146 48232
rect 340138 48220 340144 48232
rect 340196 48220 340202 48272
rect 189718 47676 189724 47728
rect 189776 47716 189782 47728
rect 315298 47716 315304 47728
rect 189776 47688 315304 47716
rect 189776 47676 189782 47688
rect 315298 47676 315304 47688
rect 315356 47676 315362 47728
rect 99374 47608 99380 47660
rect 99432 47648 99438 47660
rect 254670 47648 254676 47660
rect 99432 47620 254676 47648
rect 99432 47608 99438 47620
rect 254670 47608 254676 47620
rect 254728 47608 254734 47660
rect 110414 47540 110420 47592
rect 110472 47580 110478 47592
rect 273990 47580 273996 47592
rect 110472 47552 273996 47580
rect 110472 47540 110478 47552
rect 273990 47540 273996 47552
rect 274048 47540 274054 47592
rect 340874 47540 340880 47592
rect 340932 47580 340938 47592
rect 498194 47580 498200 47592
rect 340932 47552 498200 47580
rect 340932 47540 340938 47552
rect 498194 47540 498200 47552
rect 498252 47540 498258 47592
rect 273254 47336 273260 47388
rect 273312 47376 273318 47388
rect 274082 47376 274088 47388
rect 273312 47348 274088 47376
rect 273312 47336 273318 47348
rect 274082 47336 274088 47348
rect 274140 47336 274146 47388
rect 367830 46860 367836 46912
rect 367888 46900 367894 46912
rect 422294 46900 422300 46912
rect 367888 46872 422300 46900
rect 367888 46860 367894 46872
rect 422294 46860 422300 46872
rect 422352 46860 422358 46912
rect 525058 46860 525064 46912
rect 525116 46900 525122 46912
rect 580166 46900 580172 46912
rect 525116 46872 580172 46900
rect 525116 46860 525122 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 115934 46316 115940 46368
rect 115992 46356 115998 46368
rect 285030 46356 285036 46368
rect 115992 46328 285036 46356
rect 115992 46316 115998 46328
rect 285030 46316 285036 46328
rect 285088 46316 285094 46368
rect 15194 46248 15200 46300
rect 15252 46288 15258 46300
rect 251818 46288 251824 46300
rect 15252 46260 251824 46288
rect 15252 46248 15258 46260
rect 251818 46248 251824 46260
rect 251876 46248 251882 46300
rect 62022 46180 62028 46232
rect 62080 46220 62086 46232
rect 327718 46220 327724 46232
rect 62080 46192 327724 46220
rect 62080 46180 62086 46192
rect 327718 46180 327724 46192
rect 327776 46180 327782 46232
rect 338114 46180 338120 46232
rect 338172 46220 338178 46232
rect 367094 46220 367100 46232
rect 338172 46192 367100 46220
rect 338172 46180 338178 46192
rect 367094 46180 367100 46192
rect 367152 46220 367158 46232
rect 367830 46220 367836 46232
rect 367152 46192 367836 46220
rect 367152 46180 367158 46192
rect 367830 46180 367836 46192
rect 367888 46180 367894 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 14458 45540 14464 45552
rect 3476 45512 14464 45540
rect 3476 45500 3482 45512
rect 14458 45500 14464 45512
rect 14516 45500 14522 45552
rect 182818 45500 182824 45552
rect 182876 45540 182882 45552
rect 296714 45540 296720 45552
rect 182876 45512 296720 45540
rect 182876 45500 182882 45512
rect 296714 45500 296720 45512
rect 296772 45540 296778 45552
rect 297634 45540 297640 45552
rect 296772 45512 297640 45540
rect 296772 45500 296778 45512
rect 297634 45500 297640 45512
rect 297692 45500 297698 45552
rect 48314 44820 48320 44872
rect 48372 44860 48378 44872
rect 258718 44860 258724 44872
rect 48372 44832 258724 44860
rect 48372 44820 48378 44832
rect 258718 44820 258724 44832
rect 258776 44820 258782 44872
rect 298830 44820 298836 44872
rect 298888 44860 298894 44872
rect 360838 44860 360844 44872
rect 298888 44832 360844 44860
rect 298888 44820 298894 44832
rect 360838 44820 360844 44832
rect 360896 44820 360902 44872
rect 113174 43460 113180 43512
rect 113232 43500 113238 43512
rect 250530 43500 250536 43512
rect 113232 43472 250536 43500
rect 113232 43460 113238 43472
rect 250530 43460 250536 43472
rect 250588 43460 250594 43512
rect 89714 43392 89720 43444
rect 89772 43432 89778 43444
rect 305822 43432 305828 43444
rect 89772 43404 305828 43432
rect 89772 43392 89778 43404
rect 305822 43392 305828 43404
rect 305880 43392 305886 43444
rect 317322 43392 317328 43444
rect 317380 43432 317386 43444
rect 427814 43432 427820 43444
rect 317380 43404 427820 43432
rect 317380 43392 317386 43404
rect 427814 43392 427820 43404
rect 427872 43392 427878 43444
rect 313274 42712 313280 42764
rect 313332 42752 313338 42764
rect 313918 42752 313924 42764
rect 313332 42724 313924 42752
rect 313332 42712 313338 42724
rect 313918 42712 313924 42724
rect 313976 42752 313982 42764
rect 429194 42752 429200 42764
rect 313976 42724 429200 42752
rect 313976 42712 313982 42724
rect 429194 42712 429200 42724
rect 429252 42712 429258 42764
rect 35986 42032 35992 42084
rect 36044 42072 36050 42084
rect 285122 42072 285128 42084
rect 36044 42044 285128 42072
rect 36044 42032 36050 42044
rect 285122 42032 285128 42044
rect 285180 42032 285186 42084
rect 342346 41352 342352 41404
rect 342404 41392 342410 41404
rect 430574 41392 430580 41404
rect 342404 41364 430580 41392
rect 342404 41352 342410 41364
rect 430574 41352 430580 41364
rect 430632 41352 430638 41404
rect 38562 40808 38568 40860
rect 38620 40848 38626 40860
rect 132494 40848 132500 40860
rect 38620 40820 132500 40848
rect 38620 40808 38626 40820
rect 132494 40808 132500 40820
rect 132552 40808 132558 40860
rect 120074 40740 120080 40792
rect 120132 40780 120138 40792
rect 253198 40780 253204 40792
rect 120132 40752 253204 40780
rect 120132 40740 120138 40752
rect 253198 40740 253204 40752
rect 253256 40740 253262 40792
rect 93946 40672 93952 40724
rect 94004 40712 94010 40724
rect 302970 40712 302976 40724
rect 94004 40684 302976 40712
rect 94004 40672 94010 40684
rect 302970 40672 302976 40684
rect 303028 40672 303034 40724
rect 309134 40060 309140 40112
rect 309192 40100 309198 40112
rect 342346 40100 342352 40112
rect 309192 40072 342352 40100
rect 309192 40060 309198 40072
rect 342346 40060 342352 40072
rect 342404 40060 342410 40112
rect 288342 39584 288348 39636
rect 288400 39624 288406 39636
rect 335998 39624 336004 39636
rect 288400 39596 336004 39624
rect 288400 39584 288406 39596
rect 335998 39584 336004 39596
rect 336056 39584 336062 39636
rect 210418 39516 210424 39568
rect 210476 39556 210482 39568
rect 302234 39556 302240 39568
rect 210476 39528 302240 39556
rect 210476 39516 210482 39528
rect 302234 39516 302240 39528
rect 302292 39516 302298 39568
rect 185578 39448 185584 39500
rect 185636 39488 185642 39500
rect 300762 39488 300768 39500
rect 185636 39460 300768 39488
rect 185636 39448 185642 39460
rect 300762 39448 300768 39460
rect 300820 39448 300826 39500
rect 117314 39380 117320 39432
rect 117372 39420 117378 39432
rect 287790 39420 287796 39432
rect 117372 39392 287796 39420
rect 117372 39380 117378 39392
rect 287790 39380 287796 39392
rect 287848 39380 287854 39432
rect 11146 39312 11152 39364
rect 11204 39352 11210 39364
rect 272610 39352 272616 39364
rect 11204 39324 272616 39352
rect 11204 39312 11210 39324
rect 272610 39312 272616 39324
rect 272668 39312 272674 39364
rect 302234 39312 302240 39364
rect 302292 39352 302298 39364
rect 433334 39352 433340 39364
rect 302292 39324 433340 39352
rect 302292 39312 302298 39324
rect 433334 39312 433340 39324
rect 433392 39312 433398 39364
rect 300762 38632 300768 38684
rect 300820 38672 300826 38684
rect 307202 38672 307208 38684
rect 300820 38644 307208 38672
rect 300820 38632 300826 38644
rect 307202 38632 307208 38644
rect 307260 38632 307266 38684
rect 232498 38020 232504 38072
rect 232556 38060 232562 38072
rect 299474 38060 299480 38072
rect 232556 38032 299480 38060
rect 232556 38020 232562 38032
rect 299474 38020 299480 38032
rect 299532 38020 299538 38072
rect 92474 37952 92480 38004
rect 92532 37992 92538 38004
rect 300118 37992 300124 38004
rect 92532 37964 300124 37992
rect 92532 37952 92538 37964
rect 300118 37952 300124 37964
rect 300176 37952 300182 38004
rect 26234 37884 26240 37936
rect 26292 37924 26298 37936
rect 264422 37924 264428 37936
rect 26292 37896 264428 37924
rect 26292 37884 26298 37896
rect 264422 37884 264428 37896
rect 264480 37884 264486 37936
rect 299474 37884 299480 37936
rect 299532 37924 299538 37936
rect 434714 37924 434720 37936
rect 299532 37896 434720 37924
rect 299532 37884 299538 37896
rect 434714 37884 434720 37896
rect 434772 37884 434778 37936
rect 222838 37204 222844 37256
rect 222896 37244 222902 37256
rect 287054 37244 287060 37256
rect 222896 37216 287060 37244
rect 222896 37204 222902 37216
rect 287054 37204 287060 37216
rect 287112 37244 287118 37256
rect 288342 37244 288348 37256
rect 287112 37216 288348 37244
rect 287112 37204 287118 37216
rect 288342 37204 288348 37216
rect 288400 37204 288406 37256
rect 211798 36592 211804 36644
rect 211856 36632 211862 36644
rect 295334 36632 295340 36644
rect 211856 36604 295340 36632
rect 211856 36592 211862 36604
rect 295334 36592 295340 36604
rect 295392 36632 295398 36644
rect 295392 36604 296714 36632
rect 295392 36592 295398 36604
rect 2774 36524 2780 36576
rect 2832 36564 2838 36576
rect 269758 36564 269764 36576
rect 2832 36536 269764 36564
rect 2832 36524 2838 36536
rect 269758 36524 269764 36536
rect 269816 36524 269822 36576
rect 296686 36564 296714 36604
rect 436186 36564 436192 36576
rect 296686 36536 436192 36564
rect 436186 36524 436192 36536
rect 436244 36524 436250 36576
rect 206278 35300 206284 35352
rect 206336 35340 206342 35352
rect 293954 35340 293960 35352
rect 206336 35312 293960 35340
rect 206336 35300 206342 35312
rect 293954 35300 293960 35312
rect 294012 35300 294018 35352
rect 111794 35232 111800 35284
rect 111852 35272 111858 35284
rect 301682 35272 301688 35284
rect 111852 35244 301688 35272
rect 111852 35232 111858 35244
rect 301682 35232 301688 35244
rect 301740 35232 301746 35284
rect 44082 35164 44088 35216
rect 44140 35204 44146 35216
rect 264330 35204 264336 35216
rect 44140 35176 264336 35204
rect 44140 35164 44146 35176
rect 264330 35164 264336 35176
rect 264388 35164 264394 35216
rect 293954 35164 293960 35216
rect 294012 35204 294018 35216
rect 436278 35204 436284 35216
rect 294012 35176 436284 35204
rect 294012 35164 294018 35176
rect 436278 35164 436284 35176
rect 436336 35164 436342 35216
rect 289078 34416 289084 34468
rect 289136 34456 289142 34468
rect 437474 34456 437480 34468
rect 289136 34428 437480 34456
rect 289136 34416 289142 34428
rect 437474 34416 437480 34428
rect 437532 34416 437538 34468
rect 41414 33804 41420 33856
rect 41472 33844 41478 33856
rect 273898 33844 273904 33856
rect 41472 33816 273904 33844
rect 41472 33804 41478 33816
rect 273898 33804 273904 33816
rect 273956 33804 273962 33856
rect 30374 33736 30380 33788
rect 30432 33776 30438 33788
rect 290458 33776 290464 33788
rect 30432 33748 290464 33776
rect 30432 33736 30438 33748
rect 290458 33736 290464 33748
rect 290516 33736 290522 33788
rect 288434 33124 288440 33176
rect 288492 33164 288498 33176
rect 289078 33164 289084 33176
rect 288492 33136 289084 33164
rect 288492 33124 288498 33136
rect 289078 33124 289084 33136
rect 289136 33124 289142 33176
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 21358 33096 21364 33108
rect 3568 33068 21364 33096
rect 3568 33056 3574 33068
rect 21358 33056 21364 33068
rect 21416 33056 21422 33108
rect 327718 33056 327724 33108
rect 327776 33096 327782 33108
rect 425054 33096 425060 33108
rect 327776 33068 425060 33096
rect 327776 33056 327782 33068
rect 425054 33056 425060 33068
rect 425112 33056 425118 33108
rect 118786 32444 118792 32496
rect 118844 32484 118850 32496
rect 304350 32484 304356 32496
rect 118844 32456 304356 32484
rect 118844 32444 118850 32456
rect 304350 32444 304356 32456
rect 304408 32444 304414 32496
rect 95234 32376 95240 32428
rect 95292 32416 95298 32428
rect 280982 32416 280988 32428
rect 95292 32388 280988 32416
rect 95292 32376 95298 32388
rect 280982 32376 280988 32388
rect 281040 32376 281046 32428
rect 327074 31764 327080 31816
rect 327132 31804 327138 31816
rect 327718 31804 327724 31816
rect 327132 31776 327724 31804
rect 327132 31764 327138 31776
rect 327718 31764 327724 31776
rect 327776 31764 327782 31816
rect 246298 31220 246304 31272
rect 246356 31260 246362 31272
rect 284386 31260 284392 31272
rect 246356 31232 284392 31260
rect 246356 31220 246362 31232
rect 284386 31220 284392 31232
rect 284444 31260 284450 31272
rect 284444 31232 287054 31260
rect 284444 31220 284450 31232
rect 85574 31152 85580 31204
rect 85632 31192 85638 31204
rect 255958 31192 255964 31204
rect 85632 31164 255964 31192
rect 85632 31152 85638 31164
rect 255958 31152 255964 31164
rect 256016 31152 256022 31204
rect 287026 31192 287054 31232
rect 438854 31192 438860 31204
rect 287026 31164 438860 31192
rect 438854 31152 438860 31164
rect 438912 31152 438918 31204
rect 100754 31084 100760 31136
rect 100812 31124 100818 31136
rect 289262 31124 289268 31136
rect 100812 31096 289268 31124
rect 100812 31084 100818 31096
rect 289262 31084 289268 31096
rect 289320 31084 289326 31136
rect 19426 31016 19432 31068
rect 19484 31056 19490 31068
rect 293218 31056 293224 31068
rect 19484 31028 293224 31056
rect 19484 31016 19490 31028
rect 293218 31016 293224 31028
rect 293276 31016 293282 31068
rect 277394 30268 277400 30320
rect 277452 30308 277458 30320
rect 278222 30308 278228 30320
rect 277452 30280 278228 30308
rect 277452 30268 277458 30280
rect 278222 30268 278228 30280
rect 278280 30308 278286 30320
rect 441614 30308 441620 30320
rect 278280 30280 441620 30308
rect 278280 30268 278286 30280
rect 441614 30268 441620 30280
rect 441672 30268 441678 30320
rect 110506 29656 110512 29708
rect 110564 29696 110570 29708
rect 250438 29696 250444 29708
rect 110564 29668 250444 29696
rect 110564 29656 110570 29668
rect 250438 29656 250444 29668
rect 250496 29656 250502 29708
rect 82814 29588 82820 29640
rect 82872 29628 82878 29640
rect 279418 29628 279424 29640
rect 82872 29600 279424 29628
rect 82872 29588 82878 29600
rect 279418 29588 279424 29600
rect 279476 29588 279482 29640
rect 59262 28908 59268 28960
rect 59320 28948 59326 28960
rect 298094 28948 298100 28960
rect 59320 28920 298100 28948
rect 59320 28908 59326 28920
rect 298094 28908 298100 28920
rect 298152 28948 298158 28960
rect 298830 28948 298836 28960
rect 298152 28920 298836 28948
rect 298152 28908 298158 28920
rect 298830 28908 298836 28920
rect 298888 28908 298894 28960
rect 213270 28296 213276 28348
rect 213328 28336 213334 28348
rect 274634 28336 274640 28348
rect 213328 28308 274640 28336
rect 213328 28296 213334 28308
rect 274634 28296 274640 28308
rect 274692 28336 274698 28348
rect 442994 28336 443000 28348
rect 274692 28308 443000 28336
rect 274692 28296 274698 28308
rect 442994 28296 443000 28308
rect 443052 28296 443058 28348
rect 44174 28228 44180 28280
rect 44232 28268 44238 28280
rect 276842 28268 276848 28280
rect 44232 28240 276848 28268
rect 44232 28228 44238 28240
rect 276842 28228 276848 28240
rect 276900 28228 276906 28280
rect 64506 27548 64512 27600
rect 64564 27588 64570 27600
rect 307754 27588 307760 27600
rect 64564 27560 307760 27588
rect 64564 27548 64570 27560
rect 307754 27548 307760 27560
rect 307812 27588 307818 27600
rect 308398 27588 308404 27600
rect 307812 27560 308404 27588
rect 307812 27548 307818 27560
rect 308398 27548 308404 27560
rect 308456 27548 308462 27600
rect 197998 26936 198004 26988
rect 198056 26976 198062 26988
rect 198056 26948 267734 26976
rect 198056 26936 198062 26948
rect 17954 26868 17960 26920
rect 18012 26908 18018 26920
rect 265710 26908 265716 26920
rect 18012 26880 265716 26908
rect 18012 26868 18018 26880
rect 265710 26868 265716 26880
rect 265768 26868 265774 26920
rect 267706 26908 267734 26948
rect 270494 26908 270500 26920
rect 267706 26880 270500 26908
rect 270494 26868 270500 26880
rect 270552 26908 270558 26920
rect 444374 26908 444380 26920
rect 270552 26880 444380 26908
rect 270552 26868 270558 26880
rect 444374 26868 444380 26880
rect 444432 26868 444438 26920
rect 216030 25576 216036 25628
rect 216088 25616 216094 25628
rect 271966 25616 271972 25628
rect 216088 25588 271972 25616
rect 216088 25576 216094 25588
rect 271966 25576 271972 25588
rect 272024 25616 272030 25628
rect 445846 25616 445852 25628
rect 272024 25588 445852 25616
rect 272024 25576 272030 25588
rect 445846 25576 445852 25588
rect 445904 25576 445910 25628
rect 20714 25508 20720 25560
rect 20772 25548 20778 25560
rect 296070 25548 296076 25560
rect 20772 25520 296076 25548
rect 20772 25508 20778 25520
rect 296070 25508 296076 25520
rect 296128 25508 296134 25560
rect 264330 24760 264336 24812
rect 264388 24800 264394 24812
rect 445938 24800 445944 24812
rect 264388 24772 445944 24800
rect 264388 24760 264394 24772
rect 445938 24760 445944 24772
rect 445996 24760 446002 24812
rect 96614 24216 96620 24268
rect 96672 24256 96678 24268
rect 302878 24256 302884 24268
rect 96672 24228 302884 24256
rect 96672 24216 96678 24228
rect 302878 24216 302884 24228
rect 302936 24216 302942 24268
rect 63494 24148 63500 24200
rect 63552 24188 63558 24200
rect 294598 24188 294604 24200
rect 63552 24160 294604 24188
rect 63552 24148 63558 24160
rect 294598 24148 294604 24160
rect 294656 24148 294662 24200
rect 2866 24080 2872 24132
rect 2924 24120 2930 24132
rect 264238 24120 264244 24132
rect 2924 24092 264244 24120
rect 2924 24080 2930 24092
rect 264238 24080 264244 24092
rect 264296 24080 264302 24132
rect 263594 23468 263600 23520
rect 263652 23508 263658 23520
rect 264330 23508 264336 23520
rect 263652 23480 264336 23508
rect 263652 23468 263658 23480
rect 264330 23468 264336 23480
rect 264388 23468 264394 23520
rect 77294 22856 77300 22908
rect 77352 22896 77358 22908
rect 260098 22896 260104 22908
rect 77352 22868 260104 22896
rect 77352 22856 77358 22868
rect 260098 22856 260104 22868
rect 260156 22856 260162 22908
rect 209038 22788 209044 22840
rect 209096 22828 209102 22840
rect 259546 22828 259552 22840
rect 209096 22800 259552 22828
rect 209096 22788 209102 22800
rect 259546 22788 259552 22800
rect 259604 22828 259610 22840
rect 447134 22828 447140 22840
rect 259604 22800 447140 22828
rect 259604 22788 259610 22800
rect 447134 22788 447140 22800
rect 447192 22788 447198 22840
rect 9674 22720 9680 22772
rect 9732 22760 9738 22772
rect 275278 22760 275284 22772
rect 9732 22732 275284 22760
rect 9732 22720 9738 22732
rect 275278 22720 275284 22732
rect 275336 22720 275342 22772
rect 253290 22040 253296 22092
rect 253348 22080 253354 22092
rect 449894 22080 449900 22092
rect 253348 22052 449900 22080
rect 253348 22040 253354 22052
rect 449894 22040 449900 22052
rect 449952 22040 449958 22092
rect 252554 21564 252560 21616
rect 252612 21604 252618 21616
rect 253290 21604 253296 21616
rect 252612 21576 253296 21604
rect 252612 21564 252618 21576
rect 253290 21564 253296 21576
rect 253348 21564 253354 21616
rect 69014 21496 69020 21548
rect 69072 21536 69078 21548
rect 257338 21536 257344 21548
rect 69072 21508 257344 21536
rect 69072 21496 69078 21508
rect 257338 21496 257344 21508
rect 257396 21496 257402 21548
rect 91094 21428 91100 21480
rect 91152 21468 91158 21480
rect 298738 21468 298744 21480
rect 91152 21440 298744 21468
rect 91152 21428 91158 21440
rect 298738 21428 298744 21440
rect 298796 21428 298802 21480
rect 67542 21360 67548 21412
rect 67600 21400 67606 21412
rect 329098 21400 329104 21412
rect 67600 21372 329104 21400
rect 67600 21360 67606 21372
rect 329098 21360 329104 21372
rect 329156 21400 329162 21412
rect 331950 21400 331956 21412
rect 329156 21372 331956 21400
rect 329156 21360 329162 21372
rect 331950 21360 331956 21372
rect 332008 21360 332014 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 22738 20652 22744 20664
rect 3476 20624 22744 20652
rect 3476 20612 3482 20624
rect 22738 20612 22744 20624
rect 22796 20612 22802 20664
rect 507118 20612 507124 20664
rect 507176 20652 507182 20664
rect 579982 20652 579988 20664
rect 507176 20624 579988 20652
rect 507176 20612 507182 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 232590 20000 232596 20052
rect 232648 20040 232654 20052
rect 249794 20040 249800 20052
rect 232648 20012 249800 20040
rect 232648 20000 232654 20012
rect 249794 20000 249800 20012
rect 249852 20040 249858 20052
rect 451274 20040 451280 20052
rect 249852 20012 451280 20040
rect 249852 20000 249858 20012
rect 451274 20000 451280 20012
rect 451332 20000 451338 20052
rect 22094 19932 22100 19984
rect 22152 19972 22158 19984
rect 307110 19972 307116 19984
rect 22152 19944 307116 19972
rect 22152 19932 22158 19944
rect 307110 19932 307116 19944
rect 307168 19932 307174 19984
rect 14 19252 20 19304
rect 72 19292 78 19304
rect 1302 19292 1308 19304
rect 72 19264 1308 19292
rect 72 19252 78 19264
rect 1302 19252 1308 19264
rect 1360 19292 1366 19304
rect 249150 19292 249156 19304
rect 1360 19264 249156 19292
rect 1360 19252 1366 19264
rect 249150 19252 249156 19264
rect 249208 19252 249214 19304
rect 104158 18708 104164 18760
rect 104216 18748 104222 18760
rect 307018 18748 307024 18760
rect 104216 18720 307024 18748
rect 104216 18708 104222 18720
rect 307018 18708 307024 18720
rect 307076 18708 307082 18760
rect 60826 18640 60832 18692
rect 60884 18680 60890 18692
rect 265618 18680 265624 18692
rect 60884 18652 265624 18680
rect 60884 18640 60890 18652
rect 265618 18640 265624 18652
rect 265676 18640 265682 18692
rect 246298 18572 246304 18624
rect 246356 18612 246362 18624
rect 452654 18612 452660 18624
rect 246356 18584 452660 18612
rect 246356 18572 246362 18584
rect 452654 18572 452660 18584
rect 452712 18572 452718 18624
rect 75914 17416 75920 17468
rect 75972 17456 75978 17468
rect 254578 17456 254584 17468
rect 75972 17428 254584 17456
rect 75972 17416 75978 17428
rect 254578 17416 254584 17428
rect 254636 17416 254642 17468
rect 244918 17348 244924 17400
rect 244976 17388 244982 17400
rect 454126 17388 454132 17400
rect 244976 17360 454132 17388
rect 244976 17348 244982 17360
rect 454126 17348 454132 17360
rect 454184 17348 454190 17400
rect 69106 17280 69112 17332
rect 69164 17320 69170 17332
rect 305730 17320 305736 17332
rect 69164 17292 305736 17320
rect 69164 17280 69170 17292
rect 305730 17280 305736 17292
rect 305788 17280 305794 17332
rect 13814 17212 13820 17264
rect 13872 17252 13878 17264
rect 283558 17252 283564 17264
rect 13872 17224 283564 17252
rect 13872 17212 13878 17224
rect 283558 17212 283564 17224
rect 283616 17212 283622 17264
rect 282270 15988 282276 16040
rect 282328 16028 282334 16040
rect 454034 16028 454040 16040
rect 282328 16000 454040 16028
rect 282328 15988 282334 16000
rect 454034 15988 454040 16000
rect 454092 15988 454098 16040
rect 85666 15920 85672 15972
rect 85724 15960 85730 15972
rect 286410 15960 286416 15972
rect 85724 15932 286416 15960
rect 85724 15920 85730 15932
rect 286410 15920 286416 15932
rect 286468 15920 286474 15972
rect 79226 15852 79232 15904
rect 79284 15892 79290 15904
rect 304258 15892 304264 15904
rect 79284 15864 304264 15892
rect 79284 15852 79290 15864
rect 304258 15852 304264 15864
rect 304316 15852 304322 15904
rect 337010 15104 337016 15156
rect 337068 15144 337074 15156
rect 501046 15144 501052 15156
rect 337068 15116 501052 15144
rect 337068 15104 337074 15116
rect 501046 15104 501052 15116
rect 501104 15104 501110 15156
rect 39114 14560 39120 14612
rect 39172 14600 39178 14612
rect 284938 14600 284944 14612
rect 39172 14572 284944 14600
rect 39172 14560 39178 14572
rect 284938 14560 284944 14572
rect 284996 14560 285002 14612
rect 17034 14492 17040 14544
rect 17092 14532 17098 14544
rect 262858 14532 262864 14544
rect 17092 14504 262864 14532
rect 17092 14492 17098 14504
rect 262858 14492 262864 14504
rect 262916 14492 262922 14544
rect 164418 14424 164424 14476
rect 164476 14464 164482 14476
rect 417418 14464 417424 14476
rect 164476 14436 417424 14464
rect 164476 14424 164482 14436
rect 417418 14424 417424 14436
rect 417476 14424 417482 14476
rect 314654 13744 314660 13796
rect 314712 13784 314718 13796
rect 315298 13784 315304 13796
rect 314712 13756 315304 13784
rect 314712 13744 314718 13756
rect 315298 13744 315304 13756
rect 315356 13784 315362 13796
rect 467834 13784 467840 13796
rect 315356 13756 467840 13784
rect 315356 13744 315362 13756
rect 467834 13744 467840 13756
rect 467892 13744 467898 13796
rect 249242 13676 249248 13728
rect 249300 13716 249306 13728
rect 358078 13716 358084 13728
rect 249300 13688 358084 13716
rect 249300 13676 249306 13688
rect 358078 13676 358084 13688
rect 358136 13676 358142 13728
rect 58434 13064 58440 13116
rect 58492 13104 58498 13116
rect 276750 13104 276756 13116
rect 58492 13076 276756 13104
rect 58492 13064 58498 13076
rect 276750 13064 276756 13076
rect 276808 13064 276814 13116
rect 248414 12452 248420 12504
rect 248472 12492 248478 12504
rect 249242 12492 249248 12504
rect 248472 12464 249248 12492
rect 248472 12452 248478 12464
rect 249242 12452 249248 12464
rect 249300 12452 249306 12504
rect 202138 11772 202144 11824
rect 202196 11812 202202 11824
rect 255866 11812 255872 11824
rect 202196 11784 255872 11812
rect 202196 11772 202202 11784
rect 255866 11772 255872 11784
rect 255924 11812 255930 11824
rect 353938 11812 353944 11824
rect 255924 11784 353944 11812
rect 255924 11772 255930 11784
rect 353938 11772 353944 11784
rect 353996 11772 354002 11824
rect 34514 11704 34520 11756
rect 34572 11744 34578 11756
rect 280890 11744 280896 11756
rect 34572 11716 280896 11744
rect 34572 11704 34578 11716
rect 280890 11704 280896 11716
rect 280948 11704 280954 11756
rect 283558 11704 283564 11756
rect 283616 11744 283622 11756
rect 478874 11744 478880 11756
rect 283616 11716 478880 11744
rect 283616 11704 283622 11716
rect 478874 11704 478880 11716
rect 478932 11704 478938 11756
rect 63034 10344 63040 10396
rect 63092 10384 63098 10396
rect 282362 10384 282368 10396
rect 63092 10356 282368 10384
rect 63092 10344 63098 10356
rect 282362 10344 282368 10356
rect 282420 10344 282426 10396
rect 305546 10344 305552 10396
rect 305604 10384 305610 10396
rect 331858 10384 331864 10396
rect 305604 10356 331864 10384
rect 305604 10344 305610 10356
rect 331858 10344 331864 10356
rect 331916 10344 331922 10396
rect 226978 10276 226984 10328
rect 227036 10316 227042 10328
rect 258258 10316 258264 10328
rect 227036 10288 258264 10316
rect 227036 10276 227042 10288
rect 258258 10276 258264 10288
rect 258316 10316 258322 10328
rect 486418 10316 486424 10328
rect 258316 10288 486424 10316
rect 258316 10276 258322 10288
rect 486418 10276 486424 10288
rect 486476 10276 486482 10328
rect 186958 9596 186964 9648
rect 187016 9636 187022 9648
rect 324958 9636 324964 9648
rect 187016 9608 324964 9636
rect 187016 9596 187022 9608
rect 324958 9596 324964 9608
rect 325016 9636 325022 9648
rect 325602 9636 325608 9648
rect 325016 9608 325608 9636
rect 325016 9596 325022 9608
rect 325602 9596 325608 9608
rect 325660 9596 325666 9648
rect 369854 9596 369860 9648
rect 369912 9636 369918 9648
rect 499758 9636 499764 9648
rect 369912 9608 499764 9636
rect 369912 9596 369918 9608
rect 499758 9596 499764 9608
rect 499816 9596 499822 9648
rect 332042 9528 332048 9580
rect 332100 9568 332106 9580
rect 423674 9568 423680 9580
rect 332100 9540 423680 9568
rect 332100 9528 332106 9540
rect 423674 9528 423680 9540
rect 423732 9528 423738 9580
rect 331582 9256 331588 9308
rect 331640 9296 331646 9308
rect 332042 9296 332048 9308
rect 331640 9268 332048 9296
rect 331640 9256 331646 9268
rect 332042 9256 332048 9268
rect 332100 9256 332106 9308
rect 3418 8984 3424 9036
rect 3476 9024 3482 9036
rect 29638 9024 29644 9036
rect 3476 8996 29644 9024
rect 3476 8984 3482 8996
rect 29638 8984 29644 8996
rect 29696 8984 29702 9036
rect 65518 8984 65524 9036
rect 65576 9024 65582 9036
rect 283650 9024 283656 9036
rect 65576 8996 283656 9024
rect 65576 8984 65582 8996
rect 283650 8984 283656 8996
rect 283708 8984 283714 9036
rect 13538 8916 13544 8968
rect 13596 8956 13602 8968
rect 249058 8956 249064 8968
rect 13596 8928 249064 8956
rect 13596 8916 13602 8928
rect 249058 8916 249064 8928
rect 249116 8916 249122 8968
rect 319714 8916 319720 8968
rect 319772 8956 319778 8968
rect 334618 8956 334624 8968
rect 319772 8928 334624 8956
rect 319772 8916 319778 8928
rect 334618 8916 334624 8928
rect 334676 8916 334682 8968
rect 340966 8916 340972 8968
rect 341024 8956 341030 8968
rect 369854 8956 369860 8968
rect 341024 8928 369860 8956
rect 341024 8916 341030 8928
rect 369854 8916 369860 8928
rect 369912 8916 369918 8968
rect 181438 8236 181444 8288
rect 181496 8276 181502 8288
rect 283558 8276 283564 8288
rect 181496 8248 283564 8276
rect 181496 8236 181502 8248
rect 283558 8236 283564 8248
rect 283616 8236 283622 8288
rect 339954 8236 339960 8288
rect 340012 8276 340018 8288
rect 431954 8276 431960 8288
rect 340012 8248 431960 8276
rect 340012 8236 340018 8248
rect 431954 8236 431960 8248
rect 432012 8236 432018 8288
rect 280798 8168 280804 8220
rect 280856 8208 280862 8220
rect 344278 8208 344284 8220
rect 280856 8180 344284 8208
rect 280856 8168 280862 8180
rect 344278 8168 344284 8180
rect 344336 8168 344342 8220
rect 215938 7624 215944 7676
rect 215996 7664 216002 7676
rect 301774 7664 301780 7676
rect 215996 7636 301780 7664
rect 215996 7624 216002 7636
rect 301774 7624 301780 7636
rect 301832 7624 301838 7676
rect 8754 7556 8760 7608
rect 8812 7596 8818 7608
rect 266998 7596 267004 7608
rect 8812 7568 267004 7596
rect 8812 7556 8818 7568
rect 266998 7556 267004 7568
rect 267056 7556 267062 7608
rect 306742 6876 306748 6928
rect 306800 6916 306806 6928
rect 339954 6916 339960 6928
rect 306800 6888 339960 6916
rect 306800 6876 306806 6888
rect 339954 6876 339960 6888
rect 340012 6876 340018 6928
rect 174538 6808 174544 6860
rect 174596 6848 174602 6860
rect 242158 6848 242164 6860
rect 174596 6820 242164 6848
rect 174596 6808 174602 6820
rect 242158 6808 242164 6820
rect 242216 6808 242222 6860
rect 281902 6808 281908 6860
rect 281960 6848 281966 6860
rect 439498 6848 439504 6860
rect 281960 6820 439504 6848
rect 281960 6808 281966 6820
rect 439498 6808 439504 6820
rect 439556 6808 439562 6860
rect 542998 6808 543004 6860
rect 543056 6848 543062 6860
rect 580166 6848 580172 6860
rect 543056 6820 580172 6848
rect 543056 6808 543062 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 301774 6740 301780 6792
rect 301832 6780 301838 6792
rect 363598 6780 363604 6792
rect 301832 6752 363604 6780
rect 301832 6740 301838 6752
rect 363598 6740 363604 6752
rect 363656 6740 363662 6792
rect 308490 6672 308496 6724
rect 308548 6712 308554 6724
rect 309870 6712 309876 6724
rect 308548 6684 309876 6712
rect 308548 6672 308554 6684
rect 309870 6672 309876 6684
rect 309928 6672 309934 6724
rect 35802 6264 35808 6316
rect 35860 6304 35866 6316
rect 136450 6304 136456 6316
rect 35860 6276 136456 6304
rect 35860 6264 35866 6276
rect 136450 6264 136456 6276
rect 136508 6264 136514 6316
rect 104526 6196 104532 6248
rect 104584 6236 104590 6248
rect 305638 6236 305644 6248
rect 104584 6208 305644 6236
rect 104584 6196 104590 6208
rect 305638 6196 305644 6208
rect 305696 6196 305702 6248
rect 28902 6128 28908 6180
rect 28960 6168 28966 6180
rect 295978 6168 295984 6180
rect 28960 6140 295984 6168
rect 28960 6128 28966 6140
rect 295978 6128 295984 6140
rect 296036 6128 296042 6180
rect 63126 5448 63132 5500
rect 63184 5488 63190 5500
rect 251174 5488 251180 5500
rect 63184 5460 251180 5488
rect 63184 5448 63190 5460
rect 251174 5448 251180 5460
rect 251232 5448 251238 5500
rect 257062 5448 257068 5500
rect 257120 5488 257126 5500
rect 257430 5488 257436 5500
rect 257120 5460 257436 5488
rect 257120 5448 257126 5460
rect 257430 5448 257436 5460
rect 257488 5488 257494 5500
rect 448514 5488 448520 5500
rect 257488 5460 448520 5488
rect 257488 5448 257494 5460
rect 448514 5448 448520 5460
rect 448572 5448 448578 5500
rect 251174 4972 251180 5024
rect 251232 5012 251238 5024
rect 251910 5012 251916 5024
rect 251232 4984 251916 5012
rect 251232 4972 251238 4984
rect 251910 4972 251916 4984
rect 251968 4972 251974 5024
rect 180058 4904 180064 4956
rect 180116 4944 180122 4956
rect 239214 4944 239220 4956
rect 180116 4916 239220 4944
rect 180116 4904 180122 4916
rect 239214 4904 239220 4916
rect 239272 4904 239278 4956
rect 213178 4836 213184 4888
rect 213236 4876 213242 4888
rect 294874 4876 294880 4888
rect 213236 4848 294880 4876
rect 213236 4836 213242 4848
rect 294874 4836 294880 4848
rect 294932 4876 294938 4888
rect 294932 4848 296714 4876
rect 294932 4836 294938 4848
rect 27706 4768 27712 4820
rect 27764 4808 27770 4820
rect 291930 4808 291936 4820
rect 27764 4780 291936 4808
rect 27764 4768 27770 4780
rect 291930 4768 291936 4780
rect 291988 4768 291994 4820
rect 296686 4808 296714 4848
rect 356790 4808 356796 4820
rect 296686 4780 356796 4808
rect 356790 4768 356796 4780
rect 356848 4768 356854 4820
rect 191098 4088 191104 4140
rect 191156 4128 191162 4140
rect 246390 4128 246396 4140
rect 191156 4100 246396 4128
rect 191156 4088 191162 4100
rect 246390 4088 246396 4100
rect 246448 4088 246454 4140
rect 300762 4088 300768 4140
rect 300820 4128 300826 4140
rect 307202 4128 307208 4140
rect 300820 4100 307208 4128
rect 300820 4088 300826 4100
rect 307202 4088 307208 4100
rect 307260 4088 307266 4140
rect 332686 4088 332692 4140
rect 332744 4128 332750 4140
rect 333238 4128 333244 4140
rect 332744 4100 333244 4128
rect 332744 4088 332750 4100
rect 333238 4088 333244 4100
rect 333296 4128 333302 4140
rect 352558 4128 352564 4140
rect 333296 4100 352564 4128
rect 333296 4088 333302 4100
rect 352558 4088 352564 4100
rect 352616 4088 352622 4140
rect 239214 4020 239220 4072
rect 239272 4060 239278 4072
rect 282270 4060 282276 4072
rect 239272 4032 282276 4060
rect 239272 4020 239278 4032
rect 282270 4020 282276 4032
rect 282328 4020 282334 4072
rect 349798 4020 349804 4072
rect 349856 4060 349862 4072
rect 350442 4060 350448 4072
rect 349856 4032 350448 4060
rect 349856 4020 349862 4032
rect 350442 4020 350448 4032
rect 350500 4060 350506 4072
rect 377398 4060 377404 4072
rect 350500 4032 377404 4060
rect 350500 4020 350506 4032
rect 377398 4020 377404 4032
rect 377456 4020 377462 4072
rect 347038 3952 347044 4004
rect 347096 3992 347102 4004
rect 354030 3992 354036 4004
rect 347096 3964 354036 3992
rect 347096 3952 347102 3964
rect 354030 3952 354036 3964
rect 354088 3952 354094 4004
rect 351178 3884 351184 3936
rect 351236 3924 351242 3936
rect 351638 3924 351644 3936
rect 351236 3896 351644 3924
rect 351236 3884 351242 3896
rect 351638 3884 351644 3896
rect 351696 3924 351702 3936
rect 495526 3924 495532 3936
rect 351696 3896 495532 3924
rect 351696 3884 351702 3896
rect 495526 3884 495532 3896
rect 495584 3884 495590 3936
rect 125870 3680 125876 3732
rect 125928 3720 125934 3732
rect 164878 3720 164884 3732
rect 125928 3692 164884 3720
rect 125928 3680 125934 3692
rect 164878 3680 164884 3692
rect 164936 3680 164942 3732
rect 78582 3612 78588 3664
rect 78640 3652 78646 3664
rect 104158 3652 104164 3664
rect 78640 3624 104164 3652
rect 78640 3612 78646 3624
rect 104158 3612 104164 3624
rect 104216 3612 104222 3664
rect 109310 3612 109316 3664
rect 109368 3652 109374 3664
rect 171778 3652 171784 3664
rect 109368 3624 171784 3652
rect 109368 3612 109374 3624
rect 171778 3612 171784 3624
rect 171836 3612 171842 3664
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 79318 3584 79324 3596
rect 6512 3556 79324 3584
rect 6512 3544 6518 3556
rect 79318 3544 79324 3556
rect 79376 3544 79382 3596
rect 85574 3544 85580 3596
rect 85632 3584 85638 3596
rect 86494 3584 86500 3596
rect 85632 3556 86500 3584
rect 85632 3544 85638 3556
rect 86494 3544 86500 3556
rect 86552 3544 86558 3596
rect 93854 3544 93860 3596
rect 93912 3584 93918 3596
rect 94774 3584 94780 3596
rect 93912 3556 94780 3584
rect 93912 3544 93918 3556
rect 94774 3544 94780 3556
rect 94832 3544 94838 3596
rect 103330 3544 103336 3596
rect 103388 3584 103394 3596
rect 195422 3584 195428 3596
rect 103388 3556 195428 3584
rect 103388 3544 103394 3556
rect 195422 3544 195428 3556
rect 195480 3544 195486 3596
rect 242986 3544 242992 3596
rect 243044 3584 243050 3596
rect 244918 3584 244924 3596
rect 243044 3556 244924 3584
rect 243044 3544 243050 3556
rect 244918 3544 244924 3556
rect 244976 3544 244982 3596
rect 267734 3544 267740 3596
rect 267792 3584 267798 3596
rect 271966 3584 271972 3596
rect 267792 3556 271972 3584
rect 267792 3544 267798 3556
rect 271966 3544 271972 3556
rect 272024 3544 272030 3596
rect 316126 3544 316132 3596
rect 316184 3584 316190 3596
rect 317322 3584 317328 3596
rect 316184 3556 317328 3584
rect 316184 3544 316190 3556
rect 317322 3544 317328 3556
rect 317380 3544 317386 3596
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3694 3516 3700 3528
rect 2832 3488 3700 3516
rect 2832 3476 2838 3488
rect 3694 3476 3700 3488
rect 3752 3476 3758 3528
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 20254 3516 20260 3528
rect 19392 3488 20260 3516
rect 19392 3476 19398 3488
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 33042 3476 33048 3528
rect 33100 3516 33106 3528
rect 150618 3516 150624 3528
rect 33100 3488 150624 3516
rect 33100 3476 33106 3488
rect 150618 3476 150624 3488
rect 150676 3476 150682 3528
rect 242894 3476 242900 3528
rect 242952 3516 242958 3528
rect 244090 3516 244096 3528
rect 242952 3488 244096 3516
rect 242952 3476 242958 3488
rect 244090 3476 244096 3488
rect 244148 3476 244154 3528
rect 307754 3476 307760 3528
rect 307812 3516 307818 3528
rect 309042 3516 309048 3528
rect 307812 3488 309048 3516
rect 307812 3476 307818 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 332594 3476 332600 3528
rect 332652 3516 332658 3528
rect 333882 3516 333888 3528
rect 332652 3488 333888 3516
rect 332652 3476 332658 3488
rect 333882 3476 333888 3488
rect 333940 3476 333946 3528
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 188522 3448 188528 3460
rect 24268 3420 188528 3448
rect 24268 3408 24274 3420
rect 188522 3408 188528 3420
rect 188580 3408 188586 3460
rect 276014 3408 276020 3460
rect 276072 3448 276078 3460
rect 276750 3448 276756 3460
rect 276072 3420 276756 3448
rect 276072 3408 276078 3420
rect 276750 3408 276756 3420
rect 276808 3408 276814 3460
rect 44174 3340 44180 3392
rect 44232 3380 44238 3392
rect 45094 3380 45100 3392
rect 44232 3352 45100 3380
rect 44232 3340 44238 3352
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 52454 3340 52460 3392
rect 52512 3380 52518 3392
rect 53374 3380 53380 3392
rect 52512 3352 53380 3380
rect 52512 3340 52518 3352
rect 53374 3340 53380 3352
rect 53432 3340 53438 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 118694 3340 118700 3392
rect 118752 3380 118758 3392
rect 119890 3380 119896 3392
rect 118752 3352 119896 3380
rect 118752 3340 118758 3352
rect 119890 3340 119896 3352
rect 119948 3340 119954 3392
rect 1670 3272 1676 3324
rect 1728 3312 1734 3324
rect 7742 3312 7748 3324
rect 1728 3284 7748 3312
rect 1728 3272 1734 3284
rect 7742 3272 7748 3284
rect 7800 3272 7806 3324
rect 235810 3068 235816 3120
rect 235868 3108 235874 3120
rect 238018 3108 238024 3120
rect 235868 3080 238024 3108
rect 235868 3068 235874 3080
rect 238018 3068 238024 3080
rect 238076 3068 238082 3120
rect 292574 3000 292580 3052
rect 292632 3040 292638 3052
rect 293954 3040 293960 3052
rect 292632 3012 293960 3040
rect 292632 3000 292638 3012
rect 293954 3000 293960 3012
rect 294012 3000 294018 3052
rect 43070 2116 43076 2168
rect 43128 2156 43134 2168
rect 301498 2156 301504 2168
rect 43128 2128 301504 2156
rect 43128 2116 43134 2128
rect 301498 2116 301504 2128
rect 301556 2116 301562 2168
rect 30098 2048 30104 2100
rect 30156 2088 30162 2100
rect 301590 2088 301596 2100
rect 30156 2060 301596 2088
rect 30156 2048 30162 2060
rect 301590 2048 301596 2060
rect 301648 2048 301654 2100
<< via1 >>
rect 201500 703264 201552 703316
rect 202788 703264 202840 703316
rect 82084 703196 82136 703248
rect 267648 703196 267700 703248
rect 99288 703128 99340 703180
rect 332508 703128 332560 703180
rect 115204 703060 115256 703112
rect 348792 703060 348844 703112
rect 79324 702992 79376 703044
rect 364340 702992 364392 703044
rect 364984 702992 365036 703044
rect 107568 702924 107620 702976
rect 413652 702924 413704 702976
rect 116584 702856 116636 702908
rect 462320 702856 462372 702908
rect 78588 702788 78640 702840
rect 429200 702788 429252 702840
rect 429844 702788 429896 702840
rect 71780 702720 71832 702772
rect 72976 702720 73028 702772
rect 113824 702720 113876 702772
rect 478512 702720 478564 702772
rect 115296 702652 115348 702704
rect 453948 702652 454000 702704
rect 492588 702652 492640 702704
rect 494796 702652 494848 702704
rect 69204 702584 69256 702636
rect 580908 702584 580960 702636
rect 113088 702516 113140 702568
rect 521568 702516 521620 702568
rect 550548 702516 550600 702568
rect 559656 702516 559708 702568
rect 80704 702448 80756 702500
rect 527180 702448 527232 702500
rect 519544 700952 519596 701004
rect 521568 700952 521620 701004
rect 40500 700340 40552 700392
rect 75184 700340 75236 700392
rect 129004 700340 129056 700392
rect 154120 700340 154172 700392
rect 188344 700340 188396 700392
rect 218980 700340 219032 700392
rect 62028 700272 62080 700324
rect 235172 700272 235224 700324
rect 238024 700272 238076 700324
rect 283840 700272 283892 700324
rect 450544 700272 450596 700324
rect 453948 700272 454000 700324
rect 492588 700272 492640 700324
rect 521568 700272 521620 700324
rect 550548 700272 550600 700324
rect 24308 697552 24360 697604
rect 110604 697552 110656 697604
rect 71044 692044 71096 692096
rect 136640 692044 136692 692096
rect 68928 690616 68980 690668
rect 169760 690616 169812 690668
rect 68652 687896 68704 687948
rect 129004 687896 129056 687948
rect 6920 686468 6972 686520
rect 89720 686468 89772 686520
rect 75184 685788 75236 685840
rect 77116 685788 77168 685840
rect 68836 685108 68888 685160
rect 238024 685108 238076 685160
rect 102232 683748 102284 683800
rect 188344 683748 188396 683800
rect 3424 683136 3476 683188
rect 75184 683136 75236 683188
rect 196624 683136 196676 683188
rect 580172 683136 580224 683188
rect 90640 681912 90692 681964
rect 59268 681844 59320 681896
rect 70032 681844 70084 681896
rect 57796 681776 57848 681828
rect 80704 681776 80756 681828
rect 4804 681708 4856 681760
rect 55128 681708 55180 681760
rect 109316 681708 109368 681760
rect 125692 681708 125744 681760
rect 53748 680960 53800 681012
rect 71780 680960 71832 681012
rect 104900 680960 104952 681012
rect 113180 680960 113232 681012
rect 69112 680348 69164 680400
rect 72608 680348 72660 680400
rect 84844 680348 84896 680400
rect 580264 680348 580316 680400
rect 69296 679328 69348 679380
rect 71044 679328 71096 679380
rect 111800 677628 111852 677680
rect 118700 677628 118752 677680
rect 64696 677560 64748 677612
rect 67640 677560 67692 677612
rect 112352 677560 112404 677612
rect 122932 677560 122984 677612
rect 111800 676268 111852 676320
rect 120356 676268 120408 676320
rect 33048 676200 33100 676252
rect 67640 676200 67692 676252
rect 112720 676200 112772 676252
rect 121552 676200 121604 676252
rect 55036 674908 55088 674960
rect 67640 674908 67692 674960
rect 111984 674840 112036 674892
rect 125784 674840 125836 674892
rect 66076 673684 66128 673736
rect 67732 673684 67784 673736
rect 48136 673480 48188 673532
rect 67640 673480 67692 673532
rect 111800 671984 111852 672036
rect 196624 671984 196676 672036
rect 65892 670760 65944 670812
rect 68652 670760 68704 670812
rect 63224 670692 63276 670744
rect 67640 670692 67692 670744
rect 111800 670692 111852 670744
rect 114560 670692 114612 670744
rect 111800 669468 111852 669520
rect 123024 669468 123076 669520
rect 66168 669400 66220 669452
rect 67824 669400 67876 669452
rect 112720 669400 112772 669452
rect 128452 669400 128504 669452
rect 64512 669332 64564 669384
rect 67640 669332 67692 669384
rect 111800 669332 111852 669384
rect 133972 669332 134024 669384
rect 67364 667904 67416 667956
rect 67732 667904 67784 667956
rect 65984 666612 66036 666664
rect 67824 666612 67876 666664
rect 61936 666544 61988 666596
rect 67640 666544 67692 666596
rect 68560 666544 68612 666596
rect 68836 666544 68888 666596
rect 111800 666544 111852 666596
rect 118792 666544 118844 666596
rect 44088 665252 44140 665304
rect 67732 665252 67784 665304
rect 42708 665184 42760 665236
rect 67640 665184 67692 665236
rect 111800 665184 111852 665236
rect 124404 665184 124456 665236
rect 61844 663824 61896 663876
rect 67640 663824 67692 663876
rect 112352 663824 112404 663876
rect 128544 663824 128596 663876
rect 52368 663756 52420 663808
rect 67732 663756 67784 663808
rect 111800 663756 111852 663808
rect 142160 663756 142212 663808
rect 62028 663008 62080 663060
rect 67640 663008 67692 663060
rect 111800 662396 111852 662448
rect 117412 662396 117464 662448
rect 53656 661648 53708 661700
rect 62028 661648 62080 661700
rect 111156 661512 111208 661564
rect 113824 661512 113876 661564
rect 60648 661036 60700 661088
rect 67640 661036 67692 661088
rect 59084 659744 59136 659796
rect 67640 659744 67692 659796
rect 112536 659744 112588 659796
rect 136732 659744 136784 659796
rect 50804 659676 50856 659728
rect 67732 659676 67784 659728
rect 112352 659676 112404 659728
rect 146300 659676 146352 659728
rect 39948 658928 40000 658980
rect 68560 658928 68612 658980
rect 109040 658384 109092 658436
rect 110604 658384 110656 658436
rect 63408 658248 63460 658300
rect 67640 658248 67692 658300
rect 2780 658180 2832 658232
rect 4804 658180 4856 658232
rect 133788 657500 133840 657552
rect 201500 657500 201552 657552
rect 56508 656956 56560 657008
rect 68192 656956 68244 657008
rect 49608 656888 49660 656940
rect 67732 656888 67784 656940
rect 112536 656888 112588 656940
rect 132500 656888 132552 656940
rect 133788 656888 133840 656940
rect 112536 655596 112588 655648
rect 121644 655596 121696 655648
rect 41236 655528 41288 655580
rect 67640 655528 67692 655580
rect 112352 655528 112404 655580
rect 139400 655528 139452 655580
rect 58624 654780 58676 654832
rect 67640 654780 67692 654832
rect 57888 652808 57940 652860
rect 67916 652808 67968 652860
rect 48044 652740 48096 652792
rect 67732 652740 67784 652792
rect 64788 651380 64840 651432
rect 67640 651380 67692 651432
rect 112536 651380 112588 651432
rect 129832 651380 129884 651432
rect 112076 650088 112128 650140
rect 119344 650088 119396 650140
rect 34428 650020 34480 650072
rect 67640 650020 67692 650072
rect 111984 650020 112036 650072
rect 143632 650020 143684 650072
rect 112996 648660 113048 648712
rect 115940 648660 115992 648712
rect 64604 648592 64656 648644
rect 67640 648592 67692 648644
rect 113088 648592 113140 648644
rect 138020 648592 138072 648644
rect 63132 647300 63184 647352
rect 67732 647300 67784 647352
rect 62028 647232 62080 647284
rect 67640 647232 67692 647284
rect 109408 647232 109460 647284
rect 112168 647232 112220 647284
rect 113088 647232 113140 647284
rect 143540 647232 143592 647284
rect 37096 645872 37148 645924
rect 67640 645872 67692 645924
rect 112996 644512 113048 644564
rect 132868 644512 132920 644564
rect 113088 644444 113140 644496
rect 135260 644444 135312 644496
rect 112812 644308 112864 644360
rect 115296 644308 115348 644360
rect 57796 643696 57848 643748
rect 69664 643696 69716 643748
rect 119344 643696 119396 643748
rect 134064 643696 134116 643748
rect 135168 643696 135220 643748
rect 135168 643084 135220 643136
rect 580172 643084 580224 643136
rect 116032 643016 116084 643068
rect 116584 643016 116636 643068
rect 112628 642064 112680 642116
rect 116032 642064 116084 642116
rect 61752 641792 61804 641844
rect 67732 641792 67784 641844
rect 37188 641724 37240 641776
rect 67640 641724 67692 641776
rect 113088 641724 113140 641776
rect 140780 641724 140832 641776
rect 63316 640364 63368 640416
rect 67640 640364 67692 640416
rect 34152 640296 34204 640348
rect 67732 640296 67784 640348
rect 108856 639616 108908 639668
rect 112260 639616 112312 639668
rect 124128 639548 124180 639600
rect 299480 639548 299532 639600
rect 38568 638936 38620 638988
rect 71320 638936 71372 638988
rect 112904 638936 112956 638988
rect 129924 638936 129976 638988
rect 46848 638868 46900 638920
rect 53748 638868 53800 638920
rect 73896 638868 73948 638920
rect 104164 638868 104216 638920
rect 122840 638868 122892 638920
rect 124128 638868 124180 638920
rect 72700 638460 72752 638512
rect 84200 638460 84252 638512
rect 95148 638460 95200 638512
rect 105544 638460 105596 638512
rect 108948 638460 109000 638512
rect 124312 638460 124364 638512
rect 57796 638392 57848 638444
rect 82268 638392 82320 638444
rect 99012 638392 99064 638444
rect 117320 638392 117372 638444
rect 54760 638324 54812 638376
rect 82912 638324 82964 638376
rect 99656 638324 99708 638376
rect 121460 638324 121512 638376
rect 48228 638256 48280 638308
rect 79048 638256 79100 638308
rect 102876 638256 102928 638308
rect 131120 638256 131172 638308
rect 3424 638188 3476 638240
rect 59176 638188 59228 638240
rect 91928 638188 91980 638240
rect 96436 638188 96488 638240
rect 124220 638188 124272 638240
rect 96528 637984 96580 638036
rect 99656 637984 99708 638036
rect 74448 637576 74500 637628
rect 93860 637576 93912 637628
rect 101404 637576 101456 637628
rect 75828 637508 75880 637560
rect 75920 637440 75972 637492
rect 77116 637440 77168 637492
rect 85580 637440 85632 637492
rect 86776 637440 86828 637492
rect 86960 637440 87012 637492
rect 88064 637440 88116 637492
rect 96620 637440 96672 637492
rect 97724 637440 97776 637492
rect 103612 637440 103664 637492
rect 104808 637440 104860 637492
rect 69204 637168 69256 637220
rect 69756 637168 69808 637220
rect 52276 636964 52328 637016
rect 78404 636964 78456 637016
rect 101588 636964 101640 637016
rect 128360 636964 128412 637016
rect 45376 636896 45428 636948
rect 74540 636896 74592 636948
rect 88708 636896 88760 636948
rect 118884 636896 118936 636948
rect 50988 636828 51040 636880
rect 84844 636828 84896 636880
rect 103520 636828 103572 636880
rect 136640 636828 136692 636880
rect 60372 635740 60424 635792
rect 71964 635740 72016 635792
rect 56324 635672 56376 635724
rect 73252 635672 73304 635724
rect 73804 635672 73856 635724
rect 92572 635672 92624 635724
rect 94504 635672 94556 635724
rect 120080 635672 120132 635724
rect 55128 635604 55180 635656
rect 80704 635604 80756 635656
rect 93216 635604 93268 635656
rect 126980 635604 127032 635656
rect 50712 635536 50764 635588
rect 80980 635536 81032 635588
rect 91284 635536 91336 635588
rect 125600 635536 125652 635588
rect 4068 635468 4120 635520
rect 96528 635468 96580 635520
rect 102232 635468 102284 635520
rect 133880 635468 133932 635520
rect 133880 634788 133932 634840
rect 579804 634788 579856 634840
rect 53748 634108 53800 634160
rect 87420 634108 87472 634160
rect 99932 634108 99984 634160
rect 132684 634108 132736 634160
rect 3424 634040 3476 634092
rect 108028 634040 108080 634092
rect 127164 634040 127216 634092
rect 107568 632952 107620 633004
rect 121552 632952 121604 633004
rect 54944 632884 54996 632936
rect 83556 632884 83608 632936
rect 57704 632816 57756 632868
rect 86132 632816 86184 632868
rect 89996 632816 90048 632868
rect 121552 632816 121604 632868
rect 52092 632748 52144 632800
rect 81624 632748 81676 632800
rect 97080 632748 97132 632800
rect 129740 632748 129792 632800
rect 39764 632680 39816 632732
rect 71780 632680 71832 632732
rect 96620 632680 96672 632732
rect 131304 632680 131356 632732
rect 45284 629960 45336 630012
rect 70676 629960 70728 630012
rect 42524 629892 42576 629944
rect 76472 629892 76524 629944
rect 98368 629892 98420 629944
rect 131764 629892 131816 629944
rect 46756 627308 46808 627360
rect 75920 627308 75972 627360
rect 49332 627240 49384 627292
rect 79692 627240 79744 627292
rect 43996 627172 44048 627224
rect 74632 627172 74684 627224
rect 3516 618604 3568 618656
rect 7564 618604 7616 618656
rect 115848 618196 115900 618248
rect 118884 618196 118936 618248
rect 580172 618196 580224 618248
rect 80796 591880 80848 591932
rect 84292 591880 84344 591932
rect 385684 590656 385736 590708
rect 579804 590656 579856 590708
rect 7564 589908 7616 589960
rect 96160 589908 96212 589960
rect 96436 589908 96488 589960
rect 96068 588548 96120 588600
rect 121736 588548 121788 588600
rect 92296 587868 92348 587920
rect 96068 587868 96120 587920
rect 97172 586576 97224 586628
rect 125968 586576 126020 586628
rect 106924 586508 106976 586560
rect 136824 586508 136876 586560
rect 47952 585760 48004 585812
rect 80796 585760 80848 585812
rect 47952 585216 48004 585268
rect 76012 585216 76064 585268
rect 85396 585216 85448 585268
rect 107016 585216 107068 585268
rect 34336 585148 34388 585200
rect 71964 585148 72016 585200
rect 75644 585148 75696 585200
rect 77392 585148 77444 585200
rect 101864 585080 101916 585132
rect 105544 585080 105596 585132
rect 113456 585148 113508 585200
rect 103888 584468 103940 584520
rect 106924 584468 106976 584520
rect 53564 584400 53616 584452
rect 81440 584400 81492 584452
rect 69664 584332 69716 584384
rect 70308 584332 70360 584384
rect 94872 584196 94924 584248
rect 97172 584196 97224 584248
rect 89628 583992 89680 584044
rect 123116 583992 123168 584044
rect 105728 583924 105780 583976
rect 118700 583924 118752 583976
rect 70308 583856 70360 583908
rect 77392 583856 77444 583908
rect 96528 583856 96580 583908
rect 114652 583856 114704 583908
rect 56416 583788 56468 583840
rect 83372 583788 83424 583840
rect 84108 583788 84160 583840
rect 96160 583788 96212 583840
rect 128636 583788 128688 583840
rect 49424 583720 49476 583772
rect 76748 583720 76800 583772
rect 102600 583720 102652 583772
rect 103428 583720 103480 583772
rect 106924 583720 106976 583772
rect 118700 583652 118752 583704
rect 119528 583652 119580 583704
rect 125692 583652 125744 583704
rect 80704 582972 80756 583024
rect 87696 582972 87748 583024
rect 56232 582564 56284 582616
rect 85120 582564 85172 582616
rect 53472 582496 53524 582548
rect 86224 582496 86276 582548
rect 91008 582496 91060 582548
rect 107108 582496 107160 582548
rect 39672 582428 39724 582480
rect 75736 582428 75788 582480
rect 87696 582428 87748 582480
rect 113364 582428 113416 582480
rect 41052 582360 41104 582412
rect 79968 582360 80020 582412
rect 92848 582360 92900 582412
rect 93768 582360 93820 582412
rect 124496 582360 124548 582412
rect 103704 581952 103756 582004
rect 69112 581884 69164 581936
rect 69756 581884 69808 581936
rect 70492 581816 70544 581868
rect 71780 581816 71832 581868
rect 57612 581612 57664 581664
rect 72424 581748 72476 581800
rect 101404 581748 101456 581800
rect 70216 581680 70268 581732
rect 73804 581680 73856 581732
rect 104440 581680 104492 581732
rect 105636 581680 105688 581732
rect 120172 581680 120224 581732
rect 121736 581476 121788 581528
rect 37004 581068 37056 581120
rect 70400 581068 70452 581120
rect 53564 581000 53616 581052
rect 70492 581000 70544 581052
rect 105636 581000 105688 581052
rect 114744 581000 114796 581052
rect 108028 580932 108080 580984
rect 122932 580932 122984 580984
rect 125876 580932 125928 580984
rect 108948 580864 109000 580916
rect 118700 580864 118752 580916
rect 105820 580252 105872 580304
rect 119344 580252 119396 580304
rect 35624 579640 35676 579692
rect 69664 579640 69716 579692
rect 59268 579572 59320 579624
rect 67640 579572 67692 579624
rect 108948 579572 109000 579624
rect 120356 579572 120408 579624
rect 121092 579572 121144 579624
rect 50896 578892 50948 578944
rect 59268 578892 59320 578944
rect 121092 578280 121144 578332
rect 123576 578280 123628 578332
rect 108672 578212 108724 578264
rect 140872 578212 140924 578264
rect 108120 578144 108172 578196
rect 125784 578144 125836 578196
rect 108948 577464 109000 577516
rect 116400 577464 116452 577516
rect 108672 576172 108724 576224
rect 116308 576172 116360 576224
rect 108764 576104 108816 576156
rect 142252 576104 142304 576156
rect 35808 575492 35860 575544
rect 67640 575492 67692 575544
rect 117136 575492 117188 575544
rect 126244 575492 126296 575544
rect 53840 574744 53892 574796
rect 55036 574744 55088 574796
rect 67640 574744 67692 574796
rect 105636 574472 105688 574524
rect 110420 574472 110472 574524
rect 48136 573996 48188 574048
rect 67640 573996 67692 574048
rect 108580 573996 108632 574048
rect 123024 573996 123076 574048
rect 108948 573928 109000 573980
rect 109684 573928 109736 573980
rect 43904 573384 43956 573436
rect 53840 573384 53892 573436
rect 32956 573316 33008 573368
rect 48136 573316 48188 573368
rect 109684 573316 109736 573368
rect 140964 573316 141016 573368
rect 108948 573180 109000 573232
rect 114560 573180 114612 573232
rect 108028 571956 108080 572008
rect 133972 571956 134024 572008
rect 134156 571956 134208 572008
rect 65892 571752 65944 571804
rect 66076 571752 66128 571804
rect 67640 571752 67692 571804
rect 64512 571276 64564 571328
rect 65892 571276 65944 571328
rect 67732 571276 67784 571328
rect 108304 571276 108356 571328
rect 128452 571276 128504 571328
rect 63224 571208 63276 571260
rect 67640 571208 67692 571260
rect 66168 569848 66220 569900
rect 66996 569848 67048 569900
rect 66996 568896 67048 568948
rect 67824 568896 67876 568948
rect 63224 568624 63276 568676
rect 67364 568624 67416 568676
rect 67640 568624 67692 568676
rect 108948 568556 109000 568608
rect 118608 568556 118660 568608
rect 108856 568488 108908 568540
rect 124404 568488 124456 568540
rect 125508 568488 125560 568540
rect 65984 568216 66036 568268
rect 67640 568216 67692 568268
rect 42800 567808 42852 567860
rect 43720 567808 43772 567860
rect 67640 567808 67692 567860
rect 125508 567808 125560 567860
rect 132592 567808 132644 567860
rect 30288 567196 30340 567248
rect 42800 567196 42852 567248
rect 60464 567196 60516 567248
rect 65984 567196 66036 567248
rect 108948 567196 109000 567248
rect 110512 567196 110564 567248
rect 113548 567196 113600 567248
rect 61936 566448 61988 566500
rect 67640 566448 67692 566500
rect 108948 566448 109000 566500
rect 128544 566448 128596 566500
rect 135168 566448 135220 566500
rect 142160 566448 142212 566500
rect 3240 565836 3292 565888
rect 25504 565836 25556 565888
rect 108948 565836 109000 565888
rect 134524 565836 134576 565888
rect 135168 565836 135220 565888
rect 108856 565768 108908 565820
rect 117412 565768 117464 565820
rect 44088 565088 44140 565140
rect 66904 565088 66956 565140
rect 67640 565088 67692 565140
rect 126244 565088 126296 565140
rect 497464 565088 497516 565140
rect 504364 565088 504416 565140
rect 42708 564340 42760 564392
rect 63500 564340 63552 564392
rect 67640 564408 67692 564460
rect 117412 564408 117464 564460
rect 119436 564408 119488 564460
rect 52368 564272 52420 564324
rect 67640 564272 67692 564324
rect 61844 564204 61896 564256
rect 67732 564204 67784 564256
rect 111708 564136 111760 564188
rect 113364 564136 113416 564188
rect 111156 563796 111208 563848
rect 114744 563796 114796 563848
rect 111248 563660 111300 563712
rect 116216 563660 116268 563712
rect 504364 563660 504416 563712
rect 580172 563660 580224 563712
rect 108948 563456 109000 563508
rect 111064 563456 111116 563508
rect 113824 563456 113876 563508
rect 60280 563184 60332 563236
rect 60648 563184 60700 563236
rect 60556 563116 60608 563168
rect 61384 563116 61436 563168
rect 49516 563048 49568 563100
rect 52368 563048 52420 563100
rect 60648 563048 60700 563100
rect 61844 563048 61896 563100
rect 53656 562300 53708 562352
rect 54484 562300 54536 562352
rect 67640 562300 67692 562352
rect 108948 562300 109000 562352
rect 142160 562300 142212 562352
rect 146300 562300 146352 562352
rect 48136 561620 48188 561672
rect 50804 561620 50856 561672
rect 67732 561620 67784 561672
rect 135904 561620 135956 561672
rect 136732 561620 136784 561672
rect 58992 561552 59044 561604
rect 60280 561552 60332 561604
rect 67640 561552 67692 561604
rect 108948 561008 109000 561060
rect 111800 561008 111852 561060
rect 117504 561008 117556 561060
rect 108856 560940 108908 560992
rect 135904 560940 135956 560992
rect 59084 560192 59136 560244
rect 59268 560192 59320 560244
rect 67640 560192 67692 560244
rect 112904 559580 112956 559632
rect 131304 559580 131356 559632
rect 42616 559512 42668 559564
rect 59268 559512 59320 559564
rect 108948 559512 109000 559564
rect 132500 559512 132552 559564
rect 132776 559512 132828 559564
rect 56416 558832 56468 558884
rect 58716 558832 58768 558884
rect 63408 558832 63460 558884
rect 64144 558832 64196 558884
rect 108028 558832 108080 558884
rect 139400 558832 139452 558884
rect 107752 558764 107804 558816
rect 111892 558764 111944 558816
rect 108948 558152 109000 558204
rect 121644 558152 121696 558204
rect 64144 557608 64196 557660
rect 67640 557608 67692 557660
rect 39948 557404 40000 557456
rect 50344 557540 50396 557592
rect 67732 557540 67784 557592
rect 49608 557472 49660 557524
rect 67824 557472 67876 557524
rect 56508 557404 56560 557456
rect 67640 557404 67692 557456
rect 108948 557132 109000 557184
rect 110604 557132 110656 557184
rect 34244 556860 34296 556912
rect 49608 556860 49660 556912
rect 39856 556792 39908 556844
rect 56508 556792 56560 556844
rect 110604 556792 110656 556844
rect 141056 556792 141108 556844
rect 56508 556180 56560 556232
rect 58624 556180 58676 556232
rect 67732 556112 67784 556164
rect 112996 555500 113048 555552
rect 119528 555500 119580 555552
rect 113088 555432 113140 555484
rect 113548 555432 113600 555484
rect 109776 555364 109828 555416
rect 121736 555364 121788 555416
rect 105636 555092 105688 555144
rect 105820 555092 105872 555144
rect 67640 554752 67692 554804
rect 108856 554752 108908 554804
rect 113272 554752 113324 554804
rect 114100 554752 114152 554804
rect 41236 554684 41288 554736
rect 62120 554684 62172 554736
rect 108948 554684 109000 554736
rect 129832 554684 129884 554736
rect 45468 554616 45520 554668
rect 48044 554616 48096 554668
rect 67640 554616 67692 554668
rect 129832 554072 129884 554124
rect 136732 554072 136784 554124
rect 108948 554004 109000 554056
rect 133972 554004 134024 554056
rect 3332 553392 3384 553444
rect 40684 553392 40736 553444
rect 67916 553392 67968 553444
rect 114100 553392 114152 553444
rect 116584 553392 116636 553444
rect 57612 553324 57664 553376
rect 57244 552644 57296 552696
rect 57888 552644 57940 552696
rect 67640 552644 67692 552696
rect 130200 552644 130252 552696
rect 138020 552644 138072 552696
rect 108948 552032 109000 552084
rect 130016 552032 130068 552084
rect 130200 552032 130252 552084
rect 64788 551964 64840 552016
rect 65616 551964 65668 552016
rect 67640 551964 67692 552016
rect 108304 551964 108356 552016
rect 143632 551964 143684 552016
rect 112628 551352 112680 551404
rect 116124 551352 116176 551404
rect 109684 551284 109736 551336
rect 117596 551284 117648 551336
rect 106740 551216 106792 551268
rect 111984 551216 112036 551268
rect 108948 550604 109000 550656
rect 59268 550536 59320 550588
rect 64604 550536 64656 550588
rect 67640 550536 67692 550588
rect 111064 550536 111116 550588
rect 115940 550536 115992 550588
rect 63132 549176 63184 549228
rect 63408 549176 63460 549228
rect 108948 549176 109000 549228
rect 132868 549176 132920 549228
rect 133788 549176 133840 549228
rect 109868 549108 109920 549160
rect 111156 549108 111208 549160
rect 63408 548564 63460 548616
rect 67640 548564 67692 548616
rect 133788 548564 133840 548616
rect 142344 548564 142396 548616
rect 108856 548496 108908 548548
rect 138664 548496 138716 548548
rect 143540 548496 143592 548548
rect 41144 547884 41196 547936
rect 67732 547884 67784 547936
rect 108948 547136 109000 547188
rect 135260 547136 135312 547188
rect 62028 546592 62080 546644
rect 64788 546592 64840 546644
rect 67640 546592 67692 546644
rect 60740 546456 60792 546508
rect 67640 546456 67692 546508
rect 108948 545640 109000 545692
rect 115204 545640 115256 545692
rect 38384 545096 38436 545148
rect 65984 545096 66036 545148
rect 67640 545096 67692 545148
rect 25504 545028 25556 545080
rect 68560 545028 68612 545080
rect 108948 544416 109000 544468
rect 116032 544416 116084 544468
rect 108856 544348 108908 544400
rect 139584 544348 139636 544400
rect 108856 543736 108908 543788
rect 109408 543736 109460 543788
rect 113272 543736 113324 543788
rect 139584 543736 139636 543788
rect 140780 543736 140832 543788
rect 60648 543668 60700 543720
rect 61752 543668 61804 543720
rect 67732 543668 67784 543720
rect 108948 543668 109000 543720
rect 129924 543668 129976 543720
rect 130752 543668 130804 543720
rect 60740 542988 60792 543040
rect 67640 542988 67692 543040
rect 130752 542988 130804 543040
rect 139400 542988 139452 543040
rect 34152 541628 34204 541680
rect 65524 541628 65576 541680
rect 67640 541628 67692 541680
rect 108856 540948 108908 541000
rect 110420 540948 110472 541000
rect 62028 540880 62080 540932
rect 63316 540880 63368 540932
rect 67640 540880 67692 540932
rect 108948 540880 109000 540932
rect 127164 540880 127216 540932
rect 131304 540880 131356 540932
rect 110420 540812 110472 540864
rect 111156 540812 111208 540864
rect 124312 540812 124364 540864
rect 37096 540336 37148 540388
rect 38568 540336 38620 540388
rect 48044 540200 48096 540252
rect 60096 540200 60148 540252
rect 60372 540200 60424 540252
rect 103704 539928 103756 539980
rect 122932 540200 122984 540252
rect 105544 539860 105596 539912
rect 105820 539860 105872 539912
rect 38476 539724 38528 539776
rect 45284 539724 45336 539776
rect 70492 539724 70544 539776
rect 60096 539656 60148 539708
rect 71964 539656 72016 539708
rect 38568 539588 38620 539640
rect 71320 539588 71372 539640
rect 108028 539588 108080 539640
rect 113180 539588 113232 539640
rect 40684 539520 40736 539572
rect 114560 539520 114612 539572
rect 115204 539520 115256 539572
rect 42708 539452 42760 539504
rect 45376 539452 45428 539504
rect 75184 539452 75236 539504
rect 97724 539452 97776 539504
rect 131764 539452 131816 539504
rect 132868 539588 132920 539640
rect 52368 539384 52420 539436
rect 77760 539384 77812 539436
rect 99656 539248 99708 539300
rect 100576 539248 100628 539300
rect 132684 539384 132736 539436
rect 104164 539316 104216 539368
rect 104716 539316 104768 539368
rect 120172 539316 120224 539368
rect 105636 538976 105688 539028
rect 105820 538976 105872 539028
rect 52092 538908 52144 538960
rect 73344 538908 73396 538960
rect 103244 538908 103296 538960
rect 106372 538908 106424 538960
rect 3424 538840 3476 538892
rect 93860 538840 93912 538892
rect 99288 538840 99340 538892
rect 111248 538840 111300 538892
rect 119344 538228 119396 538280
rect 125692 538228 125744 538280
rect 70124 538160 70176 538212
rect 86132 538160 86184 538212
rect 93860 538160 93912 538212
rect 98368 538160 98420 538212
rect 100300 538160 100352 538212
rect 128360 538160 128412 538212
rect 50712 538092 50764 538144
rect 80336 538092 80388 538144
rect 102232 538092 102284 538144
rect 131120 538092 131172 538144
rect 54944 538024 54996 538076
rect 83556 538024 83608 538076
rect 94504 538024 94556 538076
rect 119344 538024 119396 538076
rect 52276 537956 52328 538008
rect 78404 537956 78456 538008
rect 99012 537956 99064 538008
rect 121460 537956 121512 538008
rect 56324 537888 56376 537940
rect 73252 537888 73304 537940
rect 73344 537888 73396 537940
rect 80980 537888 81032 537940
rect 103520 537888 103572 537940
rect 122840 537888 122892 537940
rect 44088 537820 44140 537872
rect 74540 537820 74592 537872
rect 93216 537820 93268 537872
rect 93768 537820 93820 537872
rect 109776 537820 109828 537872
rect 43996 537548 44048 537600
rect 52276 537548 52328 537600
rect 89352 537548 89404 537600
rect 97908 537548 97960 537600
rect 103704 537548 103756 537600
rect 45376 537480 45428 537532
rect 56324 537480 56376 537532
rect 87420 537480 87472 537532
rect 99380 537480 99432 537532
rect 119436 537480 119488 537532
rect 142436 537480 142488 537532
rect 46480 536868 46532 536920
rect 50712 536868 50764 536920
rect 99472 536868 99524 536920
rect 100300 536868 100352 536920
rect 121460 536868 121512 536920
rect 124864 536868 124916 536920
rect 49608 536800 49660 536852
rect 54944 536800 54996 536852
rect 73344 536800 73396 536852
rect 73804 536800 73856 536852
rect 82820 536800 82872 536852
rect 83464 536800 83516 536852
rect 85488 536800 85540 536852
rect 97080 536800 97132 536852
rect 59176 536732 59228 536784
rect 91008 536732 91060 536784
rect 115848 536800 115900 536852
rect 121736 536800 121788 536852
rect 122840 536800 122892 536852
rect 123484 536800 123536 536852
rect 142436 536800 142488 536852
rect 580172 536800 580224 536852
rect 112260 536732 112312 536784
rect 50620 536664 50672 536716
rect 54760 536664 54812 536716
rect 82912 536664 82964 536716
rect 88064 536664 88116 536716
rect 57704 536596 57756 536648
rect 82820 536596 82872 536648
rect 93952 536596 94004 536648
rect 120080 536596 120132 536648
rect 98368 536528 98420 536580
rect 117320 536528 117372 536580
rect 95792 536460 95844 536512
rect 124220 536460 124272 536512
rect 112260 536324 112312 536376
rect 112904 536324 112956 536376
rect 113180 536324 113232 536376
rect 46848 536052 46900 536104
rect 51724 536052 51776 536104
rect 73896 536052 73948 536104
rect 120080 536052 120132 536104
rect 128452 536052 128504 536104
rect 117320 535440 117372 535492
rect 119344 535440 119396 535492
rect 124220 535440 124272 535492
rect 125784 535440 125836 535492
rect 39764 535372 39816 535424
rect 72608 535372 72660 535424
rect 92572 535372 92624 535424
rect 126980 535372 127032 535424
rect 130384 535372 130436 535424
rect 131120 535372 131172 535424
rect 53748 535304 53800 535356
rect 86776 535304 86828 535356
rect 100944 535304 100996 535356
rect 102048 535304 102100 535356
rect 133880 535304 133932 535356
rect 48228 535236 48280 535288
rect 79048 535236 79100 535288
rect 49332 535168 49384 535220
rect 79692 535168 79744 535220
rect 89996 534760 90048 534812
rect 114744 534760 114796 534812
rect 121552 534760 121604 534812
rect 96436 534692 96488 534744
rect 127164 534692 127216 534744
rect 129740 534692 129792 534744
rect 46664 534080 46716 534132
rect 48228 534080 48280 534132
rect 126980 534080 127032 534132
rect 131120 534080 131172 534132
rect 50988 534012 51040 534064
rect 55036 534012 55088 534064
rect 84844 534012 84896 534064
rect 102876 534012 102928 534064
rect 136640 534012 136692 534064
rect 57888 533944 57940 533996
rect 84200 533944 84252 533996
rect 89628 533468 89680 533520
rect 118884 533468 118936 533520
rect 56232 533400 56284 533452
rect 83556 533400 83608 533452
rect 95148 533400 95200 533452
rect 127256 533400 127308 533452
rect 42524 533332 42576 533384
rect 45284 533332 45336 533384
rect 76472 533332 76524 533384
rect 90640 533332 90692 533384
rect 124220 533332 124272 533384
rect 125600 533332 125652 533384
rect 91008 530680 91060 530732
rect 91928 530680 91980 530732
rect 109040 530680 109092 530732
rect 57336 530612 57388 530664
rect 77116 530612 77168 530664
rect 120724 530612 120776 530664
rect 45192 530544 45244 530596
rect 79324 530544 79376 530596
rect 91008 530544 91060 530596
rect 124496 530544 124548 530596
rect 46756 529864 46808 529916
rect 57336 529864 57388 529916
rect 3148 528504 3200 528556
rect 111064 528572 111116 528624
rect 3424 514768 3476 514820
rect 11704 514768 11756 514820
rect 431224 510620 431276 510672
rect 580172 510620 580224 510672
rect 11704 498788 11756 498840
rect 91100 498788 91152 498840
rect 86132 498176 86184 498228
rect 121460 498176 121512 498228
rect 3148 497428 3200 497480
rect 82912 497428 82964 497480
rect 96528 496068 96580 496120
rect 128636 496068 128688 496120
rect 132500 496068 132552 496120
rect 82820 495524 82872 495576
rect 83556 495524 83608 495576
rect 114560 495524 114612 495576
rect 85488 495388 85540 495440
rect 124312 495456 124364 495508
rect 128360 495456 128412 495508
rect 90640 494776 90692 494828
rect 114652 494776 114704 494828
rect 124312 494776 124364 494828
rect 56324 494708 56376 494760
rect 73804 494708 73856 494760
rect 95148 494708 95200 494760
rect 130108 494708 130160 494760
rect 134064 494708 134116 494760
rect 89996 494232 90048 494284
rect 96528 494232 96580 494284
rect 92480 494028 92532 494080
rect 93676 494028 93728 494080
rect 111800 494028 111852 494080
rect 82912 493960 82964 494012
rect 83556 493960 83608 494012
rect 120080 493960 120132 494012
rect 110420 493892 110472 493944
rect 111708 493892 111760 493944
rect 113916 493892 113968 493944
rect 88708 493824 88760 493876
rect 89628 493824 89680 493876
rect 80980 493348 81032 493400
rect 110420 493348 110472 493400
rect 120080 493348 120132 493400
rect 129924 493348 129976 493400
rect 82912 493280 82964 493332
rect 123116 493280 123168 493332
rect 127348 493280 127400 493332
rect 54852 492736 54904 492788
rect 55128 492736 55180 492788
rect 81900 492736 81952 492788
rect 47952 492600 48004 492652
rect 48228 492600 48280 492652
rect 53472 492600 53524 492652
rect 53656 492600 53708 492652
rect 58716 492600 58768 492652
rect 59176 492600 59228 492652
rect 77760 492600 77812 492652
rect 79324 492668 79376 492720
rect 114652 492804 114704 492856
rect 88708 492736 88760 492788
rect 110420 492736 110472 492788
rect 114468 492668 114520 492720
rect 129832 492668 129884 492720
rect 78404 492600 78456 492652
rect 82820 492600 82872 492652
rect 97816 492600 97868 492652
rect 98184 492600 98236 492652
rect 91100 492192 91152 492244
rect 131212 492192 131264 492244
rect 47860 492056 47912 492108
rect 49424 492056 49476 492108
rect 81624 492056 81676 492108
rect 92480 492056 92532 492108
rect 99656 492056 99708 492108
rect 112996 492056 113048 492108
rect 120172 492056 120224 492108
rect 70400 491988 70452 492040
rect 88064 491988 88116 492040
rect 99196 491988 99248 492040
rect 115940 491988 115992 492040
rect 41236 491920 41288 491972
rect 43812 491920 43864 491972
rect 71780 491920 71832 491972
rect 92572 491580 92624 491632
rect 99288 491580 99340 491632
rect 59176 491512 59228 491564
rect 76748 491512 76800 491564
rect 93216 491512 93268 491564
rect 100668 491512 100720 491564
rect 48228 491444 48280 491496
rect 70032 491444 70084 491496
rect 91928 491444 91980 491496
rect 95056 491444 95108 491496
rect 99196 491444 99248 491496
rect 109776 491444 109828 491496
rect 52276 491376 52328 491428
rect 74540 491376 74592 491428
rect 75460 491376 75512 491428
rect 97724 491376 97776 491428
rect 53656 491308 53708 491360
rect 80060 491308 80112 491360
rect 86776 491308 86828 491360
rect 91008 491308 91060 491360
rect 91744 491308 91796 491360
rect 96436 491308 96488 491360
rect 98184 491308 98236 491360
rect 98368 491376 98420 491428
rect 109868 491376 109920 491428
rect 110512 491308 110564 491360
rect 97908 491240 97960 491292
rect 102692 491240 102744 491292
rect 100668 491172 100720 491224
rect 127072 491240 127124 491292
rect 109132 491172 109184 491224
rect 109684 491172 109736 491224
rect 112536 491172 112588 491224
rect 91744 490628 91796 490680
rect 101404 490628 101456 490680
rect 39948 490560 40000 490612
rect 46572 490560 46624 490612
rect 72240 490560 72292 490612
rect 93768 490560 93820 490612
rect 103520 490560 103572 490612
rect 48964 489948 49016 490000
rect 74356 489948 74408 490000
rect 41052 489880 41104 489932
rect 73068 489880 73120 489932
rect 98184 489812 98236 489864
rect 99196 489812 99248 489864
rect 99288 489200 99340 489252
rect 107292 489200 107344 489252
rect 112628 489200 112680 489252
rect 99196 489132 99248 489184
rect 112444 489132 112496 489184
rect 67732 488520 67784 488572
rect 103428 488520 103480 488572
rect 117228 488520 117280 488572
rect 39672 488452 39724 488504
rect 42800 488452 42852 488504
rect 52184 488452 52236 488504
rect 67640 488452 67692 488504
rect 103336 488452 103388 488504
rect 123576 488520 123628 488572
rect 126980 488520 127032 488572
rect 52368 487772 52420 487824
rect 67640 487772 67692 487824
rect 103428 487228 103480 487280
rect 124128 487228 124180 487280
rect 104900 487160 104952 487212
rect 105728 487160 105780 487212
rect 147772 487160 147824 487212
rect 102784 487092 102836 487144
rect 140780 487092 140832 487144
rect 103336 487024 103388 487076
rect 104900 487024 104952 487076
rect 124128 487024 124180 487076
rect 125876 487024 125928 487076
rect 140780 486412 140832 486464
rect 152096 486412 152148 486464
rect 53840 485868 53892 485920
rect 67732 485868 67784 485920
rect 34336 485732 34388 485784
rect 36636 485800 36688 485852
rect 67640 485800 67692 485852
rect 41328 485732 41380 485784
rect 53840 485732 53892 485784
rect 102140 485120 102192 485172
rect 114468 485120 114520 485172
rect 53564 485052 53616 485104
rect 67640 485052 67692 485104
rect 102416 485052 102468 485104
rect 117228 485052 117280 485104
rect 64696 484372 64748 484424
rect 68468 484372 68520 484424
rect 117228 484372 117280 484424
rect 125600 484372 125652 484424
rect 286324 484372 286376 484424
rect 580172 484372 580224 484424
rect 35532 483624 35584 483676
rect 35716 483624 35768 483676
rect 67640 483624 67692 483676
rect 37004 482944 37056 482996
rect 68008 482944 68060 482996
rect 102140 482740 102192 482792
rect 105544 482740 105596 482792
rect 110604 482740 110656 482792
rect 115848 481720 115900 481772
rect 143724 481720 143776 481772
rect 40960 481652 41012 481704
rect 68928 481652 68980 481704
rect 102692 481652 102744 481704
rect 104900 481652 104952 481704
rect 107568 481652 107620 481704
rect 143540 481652 143592 481704
rect 102140 481584 102192 481636
rect 115204 481584 115256 481636
rect 115848 481584 115900 481636
rect 102232 481516 102284 481568
rect 107384 481516 107436 481568
rect 107568 481516 107620 481568
rect 66260 480836 66312 480888
rect 67640 480836 67692 480888
rect 61844 480156 61896 480208
rect 67548 480156 67600 480208
rect 102140 480156 102192 480208
rect 134156 480156 134208 480208
rect 35624 479476 35676 479528
rect 39672 479476 39724 479528
rect 66260 479476 66312 479528
rect 50896 478932 50948 478984
rect 52184 478932 52236 478984
rect 105544 478932 105596 478984
rect 115296 478932 115348 478984
rect 67640 478864 67692 478916
rect 107384 478864 107436 478916
rect 111156 478864 111208 478916
rect 134156 478864 134208 478916
rect 140872 478864 140924 478916
rect 118608 477572 118660 477624
rect 120080 477572 120132 477624
rect 61752 477504 61804 477556
rect 63040 477504 63092 477556
rect 67640 477504 67692 477556
rect 111892 477504 111944 477556
rect 113088 477504 113140 477556
rect 118700 477504 118752 477556
rect 103428 477436 103480 477488
rect 136916 477436 136968 477488
rect 102140 477368 102192 477420
rect 118608 477368 118660 477420
rect 102232 477300 102284 477352
rect 111892 477300 111944 477352
rect 38568 476076 38620 476128
rect 67640 476076 67692 476128
rect 102324 476008 102376 476060
rect 103336 476008 103388 476060
rect 139492 476008 139544 476060
rect 43904 475396 43956 475448
rect 67640 475396 67692 475448
rect 32956 475328 33008 475380
rect 67732 475328 67784 475380
rect 102140 475328 102192 475380
rect 132592 475328 132644 475380
rect 3424 474716 3476 474768
rect 11704 474716 11756 474768
rect 102140 474716 102192 474768
rect 121460 474716 121512 474768
rect 102232 474648 102284 474700
rect 134524 474648 134576 474700
rect 135444 474648 135496 474700
rect 121460 474580 121512 474632
rect 122748 474580 122800 474632
rect 128544 474580 128596 474632
rect 66076 473288 66128 473340
rect 67640 473288 67692 473340
rect 34336 472608 34388 472660
rect 66076 472608 66128 472660
rect 102140 472608 102192 472660
rect 142252 472608 142304 472660
rect 142436 472608 142488 472660
rect 102140 472064 102192 472116
rect 121460 472064 121512 472116
rect 102140 471928 102192 471980
rect 113824 471996 113876 472048
rect 133880 471996 133932 472048
rect 121460 471928 121512 471980
rect 138020 471928 138072 471980
rect 104072 471452 104124 471504
rect 107752 471452 107804 471504
rect 138020 471316 138072 471368
rect 148968 471316 149020 471368
rect 101956 471248 102008 471300
rect 135904 471248 135956 471300
rect 149244 471248 149296 471300
rect 65892 471044 65944 471096
rect 67088 471044 67140 471096
rect 67732 471044 67784 471096
rect 102140 470568 102192 470620
rect 148968 470568 149020 470620
rect 579988 470568 580040 470620
rect 139308 470500 139360 470552
rect 142160 470500 142212 470552
rect 66168 470432 66220 470484
rect 66996 470432 67048 470484
rect 67732 470432 67784 470484
rect 63316 470160 63368 470212
rect 67640 470160 67692 470212
rect 102140 469820 102192 469872
rect 117504 469820 117556 469872
rect 117504 469276 117556 469328
rect 117688 469276 117740 469328
rect 107476 469208 107528 469260
rect 145104 469208 145156 469260
rect 102140 469140 102192 469192
rect 60464 468460 60516 468512
rect 67640 468460 67692 468512
rect 64236 467916 64288 467968
rect 67640 467916 67692 467968
rect 106188 467848 106240 467900
rect 146484 467848 146536 467900
rect 61936 467780 61988 467832
rect 67456 467780 67508 467832
rect 102140 467780 102192 467832
rect 132776 467780 132828 467832
rect 137008 467780 137060 467832
rect 102232 467712 102284 467764
rect 106188 467712 106240 467764
rect 113916 467100 113968 467152
rect 128544 467100 128596 467152
rect 100576 466760 100628 466812
rect 101496 466760 101548 466812
rect 62764 466352 62816 466404
rect 63500 466352 63552 466404
rect 67640 466352 67692 466404
rect 100024 465740 100076 465792
rect 114744 465740 114796 465792
rect 54944 465672 54996 465724
rect 66904 465672 66956 465724
rect 67732 465672 67784 465724
rect 102324 465672 102376 465724
rect 141056 465672 141108 465724
rect 151912 465672 151964 465724
rect 102232 465060 102284 465112
rect 102140 464992 102192 465044
rect 107568 464992 107620 465044
rect 119988 464992 120040 465044
rect 121644 464992 121696 465044
rect 60556 464380 60608 464432
rect 67732 464380 67784 464432
rect 49516 464312 49568 464364
rect 67640 464312 67692 464364
rect 107568 464312 107620 464364
rect 143816 464312 143868 464364
rect 102140 463632 102192 463684
rect 116584 463632 116636 463684
rect 121460 463700 121512 463752
rect 117228 463632 117280 463684
rect 117504 463632 117556 463684
rect 106556 463360 106608 463412
rect 108304 463360 108356 463412
rect 54484 462952 54536 463004
rect 59084 462952 59136 463004
rect 106188 462952 106240 463004
rect 136732 462952 136784 463004
rect 146392 462952 146444 463004
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 59084 462340 59136 462392
rect 67640 462340 67692 462392
rect 102232 462272 102284 462324
rect 133972 462272 134024 462324
rect 141056 462272 141108 462324
rect 102140 462204 102192 462256
rect 106188 462204 106240 462256
rect 102140 460844 102192 460896
rect 106556 460912 106608 460964
rect 147680 460912 147732 460964
rect 48136 460164 48188 460216
rect 67640 460164 67692 460216
rect 102140 460164 102192 460216
rect 106096 460164 106148 460216
rect 130016 460164 130068 460216
rect 111064 459620 111116 459672
rect 119436 459620 119488 459672
rect 47676 459552 47728 459604
rect 48136 459552 48188 459604
rect 102232 459552 102284 459604
rect 103244 459552 103296 459604
rect 145012 459552 145064 459604
rect 63500 459484 63552 459536
rect 64144 459484 64196 459536
rect 67640 459484 67692 459536
rect 102140 459484 102192 459536
rect 111064 459484 111116 459536
rect 108304 458872 108356 458924
rect 135260 458872 135312 458924
rect 32956 458804 33008 458856
rect 63500 458804 63552 458856
rect 101312 458804 101364 458856
rect 138664 458804 138716 458856
rect 142528 458804 142580 458856
rect 50344 458124 50396 458176
rect 55864 458192 55916 458244
rect 67732 458192 67784 458244
rect 135260 458192 135312 458244
rect 136916 458192 136968 458244
rect 39856 457512 39908 457564
rect 50528 457512 50580 457564
rect 102232 457512 102284 457564
rect 108304 457512 108356 457564
rect 34244 457444 34296 457496
rect 36544 457444 36596 457496
rect 67640 457444 67692 457496
rect 103612 457444 103664 457496
rect 142344 457444 142396 457496
rect 150532 457444 150584 457496
rect 50528 456764 50580 456816
rect 50896 456764 50948 456816
rect 67640 456764 67692 456816
rect 108488 456764 108540 456816
rect 108948 456764 109000 456816
rect 150440 456764 150492 456816
rect 446404 456764 446456 456816
rect 580172 456764 580224 456816
rect 62120 456696 62172 456748
rect 67732 456696 67784 456748
rect 35716 456016 35768 456068
rect 62120 456016 62172 456068
rect 102876 456016 102928 456068
rect 121552 456016 121604 456068
rect 56508 455336 56560 455388
rect 57704 455336 57756 455388
rect 102140 455336 102192 455388
rect 108488 455336 108540 455388
rect 108948 454928 109000 454980
rect 111800 454928 111852 454980
rect 56508 454384 56560 454436
rect 57244 454384 57296 454436
rect 57704 454044 57756 454096
rect 67640 454044 67692 454096
rect 57612 453976 57664 454028
rect 68008 453976 68060 454028
rect 102140 453976 102192 454028
rect 139584 454044 139636 454096
rect 56508 453296 56560 453348
rect 67640 453296 67692 453348
rect 102876 453296 102928 453348
rect 118792 453296 118844 453348
rect 65616 452548 65668 452600
rect 67640 452548 67692 452600
rect 45468 451868 45520 451920
rect 46756 451868 46808 451920
rect 67364 451868 67416 451920
rect 102324 451868 102376 451920
rect 116032 451868 116084 451920
rect 116032 451528 116084 451580
rect 116584 451528 116636 451580
rect 30288 451256 30340 451308
rect 33784 451256 33836 451308
rect 58992 451256 59044 451308
rect 65616 451256 65668 451308
rect 102140 451256 102192 451308
rect 139400 451256 139452 451308
rect 67640 451188 67692 451240
rect 107384 449896 107436 449948
rect 138664 449896 138716 449948
rect 102140 449828 102192 449880
rect 102876 449216 102928 449268
rect 106188 449216 106240 449268
rect 107660 449216 107712 449268
rect 106004 448672 106056 448724
rect 123576 448672 123628 448724
rect 101588 448604 101640 448656
rect 107476 448604 107528 448656
rect 113272 448604 113324 448656
rect 3148 448536 3200 448588
rect 58624 448536 58676 448588
rect 59268 448536 59320 448588
rect 64144 448536 64196 448588
rect 67732 448536 67784 448588
rect 61936 448468 61988 448520
rect 63408 448468 63460 448520
rect 67640 448468 67692 448520
rect 102140 448468 102192 448520
rect 105636 448468 105688 448520
rect 106004 448468 106056 448520
rect 64788 447108 64840 447160
rect 65616 447108 65668 447160
rect 67640 447108 67692 447160
rect 102232 447108 102284 447160
rect 125876 447108 125928 447160
rect 131304 447108 131356 447160
rect 124220 446428 124272 446480
rect 124404 446428 124456 446480
rect 104808 445816 104860 445868
rect 112628 445816 112680 445868
rect 63132 445748 63184 445800
rect 67640 445748 67692 445800
rect 102600 445748 102652 445800
rect 135352 445748 135404 445800
rect 103244 445680 103296 445732
rect 104808 445680 104860 445732
rect 102508 445612 102560 445664
rect 104164 445612 104216 445664
rect 102232 445000 102284 445052
rect 136640 445000 136692 445052
rect 142160 445000 142212 445052
rect 55680 444320 55732 444372
rect 56416 444320 56468 444372
rect 67640 444320 67692 444372
rect 99656 444320 99708 444372
rect 123484 444388 123536 444440
rect 129740 444388 129792 444440
rect 41328 443640 41380 443692
rect 55680 443640 55732 443692
rect 60648 442892 60700 442944
rect 64604 442892 64656 442944
rect 37004 442688 37056 442740
rect 37188 442688 37240 442740
rect 37004 442212 37056 442264
rect 67640 442212 67692 442264
rect 102876 442212 102928 442264
rect 108764 442212 108816 442264
rect 130384 442212 130436 442264
rect 64604 441600 64656 441652
rect 67732 441600 67784 441652
rect 63408 441532 63460 441584
rect 99288 441532 99340 441584
rect 99380 441532 99432 441584
rect 65524 441464 65576 441516
rect 67640 441464 67692 441516
rect 62028 440852 62080 440904
rect 67640 440852 67692 440904
rect 117596 440852 117648 440904
rect 97908 440648 97960 440700
rect 102600 440308 102652 440360
rect 48044 440240 48096 440292
rect 50988 440240 51040 440292
rect 61844 440240 61896 440292
rect 62028 440240 62080 440292
rect 101496 440240 101548 440292
rect 102048 440240 102100 440292
rect 105544 440240 105596 440292
rect 133972 440240 134024 440292
rect 64696 439560 64748 439612
rect 75184 439560 75236 439612
rect 53748 439492 53800 439544
rect 82820 439492 82872 439544
rect 69112 439220 69164 439272
rect 71780 439220 71832 439272
rect 11704 439152 11756 439204
rect 96436 439152 96488 439204
rect 88708 439084 88760 439136
rect 121552 439084 121604 439136
rect 125508 439084 125560 439136
rect 132684 439084 132736 439136
rect 94504 439016 94556 439068
rect 128452 439016 128504 439068
rect 131488 439016 131540 439068
rect 39764 438948 39816 439000
rect 92480 438948 92532 439000
rect 93216 438948 93268 439000
rect 131120 438948 131172 439000
rect 72608 438880 72660 438932
rect 73344 438880 73396 438932
rect 119344 438880 119396 438932
rect 136824 438880 136876 438932
rect 4804 438812 4856 438864
rect 49608 438812 49660 438864
rect 99656 438812 99708 438864
rect 124864 438812 124916 438864
rect 125508 438812 125560 438864
rect 46664 438744 46716 438796
rect 78772 438744 78824 438796
rect 82820 438744 82872 438796
rect 83464 438744 83516 438796
rect 87420 438744 87472 438796
rect 91284 438744 91336 438796
rect 124220 438744 124272 438796
rect 124404 438744 124456 438796
rect 57888 438676 57940 438728
rect 82268 438676 82320 438728
rect 96436 438676 96488 438728
rect 125784 438676 125836 438728
rect 51724 438608 51776 438660
rect 73896 438608 73948 438660
rect 99012 438608 99064 438660
rect 119344 438608 119396 438660
rect 91008 438540 91060 438592
rect 100024 438540 100076 438592
rect 93860 438472 93912 438524
rect 95148 438472 95200 438524
rect 103520 438472 103572 438524
rect 58624 438404 58676 438456
rect 99748 438404 99800 438456
rect 45192 438268 45244 438320
rect 51724 438268 51776 438320
rect 45560 438200 45612 438252
rect 46204 438200 46256 438252
rect 73252 438200 73304 438252
rect 49608 438132 49660 438184
rect 50712 438132 50764 438184
rect 83556 438132 83608 438184
rect 89996 438132 90048 438184
rect 91008 438132 91060 438184
rect 97724 437996 97776 438048
rect 98644 437996 98696 438048
rect 86776 437452 86828 437504
rect 87604 437452 87656 437504
rect 97448 437384 97500 437436
rect 127164 437384 127216 437436
rect 46480 437316 46532 437368
rect 80980 437316 81032 437368
rect 88248 437316 88300 437368
rect 108396 437316 108448 437368
rect 50620 437248 50672 437300
rect 82912 437248 82964 437300
rect 88984 437248 89036 437300
rect 104900 437248 104952 437300
rect 43996 437180 44048 437232
rect 77944 437180 77996 437232
rect 78404 437180 78456 437232
rect 80152 436432 80204 436484
rect 80980 436432 81032 436484
rect 120264 436092 120316 436144
rect 120724 436092 120776 436144
rect 128452 436092 128504 436144
rect 45284 436024 45336 436076
rect 45468 436024 45520 436076
rect 76472 436024 76524 436076
rect 95056 436024 95108 436076
rect 125692 436024 125744 436076
rect 56324 435956 56376 436008
rect 81440 435956 81492 436008
rect 91928 435956 91980 436008
rect 120264 435956 120316 436008
rect 57336 435888 57388 435940
rect 76012 435888 76064 435940
rect 77116 435888 77168 435940
rect 48136 435344 48188 435396
rect 71320 435344 71372 435396
rect 42708 434664 42760 434716
rect 74724 434664 74776 434716
rect 75828 434664 75880 434716
rect 37096 434596 37148 434648
rect 47584 434596 47636 434648
rect 48136 434596 48188 434648
rect 43812 433236 43864 433288
rect 44088 433236 44140 433288
rect 74540 433236 74592 433288
rect 42708 432556 42760 432608
rect 70676 432556 70728 432608
rect 38476 431876 38528 431928
rect 42708 431876 42760 431928
rect 77944 431196 77996 431248
rect 580172 431196 580224 431248
rect 42064 430584 42116 430636
rect 42708 430584 42760 430636
rect 3424 429836 3476 429888
rect 101588 429836 101640 429888
rect 3516 422288 3568 422340
rect 120172 422220 120224 422272
rect 323584 418140 323636 418192
rect 580172 418140 580224 418192
rect 59176 410524 59228 410576
rect 89720 410524 89772 410576
rect 89720 409844 89772 409896
rect 353300 409844 353352 409896
rect 40960 406376 41012 406428
rect 71688 406376 71740 406428
rect 89812 406376 89864 406428
rect 114652 406376 114704 406428
rect 115848 406376 115900 406428
rect 92480 405016 92532 405068
rect 131304 405016 131356 405068
rect 106096 404948 106148 405000
rect 145196 404948 145248 405000
rect 544384 404336 544436 404388
rect 580172 404336 580224 404388
rect 36636 403588 36688 403640
rect 75920 403588 75972 403640
rect 75920 403044 75972 403096
rect 164884 403044 164936 403096
rect 67456 402976 67508 403028
rect 367100 402976 367152 403028
rect 64788 401616 64840 401668
rect 162124 401616 162176 401668
rect 35532 400936 35584 400988
rect 70400 400936 70452 400988
rect 34428 400868 34480 400920
rect 42800 400868 42852 400920
rect 80060 400868 80112 400920
rect 70400 400256 70452 400308
rect 74540 400256 74592 400308
rect 153844 400256 153896 400308
rect 80060 400188 80112 400240
rect 80244 400188 80296 400240
rect 320272 400188 320324 400240
rect 49424 399576 49476 399628
rect 81440 399576 81492 399628
rect 52276 399508 52328 399560
rect 88064 399508 88116 399560
rect 41052 399440 41104 399492
rect 84936 399440 84988 399492
rect 95884 399440 95936 399492
rect 108856 399440 108908 399492
rect 160744 399440 160796 399492
rect 87696 398964 87748 399016
rect 88064 398964 88116 399016
rect 159364 398964 159416 399016
rect 68652 398896 68704 398948
rect 228364 398896 228416 398948
rect 106280 398828 106332 398880
rect 106924 398828 106976 398880
rect 358820 398828 358872 398880
rect 109868 398760 109920 398812
rect 114100 398760 114152 398812
rect 53472 398148 53524 398200
rect 85764 398148 85816 398200
rect 95056 398148 95108 398200
rect 119620 398148 119672 398200
rect 52000 398080 52052 398132
rect 87604 398080 87656 398132
rect 88340 398080 88392 398132
rect 122840 398080 122892 398132
rect 157984 398080 158036 398132
rect 42616 397400 42668 397452
rect 69204 397400 69256 397452
rect 268384 397468 268436 397520
rect 107476 396856 107528 396908
rect 129832 396856 129884 396908
rect 57796 396788 57848 396840
rect 83464 396788 83516 396840
rect 97816 396788 97868 396840
rect 127256 396788 127308 396840
rect 46848 396720 46900 396772
rect 78772 396720 78824 396772
rect 93952 396720 94004 396772
rect 128544 396720 128596 396772
rect 154672 396720 154724 396772
rect 108304 396652 108356 396704
rect 114560 396652 114612 396704
rect 129832 396108 129884 396160
rect 130016 396108 130068 396160
rect 289084 396108 289136 396160
rect 46756 395972 46808 396024
rect 55956 396040 56008 396092
rect 286324 396040 286376 396092
rect 96712 395292 96764 395344
rect 130200 395292 130252 395344
rect 149152 395292 149204 395344
rect 39304 394748 39356 394800
rect 115848 394748 115900 394800
rect 118792 394748 118844 394800
rect 119988 394748 120040 394800
rect 122840 394748 122892 394800
rect 291844 394748 291896 394800
rect 385684 394748 385736 394800
rect 55864 394680 55916 394732
rect 64696 394680 64748 394732
rect 151820 394680 151872 394732
rect 304264 394680 304316 394732
rect 68744 394612 68796 394664
rect 68928 394612 68980 394664
rect 115848 394612 115900 394664
rect 118792 394612 118844 394664
rect 52092 394068 52144 394120
rect 74724 394068 74776 394120
rect 110512 394068 110564 394120
rect 130108 394068 130160 394120
rect 138112 394068 138164 394120
rect 54760 394000 54812 394052
rect 82820 394000 82872 394052
rect 100668 394000 100720 394052
rect 107660 394000 107712 394052
rect 108764 394000 108816 394052
rect 131396 394000 131448 394052
rect 47860 393932 47912 393984
rect 81440 393932 81492 393984
rect 95792 393932 95844 393984
rect 127348 393932 127400 393984
rect 152004 393932 152056 393984
rect 83004 393456 83056 393508
rect 146944 393456 146996 393508
rect 131396 393388 131448 393440
rect 316684 393388 316736 393440
rect 68928 393320 68980 393372
rect 278044 393320 278096 393372
rect 46756 392640 46808 392692
rect 77300 392640 77352 392692
rect 106188 392640 106240 392692
rect 131212 392640 131264 392692
rect 3424 392572 3476 392624
rect 52460 392572 52512 392624
rect 56416 392572 56468 392624
rect 86224 392572 86276 392624
rect 91008 392572 91060 392624
rect 120264 392572 120316 392624
rect 146300 392572 146352 392624
rect 116676 392436 116728 392488
rect 118700 392436 118752 392488
rect 43996 392164 44048 392216
rect 88984 392164 89036 392216
rect 101036 392164 101088 392216
rect 101404 392164 101456 392216
rect 135260 392164 135312 392216
rect 82912 392096 82964 392148
rect 83648 392096 83700 392148
rect 140044 392096 140096 392148
rect 67364 392028 67416 392080
rect 143632 392028 143684 392080
rect 52460 391960 52512 392012
rect 53656 391960 53708 392012
rect 116676 391960 116728 392012
rect 120264 391960 120316 392012
rect 120816 391960 120868 392012
rect 220084 391960 220136 392012
rect 41236 391892 41288 391944
rect 82912 391892 82964 391944
rect 59084 391824 59136 391876
rect 67364 391824 67416 391876
rect 53564 391212 53616 391264
rect 75460 391212 75512 391264
rect 88984 391212 89036 391264
rect 103612 391212 103664 391264
rect 110328 391212 110380 391264
rect 134064 391212 134116 391264
rect 140780 391212 140832 391264
rect 50988 390668 51040 390720
rect 79324 390668 79376 390720
rect 114100 390668 114152 390720
rect 133144 390668 133196 390720
rect 75460 390600 75512 390652
rect 134064 390600 134116 390652
rect 57704 390464 57756 390516
rect 324412 390532 324464 390584
rect 109776 390124 109828 390176
rect 114928 390124 114980 390176
rect 103336 390056 103388 390108
rect 115204 390056 115256 390108
rect 114468 389920 114520 389972
rect 124312 389920 124364 389972
rect 128544 389920 128596 389972
rect 115848 389852 115900 389904
rect 120172 389852 120224 389904
rect 147864 389852 147916 389904
rect 41236 389784 41288 389836
rect 73344 389784 73396 389836
rect 99288 389784 99340 389836
rect 128360 389784 128412 389836
rect 119436 389580 119488 389632
rect 120908 389580 120960 389632
rect 71688 389308 71740 389360
rect 73344 389308 73396 389360
rect 49608 389172 49660 389224
rect 53840 389172 53892 389224
rect 55036 389172 55088 389224
rect 95516 389172 95568 389224
rect 128360 389172 128412 389224
rect 130384 389172 130436 389224
rect 103612 389104 103664 389156
rect 110420 389104 110472 389156
rect 112536 388628 112588 388680
rect 121552 388628 121604 388680
rect 53840 388560 53892 388612
rect 77484 388560 77536 388612
rect 94872 388560 94924 388612
rect 102232 388560 102284 388612
rect 104624 388560 104676 388612
rect 114468 388560 114520 388612
rect 69664 388492 69716 388544
rect 88892 388492 88944 388544
rect 102600 388492 102652 388544
rect 115940 388492 115992 388544
rect 159456 388492 159508 388544
rect 52368 388424 52420 388476
rect 77300 388424 77352 388476
rect 110420 388424 110472 388476
rect 309140 388424 309192 388476
rect 77300 388016 77352 388068
rect 78496 388016 78548 388068
rect 95424 388084 95476 388136
rect 92848 388016 92900 388068
rect 95884 388016 95936 388068
rect 52276 387948 52328 388000
rect 69756 387948 69808 388000
rect 81440 387948 81492 388000
rect 82544 387948 82596 388000
rect 86960 387948 87012 388000
rect 93308 387948 93360 388000
rect 119344 387948 119396 388000
rect 53748 387880 53800 387932
rect 87052 387880 87104 387932
rect 91560 387880 91612 387932
rect 108304 387880 108356 387932
rect 114928 387880 114980 387932
rect 184204 387880 184256 387932
rect 4804 387812 4856 387864
rect 71780 387812 71832 387864
rect 72700 387812 72752 387864
rect 119436 387812 119488 387864
rect 121552 387812 121604 387864
rect 244924 387812 244976 387864
rect 57796 387744 57848 387796
rect 58624 387744 58676 387796
rect 107660 387744 107712 387796
rect 108488 387744 108540 387796
rect 39948 387200 40000 387252
rect 57244 387200 57296 387252
rect 57796 387200 57848 387252
rect 77944 387200 77996 387252
rect 52184 387132 52236 387184
rect 80152 387132 80204 387184
rect 86960 387132 87012 387184
rect 154580 387132 154632 387184
rect 38476 387064 38528 387116
rect 110604 387064 110656 387116
rect 115940 387064 115992 387116
rect 108488 386588 108540 386640
rect 123668 386588 123720 386640
rect 57244 386520 57296 386572
rect 84476 386520 84528 386572
rect 112168 386520 112220 386572
rect 112444 386520 112496 386572
rect 167644 386520 167696 386572
rect 48228 386452 48280 386504
rect 80612 386452 80664 386504
rect 107200 386452 107252 386504
rect 127072 386452 127124 386504
rect 154580 386452 154632 386504
rect 321560 386452 321612 386504
rect 323584 386384 323636 386436
rect 58992 386316 59044 386368
rect 60004 386316 60056 386368
rect 54852 385704 54904 385756
rect 76012 386112 76064 386164
rect 106096 386044 106148 386096
rect 53564 385636 53616 385688
rect 84292 385976 84344 386028
rect 108304 385976 108356 386028
rect 121552 385976 121604 386028
rect 134156 385704 134208 385756
rect 95424 385636 95476 385688
rect 128360 385636 128412 385688
rect 39672 385092 39724 385144
rect 71780 385296 71832 385348
rect 48136 385024 48188 385076
rect 53748 385024 53800 385076
rect 92940 385296 92992 385348
rect 104440 385296 104492 385348
rect 121552 385092 121604 385144
rect 263600 385092 263652 385144
rect 122656 385024 122708 385076
rect 61752 384956 61804 385008
rect 67640 384956 67692 385008
rect 128360 385024 128412 385076
rect 301504 385024 301556 385076
rect 132500 384956 132552 385008
rect 118516 384752 118568 384804
rect 124312 384752 124364 384804
rect 60648 384480 60700 384532
rect 61752 384480 61804 384532
rect 118608 384344 118660 384396
rect 124128 384344 124180 384396
rect 127164 384344 127216 384396
rect 39948 383664 40000 383716
rect 68744 383664 68796 383716
rect 126888 383120 126940 383172
rect 147772 383120 147824 383172
rect 118608 383052 118660 383104
rect 125508 383052 125560 383104
rect 119436 382984 119488 383036
rect 147772 382984 147824 383036
rect 124312 382916 124364 382968
rect 349804 382916 349856 382968
rect 125508 382644 125560 382696
rect 126980 382644 127032 382696
rect 42708 382236 42760 382288
rect 67640 382236 67692 382288
rect 147772 382236 147824 382288
rect 209780 382236 209832 382288
rect 118608 382168 118660 382220
rect 152096 382168 152148 382220
rect 153108 382168 153160 382220
rect 118608 381556 118660 381608
rect 126244 381556 126296 381608
rect 126888 381556 126940 381608
rect 116400 381488 116452 381540
rect 125600 381488 125652 381540
rect 137284 381488 137336 381540
rect 153108 381488 153160 381540
rect 181444 381488 181496 381540
rect 42800 380128 42852 380180
rect 43904 380128 43956 380180
rect 67916 380128 67968 380180
rect 118332 380128 118384 380180
rect 189724 380128 189776 380180
rect 3424 378768 3476 378820
rect 42800 378768 42852 378820
rect 130384 378768 130436 378820
rect 163504 378768 163556 378820
rect 118608 378700 118660 378752
rect 124128 378700 124180 378752
rect 118056 378156 118108 378208
rect 129832 378156 129884 378208
rect 213184 378156 213236 378208
rect 346400 378156 346452 378208
rect 353944 378156 353996 378208
rect 580172 378156 580224 378208
rect 118240 378088 118292 378140
rect 140964 378088 141016 378140
rect 141240 378088 141292 378140
rect 141240 377408 141292 377460
rect 155960 377408 156012 377460
rect 171784 376864 171836 376916
rect 305644 376864 305696 376916
rect 155960 376796 156012 376848
rect 313280 376796 313332 376848
rect 34336 376660 34388 376712
rect 65524 376728 65576 376780
rect 67640 376728 67692 376780
rect 263600 376728 263652 376780
rect 520924 376728 520976 376780
rect 66168 376660 66220 376712
rect 67732 376660 67784 376712
rect 118148 376660 118200 376712
rect 143540 376660 143592 376712
rect 149060 376660 149112 376712
rect 119344 376048 119396 376100
rect 297364 376048 297416 376100
rect 313280 376048 313332 376100
rect 318800 376048 318852 376100
rect 133788 375980 133840 376032
rect 143724 375980 143776 376032
rect 331220 375980 331272 376032
rect 233884 375436 233936 375488
rect 347780 375436 347832 375488
rect 62028 375368 62080 375420
rect 67088 375368 67140 375420
rect 67640 375368 67692 375420
rect 118608 375368 118660 375420
rect 132592 375368 132644 375420
rect 133788 375368 133840 375420
rect 217968 375368 218020 375420
rect 339500 375368 339552 375420
rect 138664 375300 138716 375352
rect 141148 375300 141200 375352
rect 63316 374620 63368 374672
rect 67640 374620 67692 374672
rect 129832 374620 129884 374672
rect 265624 374620 265676 374672
rect 253204 374144 253256 374196
rect 357440 374144 357492 374196
rect 141148 374076 141200 374128
rect 327264 374076 327316 374128
rect 209780 374008 209832 374060
rect 471980 374008 472032 374060
rect 60464 373940 60516 373992
rect 67732 373940 67784 373992
rect 118608 373940 118660 373992
rect 140872 373940 140924 373992
rect 64788 373260 64840 373312
rect 67640 373260 67692 373312
rect 140872 373260 140924 373312
rect 185584 373260 185636 373312
rect 220084 372988 220136 373040
rect 220728 372988 220780 373040
rect 170404 372784 170456 372836
rect 327172 372784 327224 372836
rect 117872 372716 117924 372768
rect 284300 372716 284352 372768
rect 220728 372648 220780 372700
rect 403624 372648 403676 372700
rect 59268 372580 59320 372632
rect 60464 372580 60516 372632
rect 198004 372580 198056 372632
rect 411904 372580 411956 372632
rect 3516 372512 3568 372564
rect 39304 372512 39356 372564
rect 123576 371968 123628 372020
rect 138020 371968 138072 372020
rect 139032 371968 139084 372020
rect 115848 371900 115900 371952
rect 141056 371900 141108 371952
rect 120080 371832 120132 371884
rect 135444 371832 135496 371884
rect 139492 371832 139544 371884
rect 339592 371832 339644 371884
rect 139032 371356 139084 371408
rect 135904 371288 135956 371340
rect 139492 371288 139544 371340
rect 342260 371288 342312 371340
rect 117780 371220 117832 371272
rect 338764 371220 338816 371272
rect 54944 370472 54996 370524
rect 67640 370472 67692 370524
rect 118608 370472 118660 370524
rect 120172 370472 120224 370524
rect 129832 370472 129884 370524
rect 284300 370472 284352 370524
rect 337384 370472 337436 370524
rect 249708 370132 249760 370184
rect 324964 370132 325016 370184
rect 169116 370064 169168 370116
rect 282920 370064 282972 370116
rect 174636 369996 174688 370048
rect 295340 369996 295392 370048
rect 212908 369928 212960 369980
rect 417424 369928 417476 369980
rect 37188 369860 37240 369912
rect 223488 369860 223540 369912
rect 464344 369860 464396 369912
rect 62764 369792 62816 369844
rect 67640 369792 67692 369844
rect 118424 369792 118476 369844
rect 132500 369792 132552 369844
rect 141424 369792 141476 369844
rect 121000 369180 121052 369232
rect 125876 369180 125928 369232
rect 60372 369112 60424 369164
rect 69664 369112 69716 369164
rect 118700 369112 118752 369164
rect 255320 369112 255372 369164
rect 258724 368772 258776 368824
rect 343640 368772 343692 368824
rect 194048 368704 194100 368756
rect 333980 368704 334032 368756
rect 119344 368636 119396 368688
rect 270224 368636 270276 368688
rect 282920 368636 282972 368688
rect 335452 368636 335504 368688
rect 160836 368568 160888 368620
rect 323124 368568 323176 368620
rect 49516 368500 49568 368552
rect 53656 368500 53708 368552
rect 67640 368500 67692 368552
rect 255320 368500 255372 368552
rect 457444 368500 457496 368552
rect 117780 367820 117832 367872
rect 120080 367820 120132 367872
rect 118608 367752 118660 367804
rect 122748 367752 122800 367804
rect 126428 367752 126480 367804
rect 269856 367412 269908 367464
rect 270224 367412 270276 367464
rect 340880 367412 340932 367464
rect 286324 367344 286376 367396
rect 286600 367344 286652 367396
rect 371884 367344 371936 367396
rect 166264 367276 166316 367328
rect 300124 367276 300176 367328
rect 182916 367208 182968 367260
rect 324504 367208 324556 367260
rect 126336 367140 126388 367192
rect 293224 367140 293276 367192
rect 295340 367140 295392 367192
rect 295616 367140 295668 367192
rect 350540 367140 350592 367192
rect 123484 367072 123536 367124
rect 321836 367072 321888 367124
rect 59084 367004 59136 367056
rect 67640 367004 67692 367056
rect 118148 367004 118200 367056
rect 142252 367004 142304 367056
rect 144920 367004 144972 367056
rect 189816 366052 189868 366104
rect 247040 366052 247092 366104
rect 275928 366052 275980 366104
rect 320180 366052 320232 366104
rect 176108 365984 176160 366036
rect 209044 365984 209096 366036
rect 244924 365984 244976 366036
rect 358084 365984 358136 366036
rect 162216 365916 162268 365968
rect 323032 365916 323084 365968
rect 169208 365848 169260 365900
rect 238668 365848 238720 365900
rect 297364 365848 297416 365900
rect 475384 365848 475436 365900
rect 146944 365780 146996 365832
rect 327080 365780 327132 365832
rect 124956 365712 125008 365764
rect 312728 365712 312780 365764
rect 118056 365644 118108 365696
rect 133880 365644 133932 365696
rect 196808 364692 196860 364744
rect 216588 364692 216640 364744
rect 181536 364624 181588 364676
rect 242256 364624 242308 364676
rect 309968 364624 310020 364676
rect 325792 364624 325844 364676
rect 195428 364556 195480 364608
rect 227720 364556 227772 364608
rect 171876 364488 171928 364540
rect 236092 364488 236144 364540
rect 335360 364556 335412 364608
rect 257344 364488 257396 364540
rect 395344 364488 395396 364540
rect 119528 364420 119580 364472
rect 258724 364420 258776 364472
rect 265624 364420 265676 364472
rect 414664 364420 414716 364472
rect 43904 364352 43956 364404
rect 47676 364352 47728 364404
rect 117320 364352 117372 364404
rect 67640 364284 67692 364336
rect 148968 364352 149020 364404
rect 153200 364352 153252 364404
rect 198648 364352 198700 364404
rect 579620 364352 579672 364404
rect 118148 364216 118200 364268
rect 139308 364216 139360 364268
rect 187056 363196 187108 363248
rect 206468 363196 206520 363248
rect 305644 363196 305696 363248
rect 306288 363196 306340 363248
rect 320824 363196 320876 363248
rect 191104 363128 191156 363180
rect 225788 363128 225840 363180
rect 242256 363128 242308 363180
rect 351920 363128 351972 363180
rect 195336 363060 195388 363112
rect 321652 363060 321704 363112
rect 192484 362992 192536 363044
rect 233884 362992 233936 363044
rect 268384 362992 268436 363044
rect 466460 362992 466512 363044
rect 35532 362924 35584 362976
rect 69204 362924 69256 362976
rect 123576 362924 123628 362976
rect 213184 362924 213236 362976
rect 216588 362924 216640 362976
rect 510620 362924 510672 362976
rect 64696 362856 64748 362908
rect 67640 362856 67692 362908
rect 117964 362856 118016 362908
rect 149244 362856 149296 362908
rect 217416 362856 217468 362908
rect 228364 362856 228416 362908
rect 229652 362856 229704 362908
rect 316684 362448 316736 362500
rect 317328 362448 317380 362500
rect 199384 362312 199436 362364
rect 249708 362312 249760 362364
rect 250904 362312 250956 362364
rect 149244 362244 149296 362296
rect 175924 362244 175976 362296
rect 196624 362244 196676 362296
rect 275928 362244 275980 362296
rect 276664 362244 276716 362296
rect 117688 362176 117740 362228
rect 144276 362176 144328 362228
rect 166356 362176 166408 362228
rect 309968 362176 310020 362228
rect 213184 362108 213236 362160
rect 214840 362108 214892 362160
rect 217968 362040 218020 362092
rect 219348 362040 219400 362092
rect 258724 361904 258776 361956
rect 259920 361904 259972 361956
rect 289176 361904 289228 361956
rect 319444 361904 319496 361956
rect 281172 361836 281224 361888
rect 360844 361836 360896 361888
rect 310796 361768 310848 361820
rect 399484 361768 399536 361820
rect 225788 361700 225840 361752
rect 317052 361700 317104 361752
rect 184848 361632 184900 361684
rect 202604 361632 202656 361684
rect 249708 361632 249760 361684
rect 345664 361632 345716 361684
rect 143724 361564 143776 361616
rect 144276 361564 144328 361616
rect 240600 361564 240652 361616
rect 145104 361496 145156 361548
rect 281172 361564 281224 361616
rect 301504 361564 301556 361616
rect 410524 361564 410576 361616
rect 32956 360816 33008 360868
rect 42800 360816 42852 360868
rect 118608 360816 118660 360868
rect 121644 360816 121696 360868
rect 145104 360816 145156 360868
rect 308496 360816 308548 360868
rect 309140 360816 309192 360868
rect 356704 360816 356756 360868
rect 119436 360544 119488 360596
rect 314660 360544 314712 360596
rect 278136 360476 278188 360528
rect 278596 360476 278648 360528
rect 352564 360476 352616 360528
rect 199476 360408 199528 360460
rect 310796 360408 310848 360460
rect 196716 360340 196768 360392
rect 257344 360340 257396 360392
rect 272156 360340 272208 360392
rect 406384 360340 406436 360392
rect 133144 360272 133196 360324
rect 324320 360272 324372 360324
rect 42800 360204 42852 360256
rect 44088 360204 44140 360256
rect 67640 360204 67692 360256
rect 198832 360204 198884 360256
rect 204536 360204 204588 360256
rect 312728 360204 312780 360256
rect 322940 360204 322992 360256
rect 118148 360136 118200 360188
rect 146484 360136 146536 360188
rect 317512 359592 317564 359644
rect 319536 359592 319588 359644
rect 50896 359524 50948 359576
rect 67640 359524 67692 359576
rect 36544 359456 36596 359508
rect 41052 359456 41104 359508
rect 67732 359456 67784 359508
rect 118608 359456 118660 359508
rect 120724 359456 120776 359508
rect 137008 359456 137060 359508
rect 212540 359388 212592 359440
rect 193956 358912 194008 358964
rect 199844 358912 199896 358964
rect 314844 359388 314896 359440
rect 320364 359388 320416 359440
rect 321652 358912 321704 358964
rect 167736 358844 167788 358896
rect 329840 358844 329892 358896
rect 320364 358776 320416 358828
rect 495440 358776 495492 358828
rect 118056 358708 118108 358760
rect 121000 358708 121052 358760
rect 125508 358708 125560 358760
rect 128636 358708 128688 358760
rect 57704 358028 57756 358080
rect 67640 358028 67692 358080
rect 118608 358028 118660 358080
rect 122840 358028 122892 358080
rect 146944 358028 146996 358080
rect 198832 358028 198884 358080
rect 319536 358028 319588 358080
rect 469220 358028 469272 358080
rect 3148 357416 3200 357468
rect 15844 357416 15896 357468
rect 128636 357416 128688 357468
rect 198004 357416 198056 357468
rect 35716 357348 35768 357400
rect 66904 357348 66956 357400
rect 67548 357348 67600 357400
rect 150624 357348 150676 357400
rect 151912 357348 151964 357400
rect 199844 357348 199896 357400
rect 118608 356736 118660 356788
rect 186964 356736 187016 356788
rect 124864 356668 124916 356720
rect 198280 356668 198332 356720
rect 198648 356668 198700 356720
rect 41144 356056 41196 356108
rect 68008 356056 68060 356108
rect 118608 356056 118660 356108
rect 150624 356056 150676 356108
rect 118516 355988 118568 356040
rect 143816 355988 143868 356040
rect 144828 355988 144880 356040
rect 56508 355376 56560 355428
rect 67640 355376 67692 355428
rect 55956 355308 56008 355360
rect 67732 355308 67784 355360
rect 144828 355308 144880 355360
rect 182824 355308 182876 355360
rect 319904 355308 319956 355360
rect 458180 355308 458232 355360
rect 135168 354628 135220 354680
rect 146392 354628 146444 354680
rect 198188 354628 198240 354680
rect 118608 354356 118660 354408
rect 121460 354356 121512 354408
rect 322848 354356 322900 354408
rect 324504 354356 324556 354408
rect 117780 354016 117832 354068
rect 133880 354016 133932 354068
rect 135168 354016 135220 354068
rect 121460 353948 121512 354000
rect 142252 353948 142304 354000
rect 196808 353948 196860 354000
rect 508504 353948 508556 354000
rect 579620 353948 579672 354000
rect 60004 353200 60056 353252
rect 66996 353200 67048 353252
rect 67548 353200 67600 353252
rect 41420 352520 41472 352572
rect 42616 352520 42668 352572
rect 68928 352520 68980 352572
rect 126428 352520 126480 352572
rect 140136 352520 140188 352572
rect 21364 351908 21416 351960
rect 41420 351908 41472 351960
rect 61660 351840 61712 351892
rect 64144 351840 64196 351892
rect 67640 351840 67692 351892
rect 117412 351840 117464 351892
rect 147680 351840 147732 351892
rect 118608 351772 118660 351824
rect 145196 351772 145248 351824
rect 147680 351160 147732 351212
rect 178684 351160 178736 351212
rect 319444 351160 319496 351212
rect 452660 351160 452712 351212
rect 118608 350480 118660 350532
rect 120908 350548 120960 350600
rect 132776 350548 132828 350600
rect 141424 350548 141476 350600
rect 142436 350548 142488 350600
rect 197360 350548 197412 350600
rect 322664 349800 322716 349852
rect 323124 349800 323176 349852
rect 489184 349800 489236 349852
rect 61936 349120 61988 349172
rect 64696 349120 64748 349172
rect 67640 349120 67692 349172
rect 35624 349052 35676 349104
rect 69664 349052 69716 349104
rect 118608 349052 118660 349104
rect 145012 349052 145064 349104
rect 146208 349052 146260 349104
rect 63132 348984 63184 349036
rect 65616 348984 65668 349036
rect 67640 348984 67692 349036
rect 118516 348984 118568 349036
rect 142344 348984 142396 349036
rect 143448 348984 143500 349036
rect 322204 348372 322256 348424
rect 334624 348372 334676 348424
rect 63224 347692 63276 347744
rect 66168 347692 66220 347744
rect 67640 347692 67692 347744
rect 118608 347012 118660 347064
rect 132592 347012 132644 347064
rect 133788 347012 133840 347064
rect 322296 347012 322348 347064
rect 356060 347012 356112 347064
rect 133788 346468 133840 346520
rect 180064 346468 180116 346520
rect 179328 346400 179380 346452
rect 197360 346400 197412 346452
rect 15844 346332 15896 346384
rect 68836 346332 68888 346384
rect 116584 346332 116636 346384
rect 117320 346332 117372 346384
rect 118608 346332 118660 346384
rect 136916 346332 136968 346384
rect 137192 346332 137244 346384
rect 2780 346264 2832 346316
rect 4804 346264 4856 346316
rect 137192 345652 137244 345704
rect 180156 345652 180208 345704
rect 45284 345040 45336 345092
rect 68652 345040 68704 345092
rect 118516 345040 118568 345092
rect 140872 345040 140924 345092
rect 320272 345040 320324 345092
rect 461584 345040 461636 345092
rect 118608 344972 118660 345024
rect 150440 344972 150492 345024
rect 41328 344292 41380 344344
rect 59084 344292 59136 344344
rect 150440 344292 150492 344344
rect 188344 344292 188396 344344
rect 59084 343612 59136 343664
rect 67640 343612 67692 343664
rect 117780 343544 117832 343596
rect 139584 343544 139636 343596
rect 118608 342864 118660 342916
rect 128728 342864 128780 342916
rect 139584 342864 139636 342916
rect 193864 342864 193916 342916
rect 322480 342864 322532 342916
rect 327264 342864 327316 342916
rect 352656 342864 352708 342916
rect 64604 342252 64656 342304
rect 67640 342252 67692 342304
rect 323584 342252 323636 342304
rect 493876 342252 493928 342304
rect 322848 342184 322900 342236
rect 118148 341572 118200 341624
rect 131304 341572 131356 341624
rect 37004 341504 37056 341556
rect 67916 341504 67968 341556
rect 118516 341504 118568 341556
rect 138204 341504 138256 341556
rect 63408 340892 63460 340944
rect 66168 340892 66220 340944
rect 67640 340892 67692 340944
rect 138204 340892 138256 340944
rect 190460 340892 190512 340944
rect 117320 340824 117372 340876
rect 135904 340824 135956 340876
rect 117412 340756 117464 340808
rect 130016 340756 130068 340808
rect 69296 340688 69348 340740
rect 69756 340688 69808 340740
rect 58624 340212 58676 340264
rect 70400 340212 70452 340264
rect 43812 340144 43864 340196
rect 427820 340144 427872 340196
rect 497464 340144 497516 340196
rect 75828 339872 75880 339924
rect 61844 339532 61896 339584
rect 64604 339532 64656 339584
rect 67640 339532 67692 339584
rect 111064 339532 111116 339584
rect 115664 339532 115716 339584
rect 54852 339464 54904 339516
rect 78404 339464 78456 339516
rect 107476 339464 107528 339516
rect 117412 339464 117464 339516
rect 170496 339464 170548 339516
rect 197360 339464 197412 339516
rect 46664 339396 46716 339448
rect 52184 339396 52236 339448
rect 82268 339396 82320 339448
rect 87420 339396 87472 339448
rect 87696 339396 87748 339448
rect 124864 339396 124916 339448
rect 60372 339328 60424 339380
rect 92572 339328 92624 339380
rect 93124 339328 93176 339380
rect 94596 339328 94648 339380
rect 95148 339328 95200 339380
rect 128452 339328 128504 339380
rect 194048 339396 194100 339448
rect 46204 339260 46256 339312
rect 73896 339260 73948 339312
rect 113180 339260 113232 339312
rect 113732 339260 113784 339312
rect 138020 339260 138072 339312
rect 52092 339192 52144 339244
rect 76472 339192 76524 339244
rect 105452 339192 105504 339244
rect 106188 339192 106240 339244
rect 117504 339192 117556 339244
rect 68836 338784 68888 338836
rect 98644 338784 98696 338836
rect 66996 338716 67048 338768
rect 77484 338716 77536 338768
rect 91744 338716 91796 338768
rect 121644 338716 121696 338768
rect 323032 338376 323084 338428
rect 323584 338376 323636 338428
rect 79692 338240 79744 338292
rect 83648 338240 83700 338292
rect 76472 338172 76524 338224
rect 83464 338172 83516 338224
rect 49424 337968 49476 338020
rect 83556 337968 83608 338020
rect 87604 338104 87656 338156
rect 113824 338036 113876 338088
rect 118056 338036 118108 338088
rect 112536 337968 112588 338020
rect 135352 337968 135404 338020
rect 135628 337968 135680 338020
rect 45192 337900 45244 337952
rect 74540 337900 74592 337952
rect 75276 337900 75328 337952
rect 42064 337832 42116 337884
rect 70492 337832 70544 337884
rect 57888 337764 57940 337816
rect 84200 337764 84252 337816
rect 99656 337764 99708 337816
rect 100668 337764 100720 337816
rect 119436 337900 119488 337952
rect 104808 337832 104860 337884
rect 132684 337832 132736 337884
rect 199476 338036 199528 338088
rect 136640 337968 136692 338020
rect 136824 337968 136876 338020
rect 196716 337968 196768 338020
rect 50712 337696 50764 337748
rect 86132 337696 86184 337748
rect 86868 337696 86920 337748
rect 91284 337696 91336 337748
rect 103612 337696 103664 337748
rect 109960 337696 110012 337748
rect 111800 337696 111852 337748
rect 75828 337492 75880 337544
rect 104164 337492 104216 337544
rect 107384 337492 107436 337544
rect 110236 337492 110288 337544
rect 78404 337424 78456 337476
rect 98736 337424 98788 337476
rect 103520 337424 103572 337476
rect 133880 337424 133932 337476
rect 136640 337424 136692 337476
rect 91008 337356 91060 337408
rect 91928 337356 91980 337408
rect 82820 337288 82872 337340
rect 84844 337288 84896 337340
rect 86868 337288 86920 337340
rect 131212 337356 131264 337408
rect 134524 337356 134576 337408
rect 135628 337356 135680 337408
rect 185676 337356 185728 337408
rect 103060 337220 103112 337272
rect 104808 337220 104860 337272
rect 70032 337084 70084 337136
rect 76564 337084 76616 337136
rect 111616 336744 111668 336796
rect 113824 336744 113876 336796
rect 195060 336744 195112 336796
rect 197360 336744 197412 336796
rect 46848 336676 46900 336728
rect 80796 336676 80848 336728
rect 100944 336676 100996 336728
rect 101956 336676 102008 336728
rect 56416 336608 56468 336660
rect 88984 336608 89036 336660
rect 110604 336676 110656 336728
rect 111708 336676 111760 336728
rect 111800 336676 111852 336728
rect 133972 336676 134024 336728
rect 322480 336676 322532 336728
rect 327172 336676 327224 336728
rect 328368 336676 328420 336728
rect 127256 336608 127308 336660
rect 52184 336540 52236 336592
rect 54760 336540 54812 336592
rect 82820 336540 82872 336592
rect 100300 336540 100352 336592
rect 125784 336540 125836 336592
rect 126888 336540 126940 336592
rect 70400 336472 70452 336524
rect 90364 336472 90416 336524
rect 97908 336472 97960 336524
rect 117964 336472 118016 336524
rect 50804 336404 50856 336456
rect 71964 336404 72016 336456
rect 72424 336404 72476 336456
rect 111708 336404 111760 336456
rect 124404 336404 124456 336456
rect 47584 336336 47636 336388
rect 71320 336336 71372 336388
rect 106096 336336 106148 336388
rect 111800 336336 111852 336388
rect 59084 335996 59136 336048
rect 77392 335996 77444 336048
rect 86224 335996 86276 336048
rect 121552 335996 121604 336048
rect 126888 335996 126940 336048
rect 136732 335996 136784 336048
rect 328368 335996 328420 336048
rect 388444 335996 388496 336048
rect 173164 335316 173216 335368
rect 197360 335316 197412 335368
rect 53564 335248 53616 335300
rect 87696 335248 87748 335300
rect 115112 335248 115164 335300
rect 141148 335248 141200 335300
rect 53472 335180 53524 335232
rect 86316 335180 86368 335232
rect 140688 335180 140740 335232
rect 195060 335180 195112 335232
rect 41236 335112 41288 335164
rect 71780 335112 71832 335164
rect 73068 335112 73120 335164
rect 86316 334772 86368 334824
rect 86776 334772 86828 334824
rect 98368 334704 98420 334756
rect 126428 334704 126480 334756
rect 131488 334704 131540 334756
rect 140136 334704 140188 334756
rect 140688 334704 140740 334756
rect 69664 334636 69716 334688
rect 109040 334636 109092 334688
rect 54852 334568 54904 334620
rect 103060 334568 103112 334620
rect 129740 334568 129792 334620
rect 140872 334568 140924 334620
rect 321744 334568 321796 334620
rect 328460 334568 328512 334620
rect 48044 333956 48096 334008
rect 53564 333956 53616 334008
rect 115112 333956 115164 334008
rect 115388 333956 115440 334008
rect 52000 333888 52052 333940
rect 89076 333888 89128 333940
rect 108028 333888 108080 333940
rect 131396 333888 131448 333940
rect 45468 333820 45520 333872
rect 76656 333820 76708 333872
rect 60464 333752 60516 333804
rect 81624 333752 81676 333804
rect 76656 333412 76708 333464
rect 77116 333412 77168 333464
rect 107568 333276 107620 333328
rect 115940 333276 115992 333328
rect 109040 333208 109092 333260
rect 136640 333208 136692 333260
rect 166264 333208 166316 333260
rect 352656 333208 352708 333260
rect 465080 333208 465132 333260
rect 81624 332664 81676 332716
rect 82084 332664 82136 332716
rect 73804 332596 73856 332648
rect 198832 332596 198884 332648
rect 199016 332596 199068 332648
rect 46756 332528 46808 332580
rect 79416 332528 79468 332580
rect 94504 332528 94556 332580
rect 124220 332528 124272 332580
rect 126980 332528 127032 332580
rect 188528 332528 188580 332580
rect 198096 332528 198148 332580
rect 97816 332460 97868 332512
rect 118148 332460 118200 332512
rect 97080 331916 97132 331968
rect 97816 331916 97868 331968
rect 37096 331848 37148 331900
rect 108028 331848 108080 331900
rect 322204 331712 322256 331764
rect 325700 331712 325752 331764
rect 7564 331236 7616 331288
rect 37096 331236 37148 331288
rect 122196 331236 122248 331288
rect 122656 331236 122708 331288
rect 165528 331236 165580 331288
rect 197360 331236 197412 331288
rect 93216 331168 93268 331220
rect 120816 331168 120868 331220
rect 124220 331168 124272 331220
rect 104900 330760 104952 330812
rect 128636 330760 128688 330812
rect 69112 330692 69164 330744
rect 115204 330692 115256 330744
rect 129740 330692 129792 330744
rect 169208 330692 169260 330744
rect 111800 330624 111852 330676
rect 182916 330624 182968 330676
rect 66168 330556 66220 330608
rect 151084 330556 151136 330608
rect 60556 330488 60608 330540
rect 191104 330488 191156 330540
rect 322204 330488 322256 330540
rect 325792 330488 325844 330540
rect 328552 330488 328604 330540
rect 56508 329740 56560 329792
rect 129740 329808 129792 329860
rect 123668 329740 123720 329792
rect 124312 329740 124364 329792
rect 55128 329128 55180 329180
rect 94596 329128 94648 329180
rect 85580 329060 85632 329112
rect 199384 329060 199436 329112
rect 124312 328448 124364 328500
rect 169668 328448 169720 328500
rect 197360 328448 197412 328500
rect 107752 327904 107804 327956
rect 162216 327904 162268 327956
rect 171968 327904 172020 327956
rect 198280 327904 198332 327956
rect 66904 327836 66956 327888
rect 122104 327836 122156 327888
rect 57796 327768 57848 327820
rect 111064 327768 111116 327820
rect 112444 327768 112496 327820
rect 171784 327768 171836 327820
rect 103612 327700 103664 327752
rect 169116 327700 169168 327752
rect 322848 327700 322900 327752
rect 324412 327700 324464 327752
rect 482284 327700 482336 327752
rect 195520 327088 195572 327140
rect 197360 327088 197412 327140
rect 56508 326476 56560 326528
rect 132500 326476 132552 326528
rect 88340 326408 88392 326460
rect 171876 326408 171928 326460
rect 70400 326340 70452 326392
rect 195428 326340 195480 326392
rect 110328 325660 110380 325712
rect 115296 325660 115348 325712
rect 170588 325660 170640 325712
rect 173164 325660 173216 325712
rect 104716 324980 104768 325032
rect 128544 324980 128596 325032
rect 52092 324912 52144 324964
rect 122196 324912 122248 324964
rect 162216 324912 162268 324964
rect 322756 324912 322808 324964
rect 323216 324912 323268 324964
rect 329840 324912 329892 324964
rect 334624 324912 334676 324964
rect 375932 324912 375984 324964
rect 375932 324300 375984 324352
rect 376668 324300 376720 324352
rect 580172 324300 580224 324352
rect 79324 323688 79376 323740
rect 104716 323688 104768 323740
rect 75276 323620 75328 323672
rect 114560 323620 114612 323672
rect 160836 323620 160888 323672
rect 80704 323552 80756 323604
rect 189816 323552 189868 323604
rect 322480 322940 322532 322992
rect 329840 322940 329892 322992
rect 126888 322872 126940 322924
rect 134064 322872 134116 322924
rect 197360 322872 197412 322924
rect 75276 322396 75328 322448
rect 124312 322396 124364 322448
rect 50804 322328 50856 322380
rect 107476 322328 107528 322380
rect 54944 322260 54996 322312
rect 131120 322260 131172 322312
rect 95332 322192 95384 322244
rect 174636 322192 174688 322244
rect 131120 321580 131172 321632
rect 170496 321580 170548 321632
rect 80796 320832 80848 320884
rect 191104 320832 191156 320884
rect 172428 320152 172480 320204
rect 197360 320152 197412 320204
rect 71320 319472 71372 319524
rect 135904 319472 135956 319524
rect 177948 319472 178000 319524
rect 198188 319472 198240 319524
rect 101404 319404 101456 319456
rect 181536 319404 181588 319456
rect 66168 318792 66220 318844
rect 177948 318792 178000 318844
rect 322848 318792 322900 318844
rect 323676 318792 323728 318844
rect 93216 318180 93268 318232
rect 115388 318180 115440 318232
rect 84292 318112 84344 318164
rect 113824 318112 113876 318164
rect 111248 318044 111300 318096
rect 173164 318044 173216 318096
rect 115296 317432 115348 317484
rect 197176 317432 197228 317484
rect 198648 317432 198700 317484
rect 102876 317364 102928 317416
rect 129924 317364 129976 317416
rect 322480 317364 322532 317416
rect 335544 317364 335596 317416
rect 336648 317364 336700 317416
rect 93952 316820 94004 316872
rect 116676 316820 116728 316872
rect 75184 316752 75236 316804
rect 142988 316752 143040 316804
rect 42616 316684 42668 316736
rect 122840 316684 122892 316736
rect 130384 316684 130436 316736
rect 167736 316684 167788 316736
rect 336648 316684 336700 316736
rect 454684 316684 454736 316736
rect 130292 316004 130344 316056
rect 181536 316004 181588 316056
rect 99288 315324 99340 315376
rect 142436 315324 142488 315376
rect 75920 315256 75972 315308
rect 133144 315256 133196 315308
rect 111064 314644 111116 314696
rect 175188 314644 175240 314696
rect 197360 314644 197412 314696
rect 91008 314576 91060 314628
rect 124312 314576 124364 314628
rect 125508 314576 125560 314628
rect 322480 314576 322532 314628
rect 333980 314576 334032 314628
rect 76564 313964 76616 314016
rect 176016 313964 176068 314016
rect 3424 313896 3476 313948
rect 116676 313896 116728 313948
rect 333980 313896 334032 313948
rect 500960 313896 501012 313948
rect 125508 313352 125560 313404
rect 133972 313352 134024 313404
rect 83556 313284 83608 313336
rect 108672 313284 108724 313336
rect 129188 313284 129240 313336
rect 197360 313284 197412 313336
rect 142160 313216 142212 313268
rect 143448 313216 143500 313268
rect 86316 312604 86368 312656
rect 116584 312604 116636 312656
rect 143448 312604 143500 312656
rect 195428 312604 195480 312656
rect 72424 312536 72476 312588
rect 149704 312536 149756 312588
rect 504364 312536 504416 312588
rect 580264 312536 580316 312588
rect 322848 311992 322900 312044
rect 324412 311992 324464 312044
rect 73896 311176 73948 311228
rect 120080 311176 120132 311228
rect 45376 311108 45428 311160
rect 176108 311108 176160 311160
rect 324412 311108 324464 311160
rect 413284 311108 413336 311160
rect 89720 310496 89772 310548
rect 190368 310496 190420 310548
rect 197360 310496 197412 310548
rect 100668 310428 100720 310480
rect 103612 310428 103664 310480
rect 120080 310428 120132 310480
rect 120816 310428 120868 310480
rect 195244 310428 195296 310480
rect 106096 309816 106148 309868
rect 113824 309816 113876 309868
rect 89076 309748 89128 309800
rect 142804 309748 142856 309800
rect 322480 309748 322532 309800
rect 327080 309748 327132 309800
rect 377404 309748 377456 309800
rect 56324 309136 56376 309188
rect 198096 309136 198148 309188
rect 195244 309068 195296 309120
rect 195520 309068 195572 309120
rect 101956 308524 102008 308576
rect 133144 308524 133196 308576
rect 106188 308456 106240 308508
rect 138664 308456 138716 308508
rect 93124 308388 93176 308440
rect 140136 308388 140188 308440
rect 68836 307776 68888 307828
rect 195244 307776 195296 307828
rect 322480 307708 322532 307760
rect 331220 307708 331272 307760
rect 104808 307096 104860 307148
rect 145656 307096 145708 307148
rect 79416 307028 79468 307080
rect 129004 307028 129056 307080
rect 331220 307028 331272 307080
rect 447784 307028 447836 307080
rect 71044 306416 71096 306468
rect 171784 306416 171836 306468
rect 182180 306348 182232 306400
rect 3424 306280 3476 306332
rect 21364 306280 21416 306332
rect 41052 306280 41104 306332
rect 48320 306280 48372 306332
rect 68744 305668 68796 305720
rect 120080 305668 120132 305720
rect 83648 305600 83700 305652
rect 148416 305600 148468 305652
rect 99380 304988 99432 305040
rect 169116 304988 169168 305040
rect 322480 304988 322532 305040
rect 327172 304988 327224 305040
rect 104164 304376 104216 304428
rect 137376 304376 137428 304428
rect 90364 304308 90416 304360
rect 129096 304308 129148 304360
rect 87604 304240 87656 304292
rect 167736 304240 167788 304292
rect 56416 303696 56468 303748
rect 117872 303696 117924 303748
rect 90272 303628 90324 303680
rect 171968 303628 172020 303680
rect 187240 303628 187292 303680
rect 197360 303628 197412 303680
rect 52368 302880 52420 302932
rect 70492 302880 70544 302932
rect 97356 302880 97408 302932
rect 196624 302880 196676 302932
rect 111156 302404 111208 302456
rect 111616 302404 111668 302456
rect 158076 302404 158128 302456
rect 87604 302336 87656 302388
rect 138756 302336 138808 302388
rect 79140 302268 79192 302320
rect 142896 302268 142948 302320
rect 67364 302200 67416 302252
rect 193128 302200 193180 302252
rect 197360 302200 197412 302252
rect 322480 302200 322532 302252
rect 327080 302200 327132 302252
rect 98552 301588 98604 301640
rect 111064 301588 111116 301640
rect 82084 301520 82136 301572
rect 147036 301520 147088 301572
rect 322204 301520 322256 301572
rect 333980 301520 334032 301572
rect 53656 301452 53708 301504
rect 132592 301452 132644 301504
rect 175096 301452 175148 301504
rect 197268 301452 197320 301504
rect 322848 301452 322900 301504
rect 325056 301452 325108 301504
rect 429200 301452 429252 301504
rect 125784 300976 125836 301028
rect 126244 300976 126296 301028
rect 152556 300976 152608 301028
rect 109684 300908 109736 300960
rect 110328 300908 110380 300960
rect 175096 300908 175148 300960
rect 84200 300840 84252 300892
rect 166264 300840 166316 300892
rect 333980 300840 334032 300892
rect 468484 300840 468536 300892
rect 117872 300772 117924 300824
rect 132776 300772 132828 300824
rect 133788 300772 133840 300824
rect 182180 300772 182232 300824
rect 183468 300772 183520 300824
rect 117964 300160 118016 300212
rect 125784 300160 125836 300212
rect 104992 300092 105044 300144
rect 127164 300092 127216 300144
rect 148508 300228 148560 300280
rect 133788 300160 133840 300212
rect 155316 300160 155368 300212
rect 138020 300092 138072 300144
rect 163596 300092 163648 300144
rect 183468 300092 183520 300144
rect 197360 300092 197412 300144
rect 335268 300092 335320 300144
rect 580356 300092 580408 300144
rect 87512 299684 87564 299736
rect 135996 299684 136048 299736
rect 102140 299616 102192 299668
rect 184296 299616 184348 299668
rect 22744 299548 22796 299600
rect 117964 299548 118016 299600
rect 69020 299480 69072 299532
rect 166448 299480 166500 299532
rect 65524 299412 65576 299464
rect 68652 299412 68704 299464
rect 83464 298732 83516 298784
rect 129924 298732 129976 298784
rect 322480 298732 322532 298784
rect 330484 298732 330536 298784
rect 113824 298392 113876 298444
rect 156696 298392 156748 298444
rect 82268 298324 82320 298376
rect 134616 298324 134668 298376
rect 68652 298256 68704 298308
rect 159640 298256 159692 298308
rect 93860 298188 93912 298240
rect 196716 298188 196768 298240
rect 69112 298120 69164 298172
rect 187240 298120 187292 298172
rect 17224 297372 17276 297424
rect 57244 297440 57296 297492
rect 97080 297440 97132 297492
rect 75000 297372 75052 297424
rect 147864 297372 147916 297424
rect 148140 297372 148192 297424
rect 330484 297372 330536 297424
rect 353392 297372 353444 297424
rect 407764 297372 407816 297424
rect 193036 297168 193088 297220
rect 197360 297168 197412 297220
rect 107292 296964 107344 297016
rect 123760 296964 123812 297016
rect 102876 296896 102928 296948
rect 145564 296896 145616 296948
rect 148140 296896 148192 296948
rect 152464 296896 152516 296948
rect 116676 296828 116728 296880
rect 159548 296828 159600 296880
rect 97080 296760 97132 296812
rect 160836 296760 160888 296812
rect 76472 296692 76524 296744
rect 182916 296692 182968 296744
rect 54760 295944 54812 295996
rect 71780 295944 71832 295996
rect 114468 295944 114520 295996
rect 115296 295944 115348 295996
rect 65984 295672 66036 295724
rect 196624 295672 196676 295724
rect 83556 295604 83608 295656
rect 133236 295604 133288 295656
rect 68928 295536 68980 295588
rect 125048 295536 125100 295588
rect 93216 295468 93268 295520
rect 188436 295468 188488 295520
rect 69204 295400 69256 295452
rect 195888 295400 195940 295452
rect 197452 295400 197504 295452
rect 117228 295332 117280 295384
rect 124864 295332 124916 295384
rect 322480 295332 322532 295384
rect 331220 295332 331272 295384
rect 80336 295264 80388 295316
rect 86224 295264 86276 295316
rect 117044 295264 117096 295316
rect 123484 295264 123536 295316
rect 111248 294924 111300 294976
rect 124956 294924 125008 294976
rect 84844 294856 84896 294908
rect 91744 294856 91796 294908
rect 94504 294856 94556 294908
rect 111156 294856 111208 294908
rect 106740 294788 106792 294840
rect 126336 294788 126388 294840
rect 82912 294720 82964 294772
rect 107292 294720 107344 294772
rect 119620 294720 119672 294772
rect 147772 294720 147824 294772
rect 71320 294652 71372 294704
rect 83464 294652 83516 294704
rect 87420 294652 87472 294704
rect 117228 294652 117280 294704
rect 117688 294652 117740 294704
rect 173256 294652 173308 294704
rect 71964 294584 72016 294636
rect 101404 294584 101456 294636
rect 113824 294584 113876 294636
rect 195336 294584 195388 294636
rect 72608 294516 72660 294568
rect 75000 294516 75052 294568
rect 104900 294312 104952 294364
rect 105820 294312 105872 294364
rect 107660 294312 107712 294364
rect 108396 294312 108448 294364
rect 109316 294312 109368 294364
rect 112444 294312 112496 294364
rect 79048 294176 79100 294228
rect 79232 294176 79284 294228
rect 49608 294108 49660 294160
rect 75184 294108 75236 294160
rect 86132 294108 86184 294160
rect 87604 294108 87656 294160
rect 41236 294040 41288 294092
rect 74540 294040 74592 294092
rect 99288 294040 99340 294092
rect 101588 294040 101640 294092
rect 33784 293972 33836 294024
rect 79048 293972 79100 294024
rect 100944 293972 100996 294024
rect 118700 293972 118752 294024
rect 3424 293836 3476 293888
rect 7564 293836 7616 293888
rect 41328 293224 41380 293276
rect 99288 293224 99340 293276
rect 111708 293224 111760 293276
rect 148324 293224 148376 293276
rect 322848 293224 322900 293276
rect 324320 293224 324372 293276
rect 370504 293224 370556 293276
rect 91928 292816 91980 292868
rect 117504 292816 117556 292868
rect 115204 292748 115256 292800
rect 115756 292748 115808 292800
rect 155408 292748 155460 292800
rect 53104 292680 53156 292732
rect 92572 292680 92624 292732
rect 92940 292680 92992 292732
rect 107384 292680 107436 292732
rect 107568 292680 107620 292732
rect 151360 292680 151412 292732
rect 68744 292612 68796 292664
rect 73804 292612 73856 292664
rect 73896 292612 73948 292664
rect 124128 292612 124180 292664
rect 153476 292612 153528 292664
rect 154672 292612 154724 292664
rect 8208 292544 8260 292596
rect 96436 292544 96488 292596
rect 98368 292544 98420 292596
rect 98736 292544 98788 292596
rect 189816 292544 189868 292596
rect 194048 292544 194100 292596
rect 197452 292544 197504 292596
rect 124128 292476 124180 292528
rect 129832 292476 129884 292528
rect 71688 292340 71740 292392
rect 75368 292340 75420 292392
rect 121460 291932 121512 291984
rect 153476 291932 153528 291984
rect 153936 291932 153988 291984
rect 61844 291796 61896 291848
rect 71044 291864 71096 291916
rect 110880 291864 110932 291916
rect 112812 291864 112864 291916
rect 117504 291864 117556 291916
rect 118700 291864 118752 291916
rect 151176 291864 151228 291916
rect 177396 291796 177448 291848
rect 123668 291252 123720 291304
rect 188528 291184 188580 291236
rect 322848 291184 322900 291236
rect 324320 291184 324372 291236
rect 499672 291184 499724 291236
rect 38108 291116 38160 291168
rect 38476 291116 38528 291168
rect 67640 291116 67692 291168
rect 148416 291116 148468 291168
rect 148600 291116 148652 291168
rect 25504 290436 25556 290488
rect 38108 290436 38160 290488
rect 325056 290436 325108 290488
rect 420920 290436 420972 290488
rect 148600 289960 148652 290012
rect 179236 289960 179288 290012
rect 121552 289892 121604 289944
rect 156604 289892 156656 289944
rect 59084 289824 59136 289876
rect 67640 289824 67692 289876
rect 121460 289824 121512 289876
rect 169208 289824 169260 289876
rect 197452 289824 197504 289876
rect 121552 289756 121604 289808
rect 187056 289756 187108 289808
rect 69020 289144 69072 289196
rect 69756 289144 69808 289196
rect 123576 289144 123628 289196
rect 126428 289144 126480 289196
rect 168288 289144 168340 289196
rect 123668 289076 123720 289128
rect 185768 289076 185820 289128
rect 60372 288396 60424 288448
rect 67640 288396 67692 288448
rect 168288 288396 168340 288448
rect 197452 288396 197504 288448
rect 322848 288396 322900 288448
rect 327264 288396 327316 288448
rect 121460 288328 121512 288380
rect 166356 288328 166408 288380
rect 121552 288260 121604 288312
rect 152004 288260 152056 288312
rect 153108 288260 153160 288312
rect 153108 287648 153160 287700
rect 165068 287648 165120 287700
rect 46756 287036 46808 287088
rect 67640 287036 67692 287088
rect 362960 287036 363012 287088
rect 364248 287036 364300 287088
rect 506480 287036 506532 287088
rect 55128 286968 55180 287020
rect 67732 286968 67784 287020
rect 121552 286968 121604 287020
rect 124220 286968 124272 287020
rect 60556 286900 60608 286952
rect 67640 286900 67692 286952
rect 322204 286288 322256 286340
rect 362960 286288 363012 286340
rect 182088 285744 182140 285796
rect 197452 285744 197504 285796
rect 57520 285676 57572 285728
rect 67824 285676 67876 285728
rect 120724 285676 120776 285728
rect 196808 285676 196860 285728
rect 57796 285608 57848 285660
rect 67640 285608 67692 285660
rect 121460 285608 121512 285660
rect 193956 285608 194008 285660
rect 121552 285540 121604 285592
rect 153200 285540 153252 285592
rect 43812 284316 43864 284368
rect 67640 284316 67692 284368
rect 121460 284248 121512 284300
rect 147128 284248 147180 284300
rect 127072 283568 127124 283620
rect 179420 283568 179472 283620
rect 123576 282956 123628 283008
rect 127072 282956 127124 283008
rect 121460 282888 121512 282940
rect 127716 282888 127768 282940
rect 179420 282888 179472 282940
rect 180708 282888 180760 282940
rect 197452 282888 197504 282940
rect 322480 282888 322532 282940
rect 329932 282888 329984 282940
rect 43996 282820 44048 282872
rect 67640 282820 67692 282872
rect 124956 282140 125008 282192
rect 150624 282140 150676 282192
rect 184756 281596 184808 281648
rect 190460 281596 190512 281648
rect 191748 281596 191800 281648
rect 121460 281528 121512 281580
rect 170404 281528 170456 281580
rect 173348 281528 173400 281580
rect 197452 281528 197504 281580
rect 121552 281460 121604 281512
rect 192484 281460 192536 281512
rect 191748 281392 191800 281444
rect 197452 281392 197504 281444
rect 45468 280168 45520 280220
rect 67640 280168 67692 280220
rect 121460 280168 121512 280220
rect 148416 280168 148468 280220
rect 322480 280168 322532 280220
rect 336004 280168 336056 280220
rect 40868 280100 40920 280152
rect 41144 280100 41196 280152
rect 67732 280100 67784 280152
rect 121552 280100 121604 280152
rect 130384 280100 130436 280152
rect 29644 279420 29696 279472
rect 40868 279420 40920 279472
rect 52276 279420 52328 279472
rect 57796 279420 57848 279472
rect 67640 279420 67692 279472
rect 123760 279420 123812 279472
rect 163688 279420 163740 279472
rect 121460 278740 121512 278792
rect 192484 278740 192536 278792
rect 121552 278672 121604 278724
rect 184848 278672 184900 278724
rect 184848 278196 184900 278248
rect 187056 278196 187108 278248
rect 195796 277448 195848 277500
rect 197452 277448 197504 277500
rect 47952 277380 48004 277432
rect 67640 277380 67692 277432
rect 121460 277312 121512 277364
rect 131120 277312 131172 277364
rect 61844 276632 61896 276684
rect 67640 276632 67692 276684
rect 322204 276088 322256 276140
rect 121460 276020 121512 276072
rect 130568 276020 130620 276072
rect 322848 276020 322900 276072
rect 325056 276020 325108 276072
rect 521660 276020 521712 276072
rect 191748 275408 191800 275460
rect 197360 275408 197412 275460
rect 121552 274796 121604 274848
rect 128268 274796 128320 274848
rect 129924 274796 129976 274848
rect 121460 274728 121512 274780
rect 131856 274728 131908 274780
rect 53656 274660 53708 274712
rect 67640 274660 67692 274712
rect 121552 274660 121604 274712
rect 122104 274660 122156 274712
rect 162400 274660 162452 274712
rect 187148 274660 187200 274712
rect 197360 274660 197412 274712
rect 52092 274592 52144 274644
rect 67732 274592 67784 274644
rect 322388 274592 322440 274644
rect 339592 274592 339644 274644
rect 339592 273912 339644 273964
rect 382924 273912 382976 273964
rect 121460 273300 121512 273352
rect 171876 273300 171928 273352
rect 52276 273232 52328 273284
rect 67640 273232 67692 273284
rect 123484 273232 123536 273284
rect 194508 273232 194560 273284
rect 197360 273232 197412 273284
rect 121460 273164 121512 273216
rect 133880 273164 133932 273216
rect 125140 271872 125192 271924
rect 187148 271872 187200 271924
rect 336004 271872 336056 271924
rect 400864 271872 400916 271924
rect 417424 271872 417476 271924
rect 419540 271872 419592 271924
rect 580172 271872 580224 271924
rect 57704 271804 57756 271856
rect 67732 271804 67784 271856
rect 127716 271124 127768 271176
rect 197360 271124 197412 271176
rect 63224 270512 63276 270564
rect 67640 270512 67692 270564
rect 121460 270512 121512 270564
rect 173256 270512 173308 270564
rect 322848 270512 322900 270564
rect 331312 270512 331364 270564
rect 56324 270444 56376 270496
rect 67732 270444 67784 270496
rect 57704 269764 57756 269816
rect 67824 269764 67876 269816
rect 66076 269084 66128 269136
rect 68192 269084 68244 269136
rect 121552 269084 121604 269136
rect 130384 269084 130436 269136
rect 322848 269084 322900 269136
rect 326344 269084 326396 269136
rect 52460 269016 52512 269068
rect 53564 269016 53616 269068
rect 67640 269016 67692 269068
rect 121460 269016 121512 269068
rect 149152 269016 149204 269068
rect 149336 269016 149388 269068
rect 45284 268404 45336 268456
rect 52092 268404 52144 268456
rect 149336 268404 149388 268456
rect 181628 268404 181680 268456
rect 21364 268336 21416 268388
rect 52460 268336 52512 268388
rect 125048 268336 125100 268388
rect 183376 268336 183428 268388
rect 183376 267792 183428 267844
rect 197360 267792 197412 267844
rect 121460 267724 121512 267776
rect 191196 267724 191248 267776
rect 48136 267656 48188 267708
rect 67732 267656 67784 267708
rect 322480 267656 322532 267708
rect 342260 267656 342312 267708
rect 52092 266976 52144 267028
rect 67640 266976 67692 267028
rect 160836 266976 160888 267028
rect 176660 266976 176712 267028
rect 342260 266976 342312 267028
rect 499856 266976 499908 267028
rect 121460 266432 121512 266484
rect 147220 266432 147272 266484
rect 3056 266364 3108 266416
rect 54484 266364 54536 266416
rect 121552 266364 121604 266416
rect 149796 266364 149848 266416
rect 176660 266364 176712 266416
rect 177856 266364 177908 266416
rect 197360 266364 197412 266416
rect 54852 266296 54904 266348
rect 67732 266296 67784 266348
rect 121460 265004 121512 265056
rect 152648 265004 152700 265056
rect 54944 264936 54996 264988
rect 67640 264936 67692 264988
rect 68560 264936 68612 264988
rect 68836 264936 68888 264988
rect 121552 264936 121604 264988
rect 158168 264936 158220 264988
rect 322480 264936 322532 264988
rect 330024 264936 330076 264988
rect 14464 264188 14516 264240
rect 43904 264188 43956 264240
rect 55864 264188 55916 264240
rect 124128 264188 124180 264240
rect 195704 264188 195756 264240
rect 197360 264188 197412 264240
rect 56232 263644 56284 263696
rect 67640 263644 67692 263696
rect 55864 263576 55916 263628
rect 56324 263576 56376 263628
rect 67732 263576 67784 263628
rect 121552 263576 121604 263628
rect 134708 263576 134760 263628
rect 335268 263576 335320 263628
rect 490564 263576 490616 263628
rect 56508 263508 56560 263560
rect 67640 263508 67692 263560
rect 121460 263508 121512 263560
rect 136732 263508 136784 263560
rect 137100 263508 137152 263560
rect 332600 263508 332652 263560
rect 68560 262896 68612 262948
rect 68928 262896 68980 262948
rect 137100 262828 137152 262880
rect 178776 262828 178828 262880
rect 121460 262760 121512 262812
rect 125140 262760 125192 262812
rect 56508 262216 56560 262268
rect 67640 262216 67692 262268
rect 322480 262216 322532 262268
rect 332600 262216 332652 262268
rect 65984 262148 66036 262200
rect 67732 262148 67784 262200
rect 121552 262148 121604 262200
rect 126888 262148 126940 262200
rect 121460 261876 121512 261928
rect 123484 261876 123536 261928
rect 126888 261468 126940 261520
rect 160928 261468 160980 261520
rect 140044 260856 140096 260908
rect 190276 260856 190328 260908
rect 197360 260856 197412 260908
rect 56416 260788 56468 260840
rect 67640 260788 67692 260840
rect 121460 260788 121512 260840
rect 139584 260788 139636 260840
rect 140688 260788 140740 260840
rect 370504 260108 370556 260160
rect 548524 260108 548576 260160
rect 139584 259496 139636 259548
rect 144184 259496 144236 259548
rect 121460 259428 121512 259480
rect 170680 259428 170732 259480
rect 179880 259428 179932 259480
rect 197360 259428 197412 259480
rect 322572 259428 322624 259480
rect 327356 259428 327408 259480
rect 121552 259360 121604 259412
rect 143632 259360 143684 259412
rect 144828 259360 144880 259412
rect 144828 258680 144880 258732
rect 166540 258680 166592 258732
rect 548524 258680 548576 258732
rect 579988 258680 580040 258732
rect 61844 258068 61896 258120
rect 67732 258068 67784 258120
rect 121644 258068 121696 258120
rect 154120 258068 154172 258120
rect 324412 258068 324464 258120
rect 425060 258068 425112 258120
rect 34428 258000 34480 258052
rect 67640 258000 67692 258052
rect 121460 258000 121512 258052
rect 154580 258000 154632 258052
rect 15844 257320 15896 257372
rect 34428 257320 34480 257372
rect 131764 257320 131816 257372
rect 197360 257320 197412 257372
rect 65984 256708 66036 256760
rect 68008 256708 68060 256760
rect 121552 256708 121604 256760
rect 134524 256708 134576 256760
rect 121460 256640 121512 256692
rect 148600 256640 148652 256692
rect 121552 256572 121604 256624
rect 133880 256572 133932 256624
rect 135168 256572 135220 256624
rect 135168 255960 135220 256012
rect 166356 255960 166408 256012
rect 178776 255348 178828 255400
rect 180616 255348 180668 255400
rect 53564 255280 53616 255332
rect 67640 255280 67692 255332
rect 176108 255280 176160 255332
rect 179880 255280 179932 255332
rect 197360 255280 197412 255332
rect 50988 255212 51040 255264
rect 67732 255212 67784 255264
rect 143448 255212 143500 255264
rect 194048 255212 194100 255264
rect 52184 255144 52236 255196
rect 67640 255144 67692 255196
rect 142988 254804 143040 254856
rect 143448 254804 143500 254856
rect 121460 253920 121512 253972
rect 161020 253920 161072 253972
rect 48320 253852 48372 253904
rect 48964 253852 49016 253904
rect 67640 253852 67692 253904
rect 32404 253172 32456 253224
rect 48964 253172 49016 253224
rect 121460 252628 121512 252680
rect 126336 252628 126388 252680
rect 121552 252560 121604 252612
rect 155500 252560 155552 252612
rect 191288 252560 191340 252612
rect 197360 252560 197412 252612
rect 121460 252492 121512 252544
rect 155960 252492 156012 252544
rect 322480 251268 322532 251320
rect 325792 251268 325844 251320
rect 61752 251200 61804 251252
rect 67640 251200 67692 251252
rect 121460 251200 121512 251252
rect 188620 251200 188672 251252
rect 66168 251132 66220 251184
rect 67732 251132 67784 251184
rect 120632 251132 120684 251184
rect 140964 251132 141016 251184
rect 121460 249772 121512 249824
rect 137468 249772 137520 249824
rect 121552 249704 121604 249756
rect 129188 249704 129240 249756
rect 39856 249024 39908 249076
rect 57612 249024 57664 249076
rect 189816 249024 189868 249076
rect 194416 249024 194468 249076
rect 194416 248752 194468 248804
rect 197360 248752 197412 248804
rect 57612 248480 57664 248532
rect 67640 248480 67692 248532
rect 120080 248412 120132 248464
rect 176200 248412 176252 248464
rect 320272 248412 320324 248464
rect 434720 248412 434772 248464
rect 121552 248344 121604 248396
rect 146300 248344 146352 248396
rect 121460 247936 121512 247988
rect 123484 247936 123536 247988
rect 134616 247868 134668 247920
rect 147128 247868 147180 247920
rect 146300 247800 146352 247852
rect 173440 247800 173492 247852
rect 122288 247732 122340 247784
rect 160836 247732 160888 247784
rect 122196 247664 122248 247716
rect 164976 247664 165028 247716
rect 65892 247120 65944 247172
rect 67732 247120 67784 247172
rect 60464 247052 60516 247104
rect 67640 247052 67692 247104
rect 120080 246304 120132 246356
rect 135260 246304 135312 246356
rect 192944 246304 192996 246356
rect 197360 246304 197412 246356
rect 121552 245760 121604 245812
rect 123760 245760 123812 245812
rect 64788 245692 64840 245744
rect 67640 245692 67692 245744
rect 56416 245624 56468 245676
rect 67732 245624 67784 245676
rect 121460 245624 121512 245676
rect 151268 245624 151320 245676
rect 320364 245624 320416 245676
rect 374644 245624 374696 245676
rect 50804 245556 50856 245608
rect 67640 245556 67692 245608
rect 121552 245556 121604 245608
rect 138204 245556 138256 245608
rect 46664 245488 46716 245540
rect 55864 245488 55916 245540
rect 56416 245488 56468 245540
rect 121460 244264 121512 244316
rect 154028 244264 154080 244316
rect 322848 244264 322900 244316
rect 324412 244264 324464 244316
rect 378784 244264 378836 244316
rect 37096 244196 37148 244248
rect 67732 244196 67784 244248
rect 45376 244128 45428 244180
rect 67640 244128 67692 244180
rect 68468 243516 68520 243568
rect 68928 243516 68980 243568
rect 137284 242972 137336 243024
rect 184388 242972 184440 243024
rect 121460 242904 121512 242956
rect 185860 242904 185912 242956
rect 321744 242904 321796 242956
rect 449164 242904 449216 242956
rect 121552 242836 121604 242888
rect 137284 242836 137336 242888
rect 121460 242768 121512 242820
rect 132592 242768 132644 242820
rect 133788 242768 133840 242820
rect 196808 242496 196860 242548
rect 197268 242496 197320 242548
rect 198464 242496 198516 242548
rect 154120 242156 154172 242208
rect 189816 242156 189868 242208
rect 3424 241408 3476 241460
rect 34612 241408 34664 241460
rect 34612 240728 34664 240780
rect 35532 240728 35584 240780
rect 58900 240728 58952 240780
rect 158168 240728 158220 240780
rect 194324 240728 194376 240780
rect 536840 240728 536892 240780
rect 580264 240728 580316 240780
rect 121460 240184 121512 240236
rect 126428 240184 126480 240236
rect 325056 240184 325108 240236
rect 502432 240184 502484 240236
rect 119988 240116 120040 240168
rect 199660 240116 199712 240168
rect 320088 240116 320140 240168
rect 536840 240116 536892 240168
rect 3516 240048 3568 240100
rect 39948 240048 40000 240100
rect 55036 240048 55088 240100
rect 68652 240048 68704 240100
rect 120816 240048 120868 240100
rect 329840 240048 329892 240100
rect 130568 239980 130620 240032
rect 327080 239980 327132 240032
rect 71780 239912 71832 239964
rect 201408 239912 201460 239964
rect 320272 239912 320324 239964
rect 70400 239776 70452 239828
rect 71308 239776 71360 239828
rect 75920 239776 75972 239828
rect 77104 239776 77156 239828
rect 77300 239776 77352 239828
rect 78392 239776 78444 239828
rect 84292 239776 84344 239828
rect 85476 239776 85528 239828
rect 86960 239776 87012 239828
rect 88052 239776 88104 239828
rect 92480 239776 92532 239828
rect 93204 239776 93256 239828
rect 95240 239776 95292 239828
rect 96424 239776 96476 239828
rect 99380 239776 99432 239828
rect 100288 239776 100340 239828
rect 100760 239776 100812 239828
rect 101576 239776 101628 239828
rect 102140 239776 102192 239828
rect 102864 239776 102916 239828
rect 110420 239776 110472 239828
rect 111236 239776 111288 239828
rect 114560 239776 114612 239828
rect 115744 239776 115796 239828
rect 238760 239776 238812 239828
rect 239910 239776 239962 239828
rect 247040 239776 247092 239828
rect 248282 239776 248334 239828
rect 258080 239776 258132 239828
rect 259230 239776 259282 239828
rect 266360 239776 266412 239828
rect 267602 239776 267654 239828
rect 285680 239776 285732 239828
rect 286922 239776 286974 239828
rect 195888 239640 195940 239692
rect 200856 239640 200908 239692
rect 193036 239504 193088 239556
rect 201592 239504 201644 239556
rect 69848 239436 69900 239488
rect 76564 239436 76616 239488
rect 187240 239436 187292 239488
rect 196808 239436 196860 239488
rect 65984 239368 66036 239420
rect 82084 239368 82136 239420
rect 153936 239368 153988 239420
rect 195152 239368 195204 239420
rect 512092 239368 512144 239420
rect 580172 239368 580224 239420
rect 117044 238960 117096 239012
rect 125600 238960 125652 239012
rect 85672 238892 85724 238944
rect 86776 238892 86828 238944
rect 123668 238892 123720 238944
rect 82912 238824 82964 238876
rect 120080 238824 120132 238876
rect 121460 238824 121512 238876
rect 304264 238824 304316 238876
rect 39948 238756 40000 238808
rect 111892 238756 111944 238808
rect 112536 238756 112588 238808
rect 114468 238756 114520 238808
rect 131212 238756 131264 238808
rect 252836 238756 252888 238808
rect 512092 238756 512144 238808
rect 53748 238688 53800 238740
rect 82268 238688 82320 238740
rect 83556 238688 83608 238740
rect 149060 238688 149112 238740
rect 316592 238688 316644 238740
rect 48044 238620 48096 238672
rect 72608 238620 72660 238672
rect 88708 238620 88760 238672
rect 241888 238620 241940 238672
rect 299204 238620 299256 238672
rect 320088 238620 320140 238672
rect 118332 238552 118384 238604
rect 143540 238552 143592 238604
rect 304264 238552 304316 238604
rect 312084 238552 312136 238604
rect 115112 238484 115164 238536
rect 144920 238484 144972 238536
rect 69940 238416 69992 238468
rect 119988 238416 120040 238468
rect 71964 238144 72016 238196
rect 78864 238144 78916 238196
rect 194324 238144 194376 238196
rect 204168 238144 204220 238196
rect 60372 238076 60424 238128
rect 72424 238076 72476 238128
rect 73252 238076 73304 238128
rect 83464 238076 83516 238128
rect 159640 238076 159692 238128
rect 201408 238076 201460 238128
rect 314108 238076 314160 238128
rect 320364 238076 320416 238128
rect 64788 238008 64840 238060
rect 88984 238008 89036 238060
rect 155500 238008 155552 238060
rect 204996 238008 205048 238060
rect 316592 238008 316644 238060
rect 438860 238008 438912 238060
rect 323676 237464 323728 237516
rect 332968 237464 333020 237516
rect 80980 237396 81032 237448
rect 86224 237396 86276 237448
rect 199936 237396 199988 237448
rect 202328 237396 202380 237448
rect 218704 237396 218756 237448
rect 220636 237396 220688 237448
rect 228548 237396 228600 237448
rect 229652 237396 229704 237448
rect 235264 237396 235316 237448
rect 236092 237396 236144 237448
rect 244924 237396 244976 237448
rect 246396 237396 246448 237448
rect 251640 237396 251692 237448
rect 254768 237396 254820 237448
rect 283564 237396 283616 237448
rect 284392 237396 284444 237448
rect 312084 237396 312136 237448
rect 312544 237396 312596 237448
rect 318064 237396 318116 237448
rect 318524 237396 318576 237448
rect 498292 237396 498344 237448
rect 57888 237328 57940 237380
rect 86132 237328 86184 237380
rect 128268 237328 128320 237380
rect 322204 237328 322256 237380
rect 107384 237260 107436 237312
rect 132500 237260 132552 237312
rect 162400 237260 162452 237312
rect 332600 237260 332652 237312
rect 95792 237192 95844 237244
rect 128360 237192 128412 237244
rect 166540 237192 166592 237244
rect 319352 237192 319404 237244
rect 201408 237124 201460 237176
rect 303712 237124 303764 237176
rect 181628 237056 181680 237108
rect 276020 237056 276072 237108
rect 195152 236988 195204 237040
rect 210424 236988 210476 237040
rect 276020 235968 276072 236020
rect 276664 235968 276716 236020
rect 303712 235968 303764 236020
rect 304264 235968 304316 236020
rect 326988 235968 327040 236020
rect 349160 235968 349212 236020
rect 48228 235900 48280 235952
rect 98368 235900 98420 235952
rect 106096 235900 106148 235952
rect 173348 235900 173400 235952
rect 195704 235900 195756 235952
rect 504364 235900 504416 235952
rect 54484 235832 54536 235884
rect 85672 235832 85724 235884
rect 89352 235832 89404 235884
rect 142252 235832 142304 235884
rect 149796 235832 149848 235884
rect 321560 235832 321612 235884
rect 97724 235764 97776 235816
rect 251640 235764 251692 235816
rect 58900 235696 58952 235748
rect 103520 235696 103572 235748
rect 113824 235696 113876 235748
rect 131764 235696 131816 235748
rect 165068 235696 165120 235748
rect 301504 235696 301556 235748
rect 91284 235628 91336 235680
rect 124956 235628 125008 235680
rect 191196 235628 191248 235680
rect 326344 235628 326396 235680
rect 326988 235628 327040 235680
rect 118608 235560 118660 235612
rect 129740 235560 129792 235612
rect 185768 235220 185820 235272
rect 268384 235220 268436 235272
rect 503720 234948 503772 235000
rect 504364 234948 504416 235000
rect 117688 234676 117740 234728
rect 118608 234676 118660 234728
rect 321560 234676 321612 234728
rect 322204 234676 322256 234728
rect 288900 234608 288952 234660
rect 289452 234608 289504 234660
rect 432604 234608 432656 234660
rect 61752 234540 61804 234592
rect 256700 234540 256752 234592
rect 50896 234472 50948 234524
rect 91744 234472 91796 234524
rect 95148 234472 95200 234524
rect 170588 234472 170640 234524
rect 81624 234404 81676 234456
rect 123576 234404 123628 234456
rect 151360 234404 151412 234456
rect 211804 234404 211856 234456
rect 212264 234404 212316 234456
rect 106740 234336 106792 234388
rect 140044 234336 140096 234388
rect 256700 234132 256752 234184
rect 257344 234132 257396 234184
rect 196716 233996 196768 234048
rect 224224 233996 224276 234048
rect 84200 233928 84252 233980
rect 74540 233860 74592 233912
rect 75184 233860 75236 233912
rect 171968 233928 172020 233980
rect 228364 233928 228416 233980
rect 118700 233860 118752 233912
rect 119712 233860 119764 233912
rect 188620 233860 188672 233912
rect 318708 233928 318760 233980
rect 321652 233928 321704 233980
rect 316684 233860 316736 233912
rect 319260 233860 319312 233912
rect 84292 233724 84344 233776
rect 205640 233248 205692 233300
rect 205824 233248 205876 233300
rect 307024 233248 307076 233300
rect 56324 233180 56376 233232
rect 324412 233180 324464 233232
rect 161020 233112 161072 233164
rect 325884 233112 325936 233164
rect 333980 233112 334032 233164
rect 53564 233044 53616 233096
rect 176108 233044 176160 233096
rect 189816 233044 189868 233096
rect 331312 233044 331364 233096
rect 155408 232976 155460 233028
rect 218796 232976 218848 233028
rect 183376 232568 183428 232620
rect 206468 232568 206520 232620
rect 67364 232500 67416 232552
rect 106924 232500 106976 232552
rect 198832 232500 198884 232552
rect 324412 232500 324464 232552
rect 418804 231820 418856 231872
rect 580172 231820 580224 231872
rect 99472 231752 99524 231804
rect 269120 231752 269172 231804
rect 269764 231752 269816 231804
rect 54944 231684 54996 231736
rect 205640 231684 205692 231736
rect 109868 231616 109920 231668
rect 136640 231616 136692 231668
rect 204168 231616 204220 231668
rect 329932 231616 329984 231668
rect 152464 231548 152516 231600
rect 277400 231548 277452 231600
rect 278044 231548 278096 231600
rect 182916 231480 182968 231532
rect 244924 231480 244976 231532
rect 69204 231140 69256 231192
rect 104164 231140 104216 231192
rect 103612 231072 103664 231124
rect 190184 231072 190236 231124
rect 191288 231072 191340 231124
rect 192484 231072 192536 231124
rect 226984 231072 227036 231124
rect 76012 230392 76064 230444
rect 126980 230392 127032 230444
rect 280160 230392 280212 230444
rect 281448 230392 281500 230444
rect 78864 230324 78916 230376
rect 202880 230324 202932 230376
rect 203524 230324 203576 230376
rect 211620 230324 211672 230376
rect 327172 230324 327224 230376
rect 328368 230324 328420 230376
rect 188528 229916 188580 229968
rect 213368 229916 213420 229968
rect 61844 229848 61896 229900
rect 119344 229848 119396 229900
rect 196624 229848 196676 229900
rect 233884 229848 233936 229900
rect 111892 229780 111944 229832
rect 262864 229780 262916 229832
rect 328368 229780 328420 229832
rect 340972 229780 341024 229832
rect 4804 229712 4856 229764
rect 83556 229712 83608 229764
rect 90548 229712 90600 229764
rect 255596 229712 255648 229764
rect 281448 229712 281500 229764
rect 334716 229712 334768 229764
rect 43812 229032 43864 229084
rect 327356 229032 327408 229084
rect 118792 228964 118844 229016
rect 143448 228964 143500 229016
rect 173440 228964 173492 229016
rect 324320 228964 324372 229016
rect 77392 228896 77444 228948
rect 216680 228896 216732 228948
rect 185860 228828 185912 228880
rect 321652 228828 321704 228880
rect 162216 228760 162268 228812
rect 262220 228760 262272 228812
rect 59084 228420 59136 228472
rect 166356 228420 166408 228472
rect 327356 228420 327408 228472
rect 343732 228420 343784 228472
rect 143448 228352 143500 228404
rect 495624 228352 495676 228404
rect 216680 227740 216732 227792
rect 217324 227740 217376 227792
rect 262220 227740 262272 227792
rect 262956 227740 263008 227792
rect 110512 227672 110564 227724
rect 140780 227672 140832 227724
rect 170496 227672 170548 227724
rect 418804 227672 418856 227724
rect 336004 227604 336056 227656
rect 87052 227536 87104 227588
rect 235264 227536 235316 227588
rect 204996 227468 205048 227520
rect 330024 227468 330076 227520
rect 190184 227060 190236 227112
rect 202236 227060 202288 227112
rect 96620 226992 96672 227044
rect 252836 226992 252888 227044
rect 305644 226992 305696 227044
rect 340236 226992 340288 227044
rect 110512 226312 110564 226364
rect 111064 226312 111116 226364
rect 80060 226244 80112 226296
rect 222200 226244 222252 226296
rect 155316 226176 155368 226228
rect 289820 226176 289872 226228
rect 74632 226108 74684 226160
rect 201592 226108 201644 226160
rect 202788 226108 202840 226160
rect 194416 225768 194468 225820
rect 213276 225768 213328 225820
rect 196808 225700 196860 225752
rect 314016 225700 314068 225752
rect 202788 225632 202840 225684
rect 342260 225632 342312 225684
rect 3424 225564 3476 225616
rect 120172 225564 120224 225616
rect 210424 225564 210476 225616
rect 485044 225564 485096 225616
rect 222200 224952 222252 225004
rect 222936 224952 222988 225004
rect 289820 224952 289872 225004
rect 290464 224952 290516 225004
rect 52092 224884 52144 224936
rect 318064 224884 318116 224936
rect 55864 224816 55916 224868
rect 258080 224816 258132 224868
rect 258724 224816 258776 224868
rect 141516 224748 141568 224800
rect 296720 224816 296772 224868
rect 297364 224816 297416 224868
rect 75920 224680 75972 224732
rect 213920 224680 213972 224732
rect 213920 224408 213972 224460
rect 214656 224408 214708 224460
rect 126428 224272 126480 224324
rect 231124 224272 231176 224324
rect 100852 224204 100904 224256
rect 255412 224204 255464 224256
rect 276664 224204 276716 224256
rect 478880 224204 478932 224256
rect 82084 223524 82136 223576
rect 313280 223524 313332 223576
rect 313924 223524 313976 223576
rect 70492 223456 70544 223508
rect 201500 223456 201552 223508
rect 202420 223456 202472 223508
rect 148508 223388 148560 223440
rect 238760 223388 238812 223440
rect 239404 223388 239456 223440
rect 177396 222980 177448 223032
rect 232504 222980 232556 223032
rect 122104 222912 122156 222964
rect 254032 222912 254084 222964
rect 301504 222912 301556 222964
rect 495716 222912 495768 222964
rect 60464 222844 60516 222896
rect 162216 222844 162268 222896
rect 195796 222844 195848 222896
rect 471244 222844 471296 222896
rect 154028 222096 154080 222148
rect 309140 222096 309192 222148
rect 309876 222096 309928 222148
rect 79232 222028 79284 222080
rect 218704 222028 218756 222080
rect 73804 221960 73856 222012
rect 182088 221960 182140 222012
rect 158076 221892 158128 221944
rect 237380 221892 237432 221944
rect 92572 221552 92624 221604
rect 228456 221552 228508 221604
rect 182088 221484 182140 221536
rect 347872 221484 347924 221536
rect 192944 221416 192996 221468
rect 510712 221416 510764 221468
rect 247040 220804 247092 220856
rect 323676 220804 323728 220856
rect 156696 220736 156748 220788
rect 314108 220736 314160 220788
rect 429844 220736 429896 220788
rect 431224 220736 431276 220788
rect 93952 220668 94004 220720
rect 247040 220668 247092 220720
rect 84384 220600 84436 220652
rect 230480 220600 230532 220652
rect 231216 220600 231268 220652
rect 163688 220192 163740 220244
rect 259460 220192 259512 220244
rect 167736 220124 167788 220176
rect 289084 220124 289136 220176
rect 68928 220056 68980 220108
rect 253940 220056 253992 220108
rect 293224 220056 293276 220108
rect 429844 220056 429896 220108
rect 88984 219376 89036 219428
rect 266360 219376 266412 219428
rect 84292 219308 84344 219360
rect 228548 219308 228600 219360
rect 172428 218900 172480 218952
rect 227076 218900 227128 218952
rect 134708 218832 134760 218884
rect 236644 218832 236696 218884
rect 138756 218764 138808 218816
rect 263600 218764 263652 218816
rect 147128 218696 147180 218748
rect 278780 218696 278832 218748
rect 520924 218696 520976 218748
rect 579804 218696 579856 218748
rect 266360 218016 266412 218068
rect 267004 218016 267056 218068
rect 107752 217948 107804 218000
rect 283564 217948 283616 218000
rect 131856 217540 131908 217592
rect 238208 217540 238260 217592
rect 93860 217472 93912 217524
rect 249892 217472 249944 217524
rect 77300 217404 77352 217456
rect 249064 217404 249116 217456
rect 237380 217336 237432 217388
rect 483020 217336 483072 217388
rect 177856 217268 177908 217320
rect 436100 217268 436152 217320
rect 191748 216656 191800 216708
rect 198188 216656 198240 216708
rect 114560 216588 114612 216640
rect 295340 216588 295392 216640
rect 57612 216520 57664 216572
rect 233240 216520 233292 216572
rect 198648 215976 198700 216028
rect 325884 215976 325936 216028
rect 175096 215908 175148 215960
rect 497464 215908 497516 215960
rect 295340 215296 295392 215348
rect 295984 215296 296036 215348
rect 3332 215228 3384 215280
rect 14464 215228 14516 215280
rect 103704 215228 103756 215280
rect 271880 215228 271932 215280
rect 83464 215160 83516 215212
rect 208400 215160 208452 215212
rect 208400 214820 208452 214872
rect 209044 214820 209096 214872
rect 166264 214752 166316 214804
rect 240784 214752 240836 214804
rect 271880 214752 271932 214804
rect 272524 214752 272576 214804
rect 184756 214684 184808 214736
rect 389824 214684 389876 214736
rect 41236 214616 41288 214668
rect 270500 214616 270552 214668
rect 157984 214548 158036 214600
rect 216036 214548 216088 214600
rect 233240 214548 233292 214600
rect 486424 214548 486476 214600
rect 102232 213868 102284 213920
rect 273260 213868 273312 213920
rect 273904 213868 273956 213920
rect 176016 213392 176068 213444
rect 291844 213392 291896 213444
rect 74540 213324 74592 213376
rect 246304 213324 246356 213376
rect 56508 213256 56560 213308
rect 258264 213256 258316 213308
rect 190276 213188 190328 213240
rect 393964 213188 394016 213240
rect 184296 211896 184348 211948
rect 256976 211896 257028 211948
rect 258724 211896 258776 211948
rect 342904 211896 342956 211948
rect 106924 211828 106976 211880
rect 274640 211828 274692 211880
rect 118700 211760 118752 211812
rect 307760 211760 307812 211812
rect 432604 211080 432656 211132
rect 446404 211080 446456 211132
rect 431960 210672 432012 210724
rect 432604 210672 432656 210724
rect 115940 210536 115992 210588
rect 245016 210536 245068 210588
rect 86224 210468 86276 210520
rect 224960 210468 225012 210520
rect 304264 210468 304316 210520
rect 498384 210468 498436 210520
rect 179236 210400 179288 210452
rect 417424 210400 417476 210452
rect 447784 210400 447836 210452
rect 480260 210400 480312 210452
rect 104900 209720 104952 209772
rect 281540 209720 281592 209772
rect 113180 209652 113232 209704
rect 179328 209652 179380 209704
rect 133236 209244 133288 209296
rect 240876 209244 240928 209296
rect 179328 209176 179380 209228
rect 338120 209176 338172 209228
rect 169668 209108 169720 209160
rect 367744 209108 367796 209160
rect 11704 209040 11756 209092
rect 111064 209040 111116 209092
rect 218796 209040 218848 209092
rect 494244 209040 494296 209092
rect 281540 208360 281592 208412
rect 282276 208360 282328 208412
rect 95240 208292 95292 208344
rect 260840 208292 260892 208344
rect 197268 207952 197320 208004
rect 238024 207952 238076 208004
rect 165528 207884 165580 207936
rect 222844 207884 222896 207936
rect 214656 207816 214708 207868
rect 329932 207816 329984 207868
rect 89720 207748 89772 207800
rect 252744 207748 252796 207800
rect 135904 207680 135956 207732
rect 360200 207680 360252 207732
rect 46756 207612 46808 207664
rect 214564 207612 214616 207664
rect 239404 207612 239456 207664
rect 514760 207612 514812 207664
rect 260840 207068 260892 207120
rect 261484 207068 261536 207120
rect 92480 206932 92532 206984
rect 249800 206932 249852 206984
rect 346492 207000 346544 207052
rect 100760 206388 100812 206440
rect 255504 206388 255556 206440
rect 63316 206320 63368 206372
rect 282184 206320 282236 206372
rect 180708 206252 180760 206304
rect 505100 206252 505152 206304
rect 514760 206252 514812 206304
rect 515404 206252 515456 206304
rect 580172 206252 580224 206304
rect 107660 205572 107712 205624
rect 285680 205572 285732 205624
rect 285680 205096 285732 205148
rect 286416 205096 286468 205148
rect 222936 204960 222988 205012
rect 320916 204960 320968 205012
rect 65892 204892 65944 204944
rect 240968 204892 241020 204944
rect 262956 204892 263008 204944
rect 494152 204892 494204 204944
rect 98000 204212 98052 204264
rect 146944 204212 146996 204264
rect 156604 203736 156656 203788
rect 266360 203736 266412 203788
rect 149704 203668 149756 203720
rect 280804 203668 280856 203720
rect 99380 203600 99432 203652
rect 254124 203600 254176 203652
rect 146944 203532 146996 203584
rect 392584 203532 392636 203584
rect 217324 202376 217376 202428
rect 321560 202376 321612 202428
rect 123760 202308 123812 202360
rect 262220 202308 262272 202360
rect 45468 202240 45520 202292
rect 232596 202240 232648 202292
rect 69112 202172 69164 202224
rect 280160 202172 280212 202224
rect 322204 202172 322256 202224
rect 328644 202172 328696 202224
rect 159548 202104 159600 202156
rect 381544 202104 381596 202156
rect 126336 200880 126388 200932
rect 242256 200880 242308 200932
rect 269764 200880 269816 200932
rect 327264 200880 327316 200932
rect 86960 200812 87012 200864
rect 274732 200812 274784 200864
rect 144184 200744 144236 200796
rect 509332 200744 509384 200796
rect 145656 199588 145708 199640
rect 276664 199588 276716 199640
rect 104164 199520 104216 199572
rect 260932 199520 260984 199572
rect 53656 199452 53708 199504
rect 238116 199452 238168 199504
rect 261484 199452 261536 199504
rect 321836 199452 321888 199504
rect 211804 199384 211856 199436
rect 514760 199384 514812 199436
rect 181536 198228 181588 198280
rect 213184 198228 213236 198280
rect 162216 198160 162268 198212
rect 262312 198160 262364 198212
rect 102140 198092 102192 198144
rect 250076 198092 250128 198144
rect 67456 198024 67508 198076
rect 251180 198024 251232 198076
rect 127624 197956 127676 198008
rect 195336 197956 195388 198008
rect 213276 197956 213328 198008
rect 451280 197956 451332 198008
rect 238208 196800 238260 196852
rect 271972 196800 272024 196852
rect 126244 196732 126296 196784
rect 184296 196732 184348 196784
rect 242164 196732 242216 196784
rect 328736 196732 328788 196784
rect 142896 196664 142948 196716
rect 243544 196664 243596 196716
rect 160928 196596 160980 196648
rect 502340 196596 502392 196648
rect 129096 195508 129148 195560
rect 213276 195508 213328 195560
rect 194508 195440 194560 195492
rect 336924 195440 336976 195492
rect 70400 195372 70452 195424
rect 254216 195372 254268 195424
rect 138664 195304 138716 195356
rect 352012 195304 352064 195356
rect 78680 195236 78732 195288
rect 267740 195236 267792 195288
rect 290464 195236 290516 195288
rect 507952 195236 508004 195288
rect 151084 193944 151136 193996
rect 286324 193944 286376 193996
rect 323584 193944 323636 193996
rect 341064 193944 341116 193996
rect 111800 193876 111852 193928
rect 252652 193876 252704 193928
rect 286416 193876 286468 193928
rect 330116 193876 330168 193928
rect 129004 193808 129056 193860
rect 369860 193808 369912 193860
rect 188436 192720 188488 192772
rect 245108 192720 245160 192772
rect 224868 192652 224920 192704
rect 318064 192652 318116 192704
rect 130384 192584 130436 192636
rect 264980 192584 265032 192636
rect 272524 192584 272576 192636
rect 325792 192584 325844 192636
rect 176108 192516 176160 192568
rect 343824 192516 343876 192568
rect 137376 192448 137428 192500
rect 357532 192448 357584 192500
rect 360844 192448 360896 192500
rect 517520 192448 517572 192500
rect 134524 191156 134576 191208
rect 269120 191156 269172 191208
rect 72424 191088 72476 191140
rect 273444 191088 273496 191140
rect 133144 190068 133196 190120
rect 200764 190068 200816 190120
rect 228548 190068 228600 190120
rect 309784 190068 309836 190120
rect 164976 190000 165028 190052
rect 258172 190000 258224 190052
rect 193128 189932 193180 189984
rect 335636 189932 335688 189984
rect 76564 189864 76616 189916
rect 260840 189864 260892 189916
rect 52276 189796 52328 189848
rect 267832 189796 267884 189848
rect 297364 189796 297416 189848
rect 501144 189796 501196 189848
rect 183468 189728 183520 189780
rect 460112 189728 460164 189780
rect 268384 189048 268436 189100
rect 269212 189048 269264 189100
rect 3424 188980 3476 189032
rect 53104 188980 53156 189032
rect 151176 188504 151228 188556
rect 270684 188504 270736 188556
rect 142804 188436 142856 188488
rect 196624 188436 196676 188488
rect 218704 188436 218756 188488
rect 339592 188436 339644 188488
rect 84200 188368 84252 188420
rect 249984 188368 250036 188420
rect 320824 188368 320876 188420
rect 334072 188368 334124 188420
rect 47952 188300 48004 188352
rect 256792 188300 256844 188352
rect 265624 188300 265676 188352
rect 494336 188300 494388 188352
rect 235264 187280 235316 187332
rect 308404 187280 308456 187332
rect 173256 187212 173308 187264
rect 261024 187212 261076 187264
rect 147036 187144 147088 187196
rect 189816 187144 189868 187196
rect 231216 187144 231268 187196
rect 335544 187144 335596 187196
rect 110420 187076 110472 187128
rect 249800 187076 249852 187128
rect 124864 187008 124916 187060
rect 270592 187008 270644 187060
rect 173348 186940 173400 186992
rect 342352 186940 342404 186992
rect 358084 186940 358136 186992
rect 513380 186940 513432 186992
rect 148324 185784 148376 185836
rect 210424 185784 210476 185836
rect 213368 185784 213420 185836
rect 259552 185784 259604 185836
rect 177948 185716 178000 185768
rect 345204 185716 345256 185768
rect 141424 185648 141476 185700
rect 351184 185648 351236 185700
rect 422944 185648 422996 185700
rect 450544 185648 450596 185700
rect 119344 185580 119396 185632
rect 273352 185580 273404 185632
rect 278044 185580 278096 185632
rect 503904 185580 503956 185632
rect 318616 185512 318668 185564
rect 320180 185512 320232 185564
rect 102048 184968 102100 185020
rect 169024 184968 169076 185020
rect 100668 184900 100720 184952
rect 173164 184900 173216 184952
rect 232596 184424 232648 184476
rect 266544 184424 266596 184476
rect 145564 184356 145616 184408
rect 273260 184356 273312 184408
rect 140136 184288 140188 184340
rect 278044 184288 278096 184340
rect 345664 184288 345716 184340
rect 443920 184288 443972 184340
rect 468484 184288 468536 184340
rect 510804 184288 510856 184340
rect 171784 184220 171836 184272
rect 345296 184220 345348 184272
rect 400864 184220 400916 184272
rect 505192 184220 505244 184272
rect 155224 184152 155276 184204
rect 202144 184152 202196 184204
rect 227076 184152 227128 184204
rect 507860 184152 507912 184204
rect 128268 183608 128320 183660
rect 180248 183608 180300 183660
rect 107568 183540 107620 183592
rect 196716 183540 196768 183592
rect 403624 183472 403676 183524
rect 404268 183472 404320 183524
rect 236644 183132 236696 183184
rect 263784 183132 263836 183184
rect 228364 183064 228416 183116
rect 265072 183064 265124 183116
rect 251916 182996 251968 183048
rect 345020 182996 345072 183048
rect 195244 182928 195296 182980
rect 313832 182928 313884 182980
rect 200856 182860 200908 182912
rect 338304 182860 338356 182912
rect 57704 182792 57756 182844
rect 262404 182792 262456 182844
rect 314016 182792 314068 182844
rect 331496 182792 331548 182844
rect 419356 182792 419408 182844
rect 580356 182792 580408 182844
rect 132408 182452 132460 182504
rect 164976 182452 165028 182504
rect 105728 182384 105780 182436
rect 170772 182384 170824 182436
rect 119712 182316 119764 182368
rect 204996 182316 205048 182368
rect 489184 182316 489236 182368
rect 490564 182316 490616 182368
rect 110696 182248 110748 182300
rect 196808 182248 196860 182300
rect 400864 182248 400916 182300
rect 494060 182248 494112 182300
rect 123300 182180 123352 182232
rect 214656 182180 214708 182232
rect 404268 182180 404320 182232
rect 580264 182180 580316 182232
rect 454684 182112 454736 182164
rect 455604 182112 455656 182164
rect 461584 182112 461636 182164
rect 462596 182112 462648 182164
rect 471244 182112 471296 182164
rect 476580 182112 476632 182164
rect 485044 182112 485096 182164
rect 485780 182112 485832 182164
rect 245016 181772 245068 181824
rect 263692 181772 263744 181824
rect 486424 181772 486476 181824
rect 492864 181772 492916 181824
rect 168288 181704 168340 181756
rect 216128 181704 216180 181756
rect 228456 181704 228508 181756
rect 259736 181704 259788 181756
rect 307024 181704 307076 181756
rect 336740 181704 336792 181756
rect 475384 181704 475436 181756
rect 488632 181704 488684 181756
rect 170680 181636 170732 181688
rect 251272 181636 251324 181688
rect 251824 181636 251876 181688
rect 341156 181636 341208 181688
rect 414664 181636 414716 181688
rect 441620 181636 441672 181688
rect 457444 181636 457496 181688
rect 474188 181636 474240 181688
rect 482284 181636 482336 181688
rect 505284 181636 505336 181688
rect 159364 181568 159416 181620
rect 209044 181568 209096 181620
rect 233884 181568 233936 181620
rect 334164 181568 334216 181620
rect 352564 181568 352616 181620
rect 448612 181568 448664 181620
rect 464344 181568 464396 181620
rect 503996 181568 504048 181620
rect 137468 181500 137520 181552
rect 249156 181500 249208 181552
rect 262864 181500 262916 181552
rect 446404 181500 446456 181552
rect 449164 181500 449216 181552
rect 502616 181500 502668 181552
rect 180616 181432 180668 181484
rect 497004 181432 497056 181484
rect 130936 181024 130988 181076
rect 166540 181024 166592 181076
rect 129464 180956 129516 181008
rect 167920 180956 167972 181008
rect 121184 180888 121236 180940
rect 167828 180888 167880 180940
rect 116952 180820 117004 180872
rect 170864 180820 170916 180872
rect 246304 180412 246356 180464
rect 272064 180412 272116 180464
rect 169208 180344 169260 180396
rect 251364 180344 251416 180396
rect 151268 180276 151320 180328
rect 266452 180276 266504 180328
rect 273904 180276 273956 180328
rect 332876 180276 332928 180328
rect 490656 180276 490708 180328
rect 501236 180276 501288 180328
rect 187056 180208 187108 180260
rect 324504 180208 324556 180260
rect 411904 180208 411956 180260
rect 506572 180208 506624 180260
rect 187148 180140 187200 180192
rect 349252 180140 349304 180192
rect 359464 180140 359516 180192
rect 509240 180140 509292 180192
rect 160744 180072 160796 180124
rect 195244 180072 195296 180124
rect 222844 180072 222896 180124
rect 503812 180072 503864 180124
rect 134708 179596 134760 179648
rect 165436 179596 165488 179648
rect 126060 179528 126112 179580
rect 168012 179528 168064 179580
rect 115848 179460 115900 179512
rect 166264 179460 166316 179512
rect 109960 179392 110012 179444
rect 169300 179392 169352 179444
rect 309876 178984 309928 179036
rect 325976 178984 326028 179036
rect 170404 178916 170456 178968
rect 251456 178916 251508 178968
rect 313924 178916 313976 178968
rect 332692 178916 332744 178968
rect 244924 178848 244976 178900
rect 336832 178848 336884 178900
rect 166356 178780 166408 178832
rect 267924 178780 267976 178832
rect 295984 178780 296036 178832
rect 327172 178780 327224 178832
rect 123484 178712 123536 178764
rect 249340 178712 249392 178764
rect 257344 178712 257396 178764
rect 346584 178712 346636 178764
rect 162124 178644 162176 178696
rect 198004 178644 198056 178696
rect 202328 178644 202380 178696
rect 339684 178644 339736 178696
rect 497464 178644 497516 178696
rect 502524 178644 502576 178696
rect 503628 178644 503680 178696
rect 148232 178236 148284 178288
rect 170496 178236 170548 178288
rect 114376 178168 114428 178220
rect 166448 178168 166500 178220
rect 112260 178100 112312 178152
rect 171968 178100 172020 178152
rect 97816 178032 97868 178084
rect 177396 178032 177448 178084
rect 347044 178032 347096 178084
rect 416780 178032 416832 178084
rect 503628 178032 503680 178084
rect 580172 178032 580224 178084
rect 323676 177964 323728 178016
rect 327080 177964 327132 178016
rect 242256 177624 242308 177676
rect 256884 177624 256936 177676
rect 312544 177624 312596 177676
rect 321744 177624 321796 177676
rect 226984 177556 227036 177608
rect 249248 177556 249300 177608
rect 318708 177556 318760 177608
rect 331404 177556 331456 177608
rect 231124 177488 231176 177540
rect 258356 177488 258408 177540
rect 283564 177488 283616 177540
rect 350632 177488 350684 177540
rect 190368 177420 190420 177472
rect 294696 177420 294748 177472
rect 318064 177420 318116 177472
rect 332784 177420 332836 177472
rect 202420 177352 202472 177404
rect 323124 177352 323176 177404
rect 14464 177284 14516 177336
rect 109684 177284 109736 177336
rect 203524 177284 203576 177336
rect 338212 177284 338264 177336
rect 128176 177012 128228 177064
rect 160100 177012 160152 177064
rect 124496 176944 124548 176996
rect 165252 176944 165304 176996
rect 158904 176876 158956 176928
rect 214748 176876 214800 176928
rect 108120 176808 108172 176860
rect 169116 176808 169168 176860
rect 136088 176740 136140 176792
rect 201592 176740 201644 176792
rect 496912 176740 496964 176792
rect 501052 176740 501104 176792
rect 133144 176672 133196 176724
rect 205640 176672 205692 176724
rect 342996 176672 343048 176724
rect 416780 176672 416832 176724
rect 496820 176672 496872 176724
rect 499764 176672 499816 176724
rect 201592 176604 201644 176656
rect 213920 176604 213972 176656
rect 313832 176604 313884 176656
rect 321468 176604 321520 176656
rect 118424 176264 118476 176316
rect 166356 176264 166408 176316
rect 163504 176196 163556 176248
rect 211804 176196 211856 176248
rect 160100 176128 160152 176180
rect 214104 176128 214156 176180
rect 102048 176060 102100 176112
rect 171784 176060 171836 176112
rect 238116 176060 238168 176112
rect 256700 176060 256752 176112
rect 307668 176060 307720 176112
rect 349344 176060 349396 176112
rect 98368 175992 98420 176044
rect 170404 175992 170456 176044
rect 171876 175992 171928 176044
rect 258080 175992 258132 176044
rect 267004 175992 267056 176044
rect 323032 175992 323084 176044
rect 121920 175924 121972 175976
rect 195428 175924 195480 175976
rect 238024 175924 238076 175976
rect 396724 175924 396776 175976
rect 240784 175788 240836 175840
rect 248052 175788 248104 175840
rect 496820 175584 496872 175636
rect 498476 175584 498528 175636
rect 165436 175176 165488 175228
rect 213920 175176 213972 175228
rect 205640 175108 205692 175160
rect 214012 175108 214064 175160
rect 252468 175108 252520 175160
rect 258172 175108 258224 175160
rect 165252 174496 165304 174548
rect 214932 174496 214984 174548
rect 284944 174020 284996 174072
rect 307576 174020 307628 174072
rect 265808 173952 265860 174004
rect 307668 173952 307720 174004
rect 263048 173884 263100 173936
rect 307484 173884 307536 173936
rect 358084 173884 358136 173936
rect 416780 173884 416832 173936
rect 164976 173816 165028 173868
rect 213920 173816 213972 173868
rect 252468 173816 252520 173868
rect 262404 173816 262456 173868
rect 166540 173748 166592 173800
rect 214012 173748 214064 173800
rect 302884 172660 302936 172712
rect 307484 172660 307536 172712
rect 298744 172592 298796 172644
rect 307668 172592 307720 172644
rect 276756 172524 276808 172576
rect 307300 172524 307352 172576
rect 167920 172456 167972 172508
rect 213920 172456 213972 172508
rect 252376 172456 252428 172508
rect 261024 172456 261076 172508
rect 252468 172116 252520 172168
rect 258080 172116 258132 172168
rect 261484 171776 261536 171828
rect 307392 171776 307444 171828
rect 278228 171164 278280 171216
rect 307668 171164 307720 171216
rect 265716 171096 265768 171148
rect 307116 171096 307168 171148
rect 324964 171096 325016 171148
rect 327080 171096 327132 171148
rect 353944 171096 353996 171148
rect 416780 171096 416832 171148
rect 168012 171028 168064 171080
rect 214012 171028 214064 171080
rect 252468 171028 252520 171080
rect 263600 171028 263652 171080
rect 180248 170960 180300 171012
rect 213920 170960 213972 171012
rect 252376 170960 252428 171012
rect 262312 170960 262364 171012
rect 252468 170552 252520 170604
rect 256700 170552 256752 170604
rect 297456 169872 297508 169924
rect 306748 169872 306800 169924
rect 267188 169804 267240 169856
rect 307668 169804 307720 169856
rect 261668 169736 261720 169788
rect 307484 169736 307536 169788
rect 324320 169668 324372 169720
rect 335636 169668 335688 169720
rect 300308 168444 300360 168496
rect 307668 168444 307720 168496
rect 259000 168376 259052 168428
rect 307576 168376 307628 168428
rect 414664 168376 414716 168428
rect 416780 168376 416832 168428
rect 167828 168308 167880 168360
rect 214012 168308 214064 168360
rect 252376 168308 252428 168360
rect 256884 168308 256936 168360
rect 324320 168308 324372 168360
rect 357440 168308 357492 168360
rect 496820 168308 496872 168360
rect 502432 168308 502484 168360
rect 503628 168308 503680 168360
rect 195428 168240 195480 168292
rect 213920 168240 213972 168292
rect 252468 168036 252520 168088
rect 259460 168036 259512 168088
rect 291936 167628 291988 167680
rect 306564 167628 306616 167680
rect 338764 167628 338816 167680
rect 348424 167628 348476 167680
rect 503628 167628 503680 167680
rect 543004 167628 543056 167680
rect 251272 167220 251324 167272
rect 251548 167220 251600 167272
rect 268384 167084 268436 167136
rect 307668 167084 307720 167136
rect 264428 167016 264480 167068
rect 307300 167016 307352 167068
rect 166356 166948 166408 167000
rect 214104 166948 214156 167000
rect 170864 166880 170916 166932
rect 214012 166880 214064 166932
rect 204996 166812 205048 166864
rect 213920 166812 213972 166864
rect 252376 166676 252428 166728
rect 258264 166676 258316 166728
rect 252468 166608 252520 166660
rect 258356 166608 258408 166660
rect 295984 166336 296036 166388
rect 306656 166336 306708 166388
rect 264336 166268 264388 166320
rect 306932 166268 306984 166320
rect 496820 166268 496872 166320
rect 504088 166268 504140 166320
rect 252468 166064 252520 166116
rect 259736 166064 259788 166116
rect 271144 165588 271196 165640
rect 306748 165588 306800 165640
rect 338764 165588 338816 165640
rect 416780 165588 416832 165640
rect 504088 165588 504140 165640
rect 525064 165588 525116 165640
rect 535460 165588 535512 165640
rect 580172 165588 580224 165640
rect 166264 165520 166316 165572
rect 213920 165520 213972 165572
rect 252468 165520 252520 165572
rect 259552 165520 259604 165572
rect 324320 165520 324372 165572
rect 339684 165520 339736 165572
rect 166448 165452 166500 165504
rect 214012 165452 214064 165504
rect 252376 165452 252428 165504
rect 256792 165452 256844 165504
rect 324412 165452 324464 165504
rect 332876 165452 332928 165504
rect 258724 164840 258776 164892
rect 307484 164840 307536 164892
rect 496820 164840 496872 164892
rect 503996 164840 504048 164892
rect 301596 164296 301648 164348
rect 307116 164296 307168 164348
rect 269856 164228 269908 164280
rect 307668 164228 307720 164280
rect 359464 164228 359516 164280
rect 416780 164228 416832 164280
rect 496360 164228 496412 164280
rect 530584 164228 530636 164280
rect 3240 164160 3292 164212
rect 33784 164160 33836 164212
rect 171968 164160 172020 164212
rect 213920 164160 213972 164212
rect 252468 164160 252520 164212
rect 270500 164160 270552 164212
rect 324320 164160 324372 164212
rect 334164 164160 334216 164212
rect 496820 164160 496872 164212
rect 509332 164160 509384 164212
rect 535460 164160 535512 164212
rect 252376 164092 252428 164144
rect 263784 164092 263836 164144
rect 324412 164092 324464 164144
rect 331496 164092 331548 164144
rect 272524 163548 272576 163600
rect 306564 163548 306616 163600
rect 257620 163480 257672 163532
rect 307576 163480 307628 163532
rect 293316 162868 293368 162920
rect 307668 162868 307720 162920
rect 340144 162868 340196 162920
rect 416780 162868 416832 162920
rect 169300 162800 169352 162852
rect 214012 162800 214064 162852
rect 252376 162800 252428 162852
rect 266544 162800 266596 162852
rect 324320 162800 324372 162852
rect 334072 162800 334124 162852
rect 496820 162800 496872 162852
rect 515404 162800 515456 162852
rect 196808 162732 196860 162784
rect 213920 162732 213972 162784
rect 252468 162732 252520 162784
rect 264980 162732 265032 162784
rect 302976 161644 303028 161696
rect 307392 161644 307444 161696
rect 299020 161576 299072 161628
rect 307484 161576 307536 161628
rect 269948 161508 270000 161560
rect 307576 161508 307628 161560
rect 262864 161440 262916 161492
rect 307668 161440 307720 161492
rect 334808 161440 334860 161492
rect 416780 161440 416832 161492
rect 169116 161372 169168 161424
rect 213920 161372 213972 161424
rect 252468 161372 252520 161424
rect 263692 161372 263744 161424
rect 496912 161372 496964 161424
rect 512092 161372 512144 161424
rect 196716 161304 196768 161356
rect 214012 161304 214064 161356
rect 252376 160488 252428 160540
rect 259644 160488 259696 160540
rect 287980 160216 288032 160268
rect 307576 160216 307628 160268
rect 260472 160148 260524 160200
rect 307668 160148 307720 160200
rect 260104 160080 260156 160132
rect 306564 160080 306616 160132
rect 167736 160012 167788 160064
rect 214012 160012 214064 160064
rect 252468 160012 252520 160064
rect 273444 160012 273496 160064
rect 496912 160012 496964 160064
rect 536840 160012 536892 160064
rect 170772 159944 170824 159996
rect 213920 159944 213972 159996
rect 497004 159944 497056 159996
rect 503720 159944 503772 159996
rect 273904 158856 273956 158908
rect 306932 158856 306984 158908
rect 264520 158788 264572 158840
rect 307668 158788 307720 158840
rect 260380 158720 260432 158772
rect 307576 158720 307628 158772
rect 344284 158720 344336 158772
rect 416780 158720 416832 158772
rect 171784 158652 171836 158704
rect 213920 158652 213972 158704
rect 252468 158652 252520 158704
rect 260932 158652 260984 158704
rect 324412 158652 324464 158704
rect 335452 158652 335504 158704
rect 496912 158652 496964 158704
rect 517612 158652 517664 158704
rect 544384 158652 544436 158704
rect 324320 158516 324372 158568
rect 327448 158516 327500 158568
rect 253388 157972 253440 158024
rect 307208 157972 307260 158024
rect 283564 157428 283616 157480
rect 307484 157428 307536 157480
rect 257344 157360 257396 157412
rect 306748 157360 306800 157412
rect 169024 157292 169076 157344
rect 213920 157292 213972 157344
rect 252468 157292 252520 157344
rect 270684 157292 270736 157344
rect 496912 157292 496964 157344
rect 582380 157292 582432 157344
rect 173164 157224 173216 157276
rect 214012 157224 214064 157276
rect 253204 156612 253256 156664
rect 267832 156612 267884 156664
rect 324320 156408 324372 156460
rect 327264 156408 327316 156460
rect 281080 156068 281132 156120
rect 307668 156068 307720 156120
rect 267004 156000 267056 156052
rect 307576 156000 307628 156052
rect 260288 155932 260340 155984
rect 306564 155932 306616 155984
rect 336004 155932 336056 155984
rect 416780 155932 416832 155984
rect 170404 155864 170456 155916
rect 213920 155864 213972 155916
rect 252468 155864 252520 155916
rect 265072 155864 265124 155916
rect 496912 155864 496964 155916
rect 519544 155864 519596 155916
rect 177396 155796 177448 155848
rect 214012 155796 214064 155848
rect 252376 155796 252428 155848
rect 255412 155796 255464 155848
rect 327724 155184 327776 155236
rect 333980 155184 334032 155236
rect 304356 154708 304408 154760
rect 307668 154708 307720 154760
rect 271236 154640 271288 154692
rect 306564 154640 306616 154692
rect 261760 154572 261812 154624
rect 307300 154572 307352 154624
rect 332048 154572 332100 154624
rect 416780 154572 416832 154624
rect 252468 154504 252520 154556
rect 274732 154504 274784 154556
rect 324412 154504 324464 154556
rect 332784 154504 332836 154556
rect 497004 154504 497056 154556
rect 505284 154504 505336 154556
rect 251456 154436 251508 154488
rect 254216 154436 254268 154488
rect 324320 154436 324372 154488
rect 328736 154436 328788 154488
rect 496912 154436 496964 154488
rect 502616 154436 502668 154488
rect 167644 153824 167696 153876
rect 208400 153824 208452 153876
rect 275376 153348 275428 153400
rect 307576 153348 307628 153400
rect 258816 153280 258868 153332
rect 307668 153280 307720 153332
rect 173164 153212 173216 153264
rect 213920 153212 213972 153264
rect 258908 153212 258960 153264
rect 307300 153212 307352 153264
rect 356796 153212 356848 153264
rect 416780 153212 416832 153264
rect 252284 153144 252336 153196
rect 271972 153144 272024 153196
rect 324320 153144 324372 153196
rect 330024 153144 330076 153196
rect 496912 153144 496964 153196
rect 507952 153144 508004 153196
rect 252468 153076 252520 153128
rect 269212 153076 269264 153128
rect 252376 153008 252428 153060
rect 267924 153008 267976 153060
rect 296076 151920 296128 151972
rect 307668 151920 307720 151972
rect 206376 151852 206428 151904
rect 213920 151852 213972 151904
rect 268476 151852 268528 151904
rect 307576 151852 307628 151904
rect 199384 151784 199436 151836
rect 214012 151784 214064 151836
rect 254584 151784 254636 151836
rect 307484 151784 307536 151836
rect 324412 151716 324464 151768
rect 347872 151716 347924 151768
rect 324320 151648 324372 151700
rect 330116 151648 330168 151700
rect 252468 151444 252520 151496
rect 255596 151444 255648 151496
rect 251456 151308 251508 151360
rect 254124 151308 254176 151360
rect 251824 151104 251876 151156
rect 283564 151104 283616 151156
rect 255964 151036 256016 151088
rect 306656 151036 306708 151088
rect 279516 150560 279568 150612
rect 307576 150560 307628 150612
rect 208492 150492 208544 150544
rect 214012 150492 214064 150544
rect 298928 150492 298980 150544
rect 307668 150492 307720 150544
rect 205088 150424 205140 150476
rect 213920 150424 213972 150476
rect 360844 150424 360896 150476
rect 416780 150424 416832 150476
rect 3424 150356 3476 150408
rect 25504 150356 25556 150408
rect 170496 150356 170548 150408
rect 214012 150356 214064 150408
rect 252468 150356 252520 150408
rect 278780 150356 278832 150408
rect 324320 150356 324372 150408
rect 345296 150356 345348 150408
rect 496820 150356 496872 150408
rect 503904 150356 503956 150408
rect 208400 150288 208452 150340
rect 213920 150288 213972 150340
rect 251364 150288 251416 150340
rect 254032 150288 254084 150340
rect 324412 150288 324464 150340
rect 331404 150288 331456 150340
rect 324596 149676 324648 149728
rect 343824 149676 343876 149728
rect 304264 149200 304316 149252
rect 307668 149200 307720 149252
rect 283656 149132 283708 149184
rect 306748 149132 306800 149184
rect 254860 149064 254912 149116
rect 307576 149064 307628 149116
rect 363604 149064 363656 149116
rect 416780 149064 416832 149116
rect 252468 148996 252520 149048
rect 272064 148996 272116 149048
rect 324412 148996 324464 149048
rect 335544 148996 335596 149048
rect 252376 148928 252428 148980
rect 256976 148928 257028 148980
rect 324320 148928 324372 148980
rect 328644 148928 328696 148980
rect 289268 147772 289320 147824
rect 306932 147772 306984 147824
rect 265624 147704 265676 147756
rect 307576 147704 307628 147756
rect 254768 147636 254820 147688
rect 307668 147636 307720 147688
rect 332508 147636 332560 147688
rect 416780 147636 416832 147688
rect 252468 147568 252520 147620
rect 270592 147568 270644 147620
rect 324320 147568 324372 147620
rect 340880 147568 340932 147620
rect 496820 147568 496872 147620
rect 505192 147568 505244 147620
rect 251364 147500 251416 147552
rect 253940 147500 253992 147552
rect 252100 147432 252152 147484
rect 255504 147432 255556 147484
rect 285128 146412 285180 146464
rect 307576 146412 307628 146464
rect 200856 146344 200908 146396
rect 213920 146344 213972 146396
rect 272616 146344 272668 146396
rect 307668 146344 307720 146396
rect 171784 146276 171836 146328
rect 214012 146276 214064 146328
rect 257528 146276 257580 146328
rect 306748 146276 306800 146328
rect 345664 146276 345716 146328
rect 416780 146276 416832 146328
rect 252376 146208 252428 146260
rect 267740 146208 267792 146260
rect 324320 146208 324372 146260
rect 356060 146208 356112 146260
rect 496820 146208 496872 146260
rect 510804 146208 510856 146260
rect 252468 146140 252520 146192
rect 260840 146140 260892 146192
rect 180248 145528 180300 145580
rect 215024 145528 215076 145580
rect 277032 145528 277084 145580
rect 307116 145528 307168 145580
rect 324412 145528 324464 145580
rect 338304 145528 338356 145580
rect 166264 144916 166316 144968
rect 213920 144916 213972 144968
rect 256148 144916 256200 144968
rect 307668 144916 307720 144968
rect 252376 144848 252428 144900
rect 269120 144848 269172 144900
rect 324320 144848 324372 144900
rect 345204 144848 345256 144900
rect 252468 144780 252520 144832
rect 262220 144780 262272 144832
rect 506572 144440 506624 144492
rect 507124 144440 507176 144492
rect 167736 144168 167788 144220
rect 208492 144168 208544 144220
rect 276940 144168 276992 144220
rect 307576 144168 307628 144220
rect 496820 144168 496872 144220
rect 506572 144168 506624 144220
rect 206468 143624 206520 143676
rect 213920 143624 213972 143676
rect 251916 143624 251968 143676
rect 260104 143624 260156 143676
rect 260196 143624 260248 143676
rect 307668 143624 307720 143676
rect 198096 143556 198148 143608
rect 214012 143556 214064 143608
rect 256056 143556 256108 143608
rect 306932 143556 306984 143608
rect 352656 143556 352708 143608
rect 416780 143556 416832 143608
rect 252468 143488 252520 143540
rect 266360 143488 266412 143540
rect 324320 143488 324372 143540
rect 328552 143488 328604 143540
rect 496820 143488 496872 143540
rect 510712 143488 510764 143540
rect 512644 143488 512696 143540
rect 252376 143420 252428 143472
rect 266452 143420 266504 143472
rect 253296 142808 253348 142860
rect 307576 142808 307628 142860
rect 209228 142196 209280 142248
rect 213920 142196 213972 142248
rect 269764 142196 269816 142248
rect 307668 142196 307720 142248
rect 167644 142128 167696 142180
rect 214012 142128 214064 142180
rect 256240 142128 256292 142180
rect 306564 142128 306616 142180
rect 333244 142128 333296 142180
rect 416872 142128 416924 142180
rect 324412 142060 324464 142112
rect 343640 142060 343692 142112
rect 353300 142060 353352 142112
rect 416780 142060 416832 142112
rect 324320 141992 324372 142044
rect 329840 141992 329892 142044
rect 252192 141448 252244 141500
rect 265808 141448 265860 141500
rect 253572 141380 253624 141432
rect 307024 141380 307076 141432
rect 334624 141380 334676 141432
rect 353300 141380 353352 141432
rect 304356 140904 304408 140956
rect 307484 140904 307536 140956
rect 204996 140836 205048 140888
rect 214012 140836 214064 140888
rect 286508 140836 286560 140888
rect 306564 140836 306616 140888
rect 496820 140836 496872 140888
rect 520188 140836 520240 140888
rect 521660 140836 521712 140888
rect 178776 140768 178828 140820
rect 213920 140768 213972 140820
rect 267096 140768 267148 140820
rect 307668 140768 307720 140820
rect 495348 140768 495400 140820
rect 502800 140768 502852 140820
rect 252468 140700 252520 140752
rect 273260 140700 273312 140752
rect 496820 140700 496872 140752
rect 502524 140700 502576 140752
rect 174636 140020 174688 140072
rect 214748 140020 214800 140072
rect 502800 140020 502852 140072
rect 580172 140020 580224 140072
rect 264244 139544 264296 139596
rect 307668 139544 307720 139596
rect 211896 139476 211948 139528
rect 214656 139476 214708 139528
rect 262956 139476 263008 139528
rect 307576 139476 307628 139528
rect 166356 139408 166408 139460
rect 213920 139408 213972 139460
rect 250628 139408 250680 139460
rect 307300 139408 307352 139460
rect 367836 139408 367888 139460
rect 416780 139408 416832 139460
rect 252468 139340 252520 139392
rect 280160 139340 280212 139392
rect 324320 139340 324372 139392
rect 346584 139340 346636 139392
rect 496820 139340 496872 139392
rect 520924 139340 520976 139392
rect 287796 138116 287848 138168
rect 307300 138116 307352 138168
rect 253204 138048 253256 138100
rect 306564 138048 306616 138100
rect 170404 137980 170456 138032
rect 213920 137980 213972 138032
rect 250536 137980 250588 138032
rect 307668 137980 307720 138032
rect 3240 137912 3292 137964
rect 15844 137912 15896 137964
rect 252468 137912 252520 137964
rect 274640 137912 274692 137964
rect 324412 137912 324464 137964
rect 339592 137912 339644 137964
rect 358820 137912 358872 137964
rect 416780 137912 416832 137964
rect 496820 137912 496872 137964
rect 548524 137912 548576 137964
rect 324320 137844 324372 137896
rect 336924 137844 336976 137896
rect 290464 137232 290516 137284
rect 307208 137232 307260 137284
rect 354036 137232 354088 137284
rect 358820 137232 358872 137284
rect 202420 136688 202472 136740
rect 213920 136688 213972 136740
rect 181536 136620 181588 136672
rect 214012 136620 214064 136672
rect 250444 136620 250496 136672
rect 307668 136620 307720 136672
rect 252284 136552 252336 136604
rect 284944 136552 284996 136604
rect 324412 136552 324464 136604
rect 351920 136552 351972 136604
rect 496912 136552 496964 136604
rect 508504 136552 508556 136604
rect 252468 136484 252520 136536
rect 271880 136484 271932 136536
rect 324320 136484 324372 136536
rect 338212 136484 338264 136536
rect 252376 136416 252428 136468
rect 263048 136416 263100 136468
rect 496820 136348 496872 136400
rect 501236 136348 501288 136400
rect 300124 135464 300176 135516
rect 307668 135464 307720 135516
rect 289176 135396 289228 135448
rect 307300 135396 307352 135448
rect 280988 135328 281040 135380
rect 307576 135328 307628 135380
rect 196716 135260 196768 135312
rect 213920 135260 213972 135312
rect 254676 135260 254728 135312
rect 306564 135260 306616 135312
rect 370504 135260 370556 135312
rect 416780 135260 416832 135312
rect 252376 135192 252428 135244
rect 302884 135192 302936 135244
rect 334716 135192 334768 135244
rect 417332 135192 417384 135244
rect 252468 135124 252520 135176
rect 276756 135124 276808 135176
rect 265808 134512 265860 134564
rect 307392 134512 307444 134564
rect 198280 133968 198332 134020
rect 214012 133968 214064 134020
rect 177396 133900 177448 133952
rect 213920 133900 213972 133952
rect 286416 133900 286468 133952
rect 306564 133900 306616 133952
rect 252468 133832 252520 133884
rect 298744 133832 298796 133884
rect 374644 133832 374696 133884
rect 419448 133832 419500 133884
rect 496820 133832 496872 133884
rect 512000 133832 512052 133884
rect 252284 133764 252336 133816
rect 295984 133764 296036 133816
rect 252376 133696 252428 133748
rect 265716 133696 265768 133748
rect 404268 133152 404320 133204
rect 419632 133152 419684 133204
rect 210516 132880 210568 132932
rect 213920 132880 213972 132932
rect 300216 132608 300268 132660
rect 306932 132608 306984 132660
rect 297364 132540 297416 132592
rect 307300 132540 307352 132592
rect 171968 132472 172020 132524
rect 213920 132472 213972 132524
rect 292028 132472 292080 132524
rect 306564 132472 306616 132524
rect 252284 132404 252336 132456
rect 297456 132404 297508 132456
rect 367744 132404 367796 132456
rect 417516 132404 417568 132456
rect 252468 132336 252520 132388
rect 278228 132336 278280 132388
rect 252376 132268 252428 132320
rect 264336 132268 264388 132320
rect 294604 131248 294656 131300
rect 307484 131248 307536 131300
rect 290556 131180 290608 131232
rect 307576 131180 307628 131232
rect 202328 131112 202380 131164
rect 213920 131112 213972 131164
rect 278136 131112 278188 131164
rect 307668 131112 307720 131164
rect 497464 131112 497516 131164
rect 498292 131112 498344 131164
rect 252468 131044 252520 131096
rect 267188 131044 267240 131096
rect 324412 131044 324464 131096
rect 346492 131044 346544 131096
rect 252376 130976 252428 131028
rect 261668 130976 261720 131028
rect 324320 130976 324372 131028
rect 331312 130976 331364 131028
rect 252468 130160 252520 130212
rect 259000 130160 259052 130212
rect 301504 129888 301556 129940
rect 307484 129888 307536 129940
rect 176016 129820 176068 129872
rect 213920 129820 213972 129872
rect 304448 129820 304500 129872
rect 306932 129820 306984 129872
rect 173348 129752 173400 129804
rect 214012 129752 214064 129804
rect 261576 129752 261628 129804
rect 306564 129752 306616 129804
rect 252284 129684 252336 129736
rect 300308 129684 300360 129736
rect 324320 129684 324372 129736
rect 349344 129684 349396 129736
rect 496820 129684 496872 129736
rect 509240 129684 509292 129736
rect 252468 129616 252520 129668
rect 291936 129616 291988 129668
rect 252376 129548 252428 129600
rect 264428 129548 264480 129600
rect 298836 128460 298888 128512
rect 307668 128460 307720 128512
rect 284944 128392 284996 128444
rect 306932 128392 306984 128444
rect 177488 128324 177540 128376
rect 213920 128324 213972 128376
rect 264336 128324 264388 128376
rect 307576 128324 307628 128376
rect 252376 128256 252428 128308
rect 271144 128256 271196 128308
rect 324320 128256 324372 128308
rect 350632 128256 350684 128308
rect 382924 128256 382976 128308
rect 418712 128256 418764 128308
rect 496820 128256 496872 128308
rect 507860 128256 507912 128308
rect 252468 128188 252520 128240
rect 268384 128188 268436 128240
rect 324412 128188 324464 128240
rect 329932 128188 329984 128240
rect 252284 128120 252336 128172
rect 257620 128120 257672 128172
rect 268568 127644 268620 127696
rect 307392 127644 307444 127696
rect 252192 127576 252244 127628
rect 305644 127576 305696 127628
rect 530584 127576 530636 127628
rect 580172 127576 580224 127628
rect 496912 127236 496964 127288
rect 499856 127236 499908 127288
rect 184388 127032 184440 127084
rect 214012 127032 214064 127084
rect 295984 127032 296036 127084
rect 307576 127032 307628 127084
rect 57796 126964 57848 127016
rect 65524 126964 65576 127016
rect 173256 126964 173308 127016
rect 213920 126964 213972 127016
rect 293224 126964 293276 127016
rect 307668 126964 307720 127016
rect 252468 126896 252520 126948
rect 272524 126896 272576 126948
rect 496820 126896 496872 126948
rect 514760 126896 514812 126948
rect 251180 126828 251232 126880
rect 253388 126828 253440 126880
rect 252468 126420 252520 126472
rect 258724 126420 258776 126472
rect 252284 126216 252336 126268
rect 293316 126216 293368 126268
rect 296168 125740 296220 125792
rect 307668 125740 307720 125792
rect 192484 125672 192536 125724
rect 214012 125672 214064 125724
rect 283564 125672 283616 125724
rect 307484 125672 307536 125724
rect 169116 125604 169168 125656
rect 213920 125604 213972 125656
rect 275284 125604 275336 125656
rect 307576 125604 307628 125656
rect 252100 125536 252152 125588
rect 253572 125536 253624 125588
rect 324412 125536 324464 125588
rect 346400 125536 346452 125588
rect 496820 125536 496872 125588
rect 513380 125536 513432 125588
rect 252468 125468 252520 125520
rect 269856 125468 269908 125520
rect 324320 125468 324372 125520
rect 327724 125468 327776 125520
rect 252376 125400 252428 125452
rect 301596 125400 301648 125452
rect 301688 124312 301740 124364
rect 307668 124312 307720 124364
rect 180340 124244 180392 124296
rect 213920 124244 213972 124296
rect 285036 124244 285088 124296
rect 307576 124244 307628 124296
rect 171876 124176 171928 124228
rect 214012 124176 214064 124228
rect 272524 124176 272576 124228
rect 307484 124176 307536 124228
rect 252468 124108 252520 124160
rect 302976 124108 303028 124160
rect 324412 124108 324464 124160
rect 349252 124108 349304 124160
rect 324320 124040 324372 124092
rect 347780 124040 347832 124092
rect 496820 124040 496872 124092
rect 499580 124040 499632 124092
rect 251732 123428 251784 123480
rect 264520 123428 264572 123480
rect 293316 122952 293368 123004
rect 307576 122952 307628 123004
rect 196808 122884 196860 122936
rect 213920 122884 213972 122936
rect 56508 122816 56560 122868
rect 66076 122816 66128 122868
rect 170496 122816 170548 122868
rect 214012 122816 214064 122868
rect 303068 122816 303120 122868
rect 307668 122816 307720 122868
rect 252468 122748 252520 122800
rect 299020 122748 299072 122800
rect 324320 122748 324372 122800
rect 347964 122748 348016 122800
rect 376668 122748 376720 122800
rect 416780 122748 416832 122800
rect 496820 122748 496872 122800
rect 505100 122748 505152 122800
rect 252376 122680 252428 122732
rect 269948 122680 270000 122732
rect 324412 122680 324464 122732
rect 342260 122680 342312 122732
rect 252284 122612 252336 122664
rect 262864 122612 262916 122664
rect 279424 122068 279476 122120
rect 308496 122068 308548 122120
rect 298744 121592 298796 121644
rect 307668 121592 307720 121644
rect 203524 121524 203576 121576
rect 214012 121524 214064 121576
rect 297456 121524 297508 121576
rect 307484 121524 307536 121576
rect 166448 121456 166500 121508
rect 213920 121456 213972 121508
rect 269856 121456 269908 121508
rect 307576 121456 307628 121508
rect 252468 121388 252520 121440
rect 287980 121388 288032 121440
rect 324320 121388 324372 121440
rect 335360 121388 335412 121440
rect 407764 121388 407816 121440
rect 416780 121388 416832 121440
rect 252468 120300 252520 120352
rect 260472 120300 260524 120352
rect 287888 120232 287940 120284
rect 307668 120232 307720 120284
rect 183008 120164 183060 120216
rect 214012 120164 214064 120216
rect 268384 120164 268436 120216
rect 307484 120164 307536 120216
rect 57888 120096 57940 120148
rect 65156 120096 65208 120148
rect 169024 120096 169076 120148
rect 213920 120096 213972 120148
rect 260104 120096 260156 120148
rect 307576 120096 307628 120148
rect 252468 120028 252520 120080
rect 273904 120028 273956 120080
rect 324320 119960 324372 120012
rect 325976 119960 326028 120012
rect 496912 119552 496964 119604
rect 500960 119552 501012 119604
rect 263048 119416 263100 119468
rect 307116 119416 307168 119468
rect 251916 119348 251968 119400
rect 304356 119348 304408 119400
rect 252468 118940 252520 118992
rect 260380 118940 260432 118992
rect 170588 118804 170640 118856
rect 214012 118804 214064 118856
rect 278320 118804 278372 118856
rect 307668 118804 307720 118856
rect 178868 118736 178920 118788
rect 213920 118736 213972 118788
rect 300308 118668 300360 118720
rect 307484 118668 307536 118720
rect 252468 118600 252520 118652
rect 290464 118600 290516 118652
rect 324412 118600 324464 118652
rect 345112 118600 345164 118652
rect 371884 118600 371936 118652
rect 416780 118600 416832 118652
rect 496820 118600 496872 118652
rect 517520 118600 517572 118652
rect 252376 118532 252428 118584
rect 257344 118532 257396 118584
rect 324320 118532 324372 118584
rect 342352 118532 342404 118584
rect 252100 117920 252152 117972
rect 275376 117920 275428 117972
rect 304540 117444 304592 117496
rect 307576 117444 307628 117496
rect 203616 117376 203668 117428
rect 213920 117376 213972 117428
rect 282368 117376 282420 117428
rect 306564 117376 306616 117428
rect 173440 117308 173492 117360
rect 214012 117308 214064 117360
rect 261668 117308 261720 117360
rect 307668 117308 307720 117360
rect 252376 117240 252428 117292
rect 277032 117240 277084 117292
rect 340236 117240 340288 117292
rect 416780 117240 416832 117292
rect 496820 117240 496872 117292
rect 503812 117240 503864 117292
rect 252284 117172 252336 117224
rect 267004 117172 267056 117224
rect 324412 117172 324464 117224
rect 338120 117172 338172 117224
rect 324320 117104 324372 117156
rect 340972 117104 341024 117156
rect 252468 116832 252520 116884
rect 260288 116832 260340 116884
rect 276848 116084 276900 116136
rect 306748 116084 306800 116136
rect 207848 116016 207900 116068
rect 213920 116016 213972 116068
rect 273904 116016 273956 116068
rect 307668 116016 307720 116068
rect 181628 115948 181680 116000
rect 214012 115948 214064 116000
rect 258724 115948 258776 116000
rect 307576 115948 307628 116000
rect 252468 115880 252520 115932
rect 281080 115880 281132 115932
rect 324412 115880 324464 115932
rect 343732 115880 343784 115932
rect 252376 115812 252428 115864
rect 271236 115812 271288 115864
rect 324320 115812 324372 115864
rect 332692 115812 332744 115864
rect 290464 114656 290516 114708
rect 307668 114656 307720 114708
rect 280896 114588 280948 114640
rect 307576 114588 307628 114640
rect 195520 114520 195572 114572
rect 213920 114520 213972 114572
rect 252376 114520 252428 114572
rect 258908 114520 258960 114572
rect 271144 114520 271196 114572
rect 307484 114520 307536 114572
rect 252468 114452 252520 114504
rect 261760 114452 261812 114504
rect 324412 114452 324464 114504
rect 345020 114452 345072 114504
rect 385684 114452 385736 114504
rect 416780 114452 416832 114504
rect 324320 114384 324372 114436
rect 341156 114384 341208 114436
rect 496820 114180 496872 114232
rect 499672 114180 499724 114232
rect 252468 113772 252520 113824
rect 268476 113772 268528 113824
rect 291936 113296 291988 113348
rect 307668 113296 307720 113348
rect 200948 113228 201000 113280
rect 214012 113228 214064 113280
rect 265716 113228 265768 113280
rect 307576 113228 307628 113280
rect 196900 113160 196952 113212
rect 213920 113160 213972 113212
rect 249064 113160 249116 113212
rect 307668 113160 307720 113212
rect 324320 113092 324372 113144
rect 349160 113092 349212 113144
rect 252468 112888 252520 112940
rect 255964 112888 256016 112940
rect 413284 112888 413336 112940
rect 416780 112888 416832 112940
rect 252100 112480 252152 112532
rect 289268 112480 289320 112532
rect 252192 112412 252244 112464
rect 304264 112412 304316 112464
rect 205180 111868 205232 111920
rect 213920 111868 213972 111920
rect 252468 111868 252520 111920
rect 258816 111868 258868 111920
rect 304356 111868 304408 111920
rect 307668 111868 307720 111920
rect 174728 111800 174780 111852
rect 214012 111800 214064 111852
rect 267004 111800 267056 111852
rect 306932 111800 306984 111852
rect 3424 111732 3476 111784
rect 11704 111732 11756 111784
rect 167920 111732 167972 111784
rect 205088 111732 205140 111784
rect 252468 111732 252520 111784
rect 296076 111732 296128 111784
rect 324320 111732 324372 111784
rect 336832 111732 336884 111784
rect 388444 111732 388496 111784
rect 416780 111732 416832 111784
rect 496820 111732 496872 111784
rect 506480 111732 506532 111784
rect 252284 111664 252336 111716
rect 254584 111664 254636 111716
rect 324412 111664 324464 111716
rect 336740 111664 336792 111716
rect 496820 111596 496872 111648
rect 501144 111596 501196 111648
rect 294788 110576 294840 110628
rect 307484 110576 307536 110628
rect 176200 110508 176252 110560
rect 213920 110508 213972 110560
rect 273996 110508 274048 110560
rect 307576 110508 307628 110560
rect 166540 110440 166592 110492
rect 214012 110440 214064 110492
rect 253388 110440 253440 110492
rect 307668 110440 307720 110492
rect 252284 110372 252336 110424
rect 305828 110372 305880 110424
rect 324320 110372 324372 110424
rect 341064 110372 341116 110424
rect 377404 110372 377456 110424
rect 416780 110372 416832 110424
rect 496820 110372 496872 110424
rect 510620 110372 510672 110424
rect 252376 110304 252428 110356
rect 298928 110304 298980 110356
rect 252468 110236 252520 110288
rect 279516 110236 279568 110288
rect 324412 109692 324464 109744
rect 328460 109692 328512 109744
rect 174820 109080 174872 109132
rect 213920 109080 213972 109132
rect 302884 109080 302936 109132
rect 306932 109080 306984 109132
rect 167828 109012 167880 109064
rect 214012 109012 214064 109064
rect 289268 109012 289320 109064
rect 307668 109012 307720 109064
rect 168104 108944 168156 108996
rect 180248 108944 180300 108996
rect 252468 108944 252520 108996
rect 283656 108944 283708 108996
rect 251732 108876 251784 108928
rect 254860 108876 254912 108928
rect 251824 108332 251876 108384
rect 256240 108332 256292 108384
rect 324320 108196 324372 108248
rect 327172 108196 327224 108248
rect 255964 107856 256016 107908
rect 307668 107856 307720 107908
rect 180432 107720 180484 107772
rect 214012 107720 214064 107772
rect 279424 107720 279476 107772
rect 307668 107720 307720 107772
rect 169208 107652 169260 107704
rect 213920 107652 213972 107704
rect 302976 107652 303028 107704
rect 307576 107652 307628 107704
rect 252468 107584 252520 107636
rect 265624 107584 265676 107636
rect 324320 107584 324372 107636
rect 354680 107584 354732 107636
rect 389824 107584 389876 107636
rect 416780 107584 416832 107636
rect 496820 107584 496872 107636
rect 502340 107584 502392 107636
rect 251732 107516 251784 107568
rect 254768 107516 254820 107568
rect 304264 106428 304316 106480
rect 307576 106428 307628 106480
rect 176108 106360 176160 106412
rect 214012 106360 214064 106412
rect 254584 106360 254636 106412
rect 307484 106360 307536 106412
rect 170680 106292 170732 106344
rect 213920 106292 213972 106344
rect 250720 106292 250772 106344
rect 307668 106292 307720 106344
rect 252376 106224 252428 106276
rect 285128 106224 285180 106276
rect 342904 106224 342956 106276
rect 416780 106224 416832 106276
rect 252468 106156 252520 106208
rect 265808 106156 265860 106208
rect 252284 106088 252336 106140
rect 257528 106088 257580 106140
rect 283656 105000 283708 105052
rect 307484 105000 307536 105052
rect 192576 104932 192628 104984
rect 213920 104932 213972 104984
rect 265624 104932 265676 104984
rect 307668 104932 307720 104984
rect 172060 104864 172112 104916
rect 214012 104864 214064 104916
rect 257344 104864 257396 104916
rect 306932 104864 306984 104916
rect 252376 104796 252428 104848
rect 276940 104796 276992 104848
rect 356704 104796 356756 104848
rect 416780 104796 416832 104848
rect 252468 104728 252520 104780
rect 272616 104728 272668 104780
rect 252284 104660 252336 104712
rect 256148 104660 256200 104712
rect 325700 104116 325752 104168
rect 354036 104116 354088 104168
rect 276756 103640 276808 103692
rect 306932 103640 306984 103692
rect 275376 103572 275428 103624
rect 307668 103572 307720 103624
rect 199476 103504 199528 103556
rect 213920 103504 213972 103556
rect 267188 103504 267240 103556
rect 307576 103504 307628 103556
rect 252468 103436 252520 103488
rect 303160 103436 303212 103488
rect 393964 103436 394016 103488
rect 416780 103436 416832 103488
rect 252376 103028 252428 103080
rect 256056 103028 256108 103080
rect 252468 102892 252520 102944
rect 260196 102892 260248 102944
rect 323584 102756 323636 102808
rect 367836 102756 367888 102808
rect 297548 102212 297600 102264
rect 307668 102212 307720 102264
rect 211988 102144 212040 102196
rect 213920 102144 213972 102196
rect 258908 102144 258960 102196
rect 307576 102144 307628 102196
rect 252468 102076 252520 102128
rect 269764 102076 269816 102128
rect 324320 102076 324372 102128
rect 332968 102076 333020 102128
rect 396724 102076 396776 102128
rect 416780 102076 416832 102128
rect 251364 102008 251416 102060
rect 253296 102008 253348 102060
rect 252192 101396 252244 101448
rect 267096 101396 267148 101448
rect 301596 100920 301648 100972
rect 306564 100920 306616 100972
rect 285128 100852 285180 100904
rect 307668 100852 307720 100904
rect 207756 100784 207808 100836
rect 214012 100784 214064 100836
rect 269948 100784 270000 100836
rect 307576 100784 307628 100836
rect 66168 100716 66220 100768
rect 68284 100716 68336 100768
rect 205088 100716 205140 100768
rect 213920 100716 213972 100768
rect 264428 100716 264480 100768
rect 306932 100716 306984 100768
rect 252376 100648 252428 100700
rect 286508 100648 286560 100700
rect 378784 100648 378836 100700
rect 493968 100648 494020 100700
rect 520188 100648 520240 100700
rect 580172 100648 580224 100700
rect 252284 100580 252336 100632
rect 268568 100580 268620 100632
rect 395344 100580 395396 100632
rect 494244 100580 494296 100632
rect 252468 100512 252520 100564
rect 263048 100512 263100 100564
rect 330484 99968 330536 100020
rect 370504 99968 370556 100020
rect 296076 99492 296128 99544
rect 306564 99492 306616 99544
rect 272616 99424 272668 99476
rect 307668 99424 307720 99476
rect 167736 99356 167788 99408
rect 213920 99356 213972 99408
rect 262864 99356 262916 99408
rect 307576 99356 307628 99408
rect 252468 99288 252520 99340
rect 261484 99288 261536 99340
rect 324320 99288 324372 99340
rect 339500 99288 339552 99340
rect 419632 99288 419684 99340
rect 580264 99288 580316 99340
rect 399484 99220 399536 99272
rect 496912 99220 496964 99272
rect 324412 98744 324464 98796
rect 324688 98744 324740 98796
rect 169300 98608 169352 98660
rect 214012 98608 214064 98660
rect 252468 98608 252520 98660
rect 262956 98608 263008 98660
rect 324412 98608 324464 98660
rect 331220 98608 331272 98660
rect 298928 98132 298980 98184
rect 306932 98132 306984 98184
rect 264520 98064 264572 98116
rect 307576 98064 307628 98116
rect 165252 97996 165304 98048
rect 213920 97996 213972 98048
rect 256056 97996 256108 98048
rect 307668 97996 307720 98048
rect 256700 97928 256752 97980
rect 257436 97928 257488 97980
rect 324320 97928 324372 97980
rect 350540 97928 350592 97980
rect 392584 97928 392636 97980
rect 495440 97928 495492 97980
rect 410524 97860 410576 97912
rect 497004 97860 497056 97912
rect 2780 97724 2832 97776
rect 4804 97724 4856 97776
rect 420184 97316 420236 97368
rect 427728 97316 427780 97368
rect 421564 97248 421616 97300
rect 458916 97248 458968 97300
rect 467104 97248 467156 97300
rect 492496 97248 492548 97300
rect 439504 96908 439556 96960
rect 440884 96908 440936 96960
rect 454040 96908 454092 96960
rect 455052 96908 455104 96960
rect 461584 96908 461636 96960
rect 464896 96908 464948 96960
rect 465724 96908 465776 96960
rect 467288 96908 467340 96960
rect 472624 96908 472676 96960
rect 474556 96908 474608 96960
rect 481640 96908 481692 96960
rect 482652 96908 482704 96960
rect 486424 96908 486476 96960
rect 487712 96908 487764 96960
rect 417424 96772 417476 96824
rect 420552 96772 420604 96824
rect 252468 96704 252520 96756
rect 256700 96704 256752 96756
rect 269764 96704 269816 96756
rect 307668 96704 307720 96756
rect 251824 96636 251876 96688
rect 307484 96636 307536 96688
rect 282276 96568 282328 96620
rect 321560 96568 321612 96620
rect 406384 96568 406436 96620
rect 496820 96568 496872 96620
rect 309784 96500 309836 96552
rect 322940 96500 322992 96552
rect 308404 96432 308456 96484
rect 321652 96432 321704 96484
rect 184296 95956 184348 96008
rect 222844 95956 222896 96008
rect 168288 95888 168340 95940
rect 214564 95888 214616 95940
rect 343640 95888 343692 95940
rect 498476 95888 498528 95940
rect 249248 95208 249300 95260
rect 307668 95208 307720 95260
rect 198188 95140 198240 95192
rect 321468 95140 321520 95192
rect 202236 95072 202288 95124
rect 321836 95072 321888 95124
rect 204904 95004 204956 95056
rect 321744 95004 321796 95056
rect 294696 94936 294748 94988
rect 324688 94936 324740 94988
rect 308496 94868 308548 94920
rect 324504 94868 324556 94920
rect 161480 94528 161532 94580
rect 207848 94528 207900 94580
rect 130384 94460 130436 94512
rect 214012 94460 214064 94512
rect 289084 94460 289136 94512
rect 324320 94460 324372 94512
rect 426532 94460 426584 94512
rect 125416 93984 125468 94036
rect 169116 93984 169168 94036
rect 112352 93916 112404 93968
rect 178868 93916 178920 93968
rect 85580 93848 85632 93900
rect 165252 93848 165304 93900
rect 67364 93780 67416 93832
rect 214840 93780 214892 93832
rect 278044 93780 278096 93832
rect 323584 93780 323636 93832
rect 198924 93712 198976 93764
rect 324596 93712 324648 93764
rect 151728 93372 151780 93424
rect 173164 93372 173216 93424
rect 118240 93304 118292 93356
rect 166448 93304 166500 93356
rect 133144 93236 133196 93288
rect 200856 93236 200908 93288
rect 129464 93168 129516 93220
rect 198096 93168 198148 93220
rect 320824 93168 320876 93220
rect 420184 93168 420236 93220
rect 98552 93100 98604 93152
rect 176200 93100 176252 93152
rect 182916 93100 182968 93152
rect 262956 93100 263008 93152
rect 419264 93100 419316 93152
rect 580264 93100 580316 93152
rect 322940 93032 322992 93084
rect 323584 93032 323636 93084
rect 110144 92420 110196 92472
rect 203616 92420 203668 92472
rect 216128 92420 216180 92472
rect 497096 92420 497148 92472
rect 120356 92352 120408 92404
rect 211896 92352 211948 92404
rect 115480 92284 115532 92336
rect 202420 92284 202472 92336
rect 88984 92216 89036 92268
rect 169300 92216 169352 92268
rect 86776 92148 86828 92200
rect 130384 92148 130436 92200
rect 130752 92148 130804 92200
rect 174636 92148 174688 92200
rect 136088 92080 136140 92132
rect 168288 92080 168340 92132
rect 85120 91060 85172 91112
rect 120724 91060 120776 91112
rect 56508 90992 56560 91044
rect 211988 90992 212040 91044
rect 114376 90924 114428 90976
rect 196716 90924 196768 90976
rect 107752 90856 107804 90908
rect 161480 90856 161532 90908
rect 122104 90788 122156 90840
rect 170496 90788 170548 90840
rect 151636 90720 151688 90772
rect 199384 90720 199436 90772
rect 135168 90652 135220 90704
rect 171784 90652 171836 90704
rect 189816 90312 189868 90364
rect 321560 90312 321612 90364
rect 465080 90312 465132 90364
rect 90548 89632 90600 89684
rect 172060 89632 172112 89684
rect 249156 89632 249208 89684
rect 256700 89632 256752 89684
rect 420920 89632 420972 89684
rect 95056 89564 95108 89616
rect 169208 89564 169260 89616
rect 103336 89496 103388 89548
rect 173348 89496 173400 89548
rect 126520 89428 126572 89480
rect 192484 89428 192536 89480
rect 122840 89360 122892 89412
rect 180340 89360 180392 89412
rect 153016 89292 153068 89344
rect 206376 89292 206428 89344
rect 280804 89020 280856 89072
rect 311900 89020 311952 89072
rect 352656 89020 352708 89072
rect 171784 88952 171836 89004
rect 307300 88952 307352 89004
rect 352564 88952 352616 89004
rect 462320 88952 462372 89004
rect 100576 88272 100628 88324
rect 205180 88272 205232 88324
rect 104440 88204 104492 88256
rect 200948 88204 201000 88256
rect 124772 88136 124824 88188
rect 204996 88136 205048 88188
rect 107292 88068 107344 88120
rect 171968 88068 172020 88120
rect 151452 88000 151504 88052
rect 213368 88000 213420 88052
rect 114928 87932 114980 87984
rect 170588 87932 170640 87984
rect 175924 87660 175976 87712
rect 257436 87660 257488 87712
rect 242164 87592 242216 87644
rect 347044 87592 347096 87644
rect 354036 87592 354088 87644
rect 456800 87592 456852 87644
rect 75368 86912 75420 86964
rect 214748 86912 214800 86964
rect 358176 86912 358228 86964
rect 421564 86912 421616 86964
rect 504364 86912 504416 86964
rect 580172 86912 580224 86964
rect 105544 86844 105596 86896
rect 216680 86844 216732 86896
rect 106096 86776 106148 86828
rect 202328 86776 202380 86828
rect 100208 86708 100260 86760
rect 166540 86708 166592 86760
rect 123300 86640 123352 86692
rect 178776 86640 178828 86692
rect 115848 86572 115900 86624
rect 169024 86572 169076 86624
rect 342260 86368 342312 86420
rect 357532 86368 357584 86420
rect 358176 86368 358228 86420
rect 177304 86300 177356 86352
rect 253296 86300 253348 86352
rect 308404 86300 308456 86352
rect 345664 86300 345716 86352
rect 209136 86232 209188 86284
rect 244280 86232 244332 86284
rect 342996 86232 343048 86284
rect 377404 86232 377456 86284
rect 455420 86232 455472 86284
rect 3148 85484 3200 85536
rect 32404 85484 32456 85536
rect 88064 85484 88116 85536
rect 167736 85484 167788 85536
rect 127624 85416 127676 85468
rect 206468 85416 206520 85468
rect 120632 85348 120684 85400
rect 196808 85348 196860 85400
rect 101864 85280 101916 85332
rect 174728 85280 174780 85332
rect 111248 85212 111300 85264
rect 173440 85212 173492 85264
rect 195336 84872 195388 84924
rect 266360 84872 266412 84924
rect 195428 84804 195480 84856
rect 307208 84804 307260 84856
rect 316040 84804 316092 84856
rect 333244 84804 333296 84856
rect 336096 84804 336148 84856
rect 460940 84804 460992 84856
rect 65984 84124 66036 84176
rect 214656 84124 214708 84176
rect 291844 84124 291896 84176
rect 332048 84124 332100 84176
rect 103428 84056 103480 84108
rect 196900 84056 196952 84108
rect 96528 83988 96580 84040
rect 174820 83988 174872 84040
rect 92388 83920 92440 83972
rect 170680 83920 170732 83972
rect 117136 83852 117188 83904
rect 181536 83852 181588 83904
rect 132408 83784 132460 83836
rect 166264 83784 166316 83836
rect 185676 83444 185728 83496
rect 254768 83444 254820 83496
rect 331956 83444 332008 83496
rect 463700 83444 463752 83496
rect 291200 82832 291252 82884
rect 291844 82832 291896 82884
rect 108948 82764 109000 82816
rect 210516 82764 210568 82816
rect 107568 82696 107620 82748
rect 195520 82696 195572 82748
rect 101956 82628 102008 82680
rect 176016 82628 176068 82680
rect 117228 82560 117280 82612
rect 183008 82560 183060 82612
rect 119896 82492 119948 82544
rect 170404 82492 170456 82544
rect 122748 82424 122800 82476
rect 166356 82424 166408 82476
rect 238024 82084 238076 82136
rect 251180 82084 251232 82136
rect 324964 82084 325016 82136
rect 461584 82084 461636 82136
rect 99196 81336 99248 81388
rect 184388 81336 184440 81388
rect 345756 81336 345808 81388
rect 465724 81336 465776 81388
rect 119988 81268 120040 81320
rect 203524 81268 203576 81320
rect 110236 81200 110288 81252
rect 181628 81200 181680 81252
rect 97816 81132 97868 81184
rect 167828 81132 167880 81184
rect 184204 80656 184256 80708
rect 313924 80656 313976 80708
rect 317420 80044 317472 80096
rect 345756 80044 345808 80096
rect 68284 79976 68336 80028
rect 199476 79976 199528 80028
rect 93768 79908 93820 79960
rect 176108 79908 176160 79960
rect 126888 79840 126940 79892
rect 209228 79840 209280 79892
rect 102048 79772 102100 79824
rect 177488 79772 177540 79824
rect 97908 79704 97960 79756
rect 173256 79704 173308 79756
rect 195244 79364 195296 79416
rect 232504 79364 232556 79416
rect 200764 79296 200816 79348
rect 246304 79296 246356 79348
rect 309784 79296 309836 79348
rect 470600 79296 470652 79348
rect 114468 78616 114520 78668
rect 213460 78616 213512 78668
rect 266360 78616 266412 78668
rect 338764 78616 338816 78668
rect 339132 78616 339184 78668
rect 471980 78616 472032 78668
rect 95148 78548 95200 78600
rect 180432 78548 180484 78600
rect 110328 78480 110380 78532
rect 177396 78480 177448 78532
rect 188436 78004 188488 78056
rect 286508 78004 286560 78056
rect 42708 77936 42760 77988
rect 128360 77936 128412 77988
rect 180156 77936 180208 77988
rect 278228 77936 278280 77988
rect 120724 77188 120776 77240
rect 205088 77188 205140 77240
rect 123944 77120 123996 77172
rect 171876 77120 171928 77172
rect 102140 76508 102192 76560
rect 305920 76508 305972 76560
rect 307208 76508 307260 76560
rect 473360 76508 473412 76560
rect 93860 75216 93912 75268
rect 297456 75216 297508 75268
rect 53840 75148 53892 75200
rect 267188 75148 267240 75200
rect 297640 75148 297692 75200
rect 472624 75148 472676 75200
rect 57888 74468 57940 74520
rect 207756 74468 207808 74520
rect 86960 73856 87012 73908
rect 269856 73856 269908 73908
rect 121460 73788 121512 73840
rect 309140 73788 309192 73840
rect 311164 73788 311216 73840
rect 469220 73788 469272 73840
rect 64604 73108 64656 73160
rect 320824 73108 320876 73160
rect 419448 73108 419500 73160
rect 579988 73108 580040 73160
rect 262956 73040 263008 73092
rect 414664 73040 414716 73092
rect 107660 72496 107712 72548
rect 253388 72496 253440 72548
rect 60740 72428 60792 72480
rect 290556 72428 290608 72480
rect 262220 71748 262272 71800
rect 262956 71748 263008 71800
rect 320180 71748 320232 71800
rect 320824 71748 320876 71800
rect 3424 71680 3476 71732
rect 41328 71680 41380 71732
rect 494152 71680 494204 71732
rect 80060 71068 80112 71120
rect 287888 71068 287940 71120
rect 66260 71000 66312 71052
rect 278320 71000 278372 71052
rect 362960 70320 363012 70372
rect 459560 70320 459612 70372
rect 178684 69776 178736 69828
rect 347044 69776 347096 69828
rect 54760 69708 54812 69760
rect 226984 69708 227036 69760
rect 55220 69640 55272 69692
rect 304540 69640 304592 69692
rect 339500 69640 339552 69692
rect 362960 69640 363012 69692
rect 60648 68960 60700 69012
rect 335360 68960 335412 69012
rect 336096 68960 336148 69012
rect 104900 68348 104952 68400
rect 293316 68348 293368 68400
rect 52368 68280 52420 68332
rect 246396 68280 246448 68332
rect 286324 68280 286376 68332
rect 292580 68280 292632 68332
rect 474740 68280 474792 68332
rect 287704 67532 287756 67584
rect 289820 67532 289872 67584
rect 114560 66988 114612 67040
rect 294788 66988 294840 67040
rect 289820 66920 289872 66972
rect 476120 66920 476172 66972
rect 35900 66852 35952 66904
rect 298836 66852 298888 66904
rect 285680 66172 285732 66224
rect 286508 66172 286560 66224
rect 477500 66172 477552 66224
rect 193864 65628 193916 65680
rect 332048 65628 332100 65680
rect 61660 65560 61712 65612
rect 269856 65560 269908 65612
rect 40040 65492 40092 65544
rect 297548 65492 297600 65544
rect 188344 64268 188396 64320
rect 333244 64268 333296 64320
rect 59176 64200 59228 64252
rect 274088 64200 274140 64252
rect 276664 64200 276716 64252
rect 278780 64200 278832 64252
rect 480260 64200 480312 64252
rect 73160 64132 73212 64184
rect 300308 64132 300360 64184
rect 98000 62840 98052 62892
rect 303068 62840 303120 62892
rect 33140 62772 33192 62824
rect 269948 62772 270000 62824
rect 278044 62772 278096 62824
rect 481732 62772 481784 62824
rect 118700 61412 118752 61464
rect 272524 61412 272576 61464
rect 273168 61344 273220 61396
rect 481640 61344 481692 61396
rect 512644 60664 512696 60716
rect 580172 60664 580224 60716
rect 52460 60052 52512 60104
rect 261576 60052 261628 60104
rect 268476 60052 268528 60104
rect 483020 60052 483072 60104
rect 56600 59984 56652 60036
rect 278136 59984 278188 60036
rect 3056 59304 3108 59356
rect 17224 59304 17276 59356
rect 332600 59304 332652 59356
rect 400864 59304 400916 59356
rect 246396 58828 246448 58880
rect 264980 58828 265032 58880
rect 84200 58760 84252 58812
rect 268384 58760 268436 58812
rect 49700 58692 49752 58744
rect 304448 58692 304500 58744
rect 6920 58624 6972 58676
rect 264520 58624 264572 58676
rect 264980 58624 265032 58676
rect 484400 58624 484452 58676
rect 261484 57876 261536 57928
rect 485780 57876 485832 57928
rect 260840 57400 260892 57452
rect 261484 57400 261536 57452
rect 52552 57196 52604 57248
rect 261668 57196 261720 57248
rect 122840 55972 122892 56024
rect 296168 55972 296220 56024
rect 46940 55904 46992 55956
rect 258908 55904 258960 55956
rect 19340 55836 19392 55888
rect 256056 55836 256108 55888
rect 254768 55768 254820 55820
rect 488540 55836 488592 55888
rect 51080 54612 51132 54664
rect 275376 54612 275428 54664
rect 67640 54544 67692 54596
rect 297364 54544 297416 54596
rect 124220 54476 124272 54528
rect 250628 54476 250680 54528
rect 251916 54476 251968 54528
rect 489920 54476 489972 54528
rect 74540 53184 74592 53236
rect 292028 53184 292080 53236
rect 31760 53116 31812 53168
rect 264336 53116 264388 53168
rect 37188 53048 37240 53100
rect 232596 53048 232648 53100
rect 247960 53048 248012 53100
rect 491300 53048 491352 53100
rect 243544 51824 243596 51876
rect 467104 51824 467156 51876
rect 70400 51756 70452 51808
rect 300216 51756 300268 51808
rect 4160 51688 4212 51740
rect 249248 51688 249300 51740
rect 196624 51008 196676 51060
rect 247040 51008 247092 51060
rect 247960 51008 248012 51060
rect 71780 50464 71832 50516
rect 250720 50464 250772 50516
rect 240784 50396 240836 50448
rect 492680 50396 492732 50448
rect 24860 50328 24912 50380
rect 298928 50328 298980 50380
rect 64696 49648 64748 49700
rect 310520 49648 310572 49700
rect 311164 49648 311216 49700
rect 349160 49648 349212 49700
rect 352012 49648 352064 49700
rect 494060 49648 494112 49700
rect 269120 49580 269172 49632
rect 269856 49580 269908 49632
rect 359464 49580 359516 49632
rect 88340 49036 88392 49088
rect 289176 49036 289228 49088
rect 37280 48968 37332 49020
rect 271144 48968 271196 49020
rect 274088 48220 274140 48272
rect 340144 48220 340196 48272
rect 189724 47676 189776 47728
rect 315304 47676 315356 47728
rect 99380 47608 99432 47660
rect 254676 47608 254728 47660
rect 110420 47540 110472 47592
rect 273996 47540 274048 47592
rect 340880 47540 340932 47592
rect 498200 47540 498252 47592
rect 273260 47336 273312 47388
rect 274088 47336 274140 47388
rect 367836 46860 367888 46912
rect 422300 46860 422352 46912
rect 525064 46860 525116 46912
rect 580172 46860 580224 46912
rect 115940 46316 115992 46368
rect 285036 46316 285088 46368
rect 15200 46248 15252 46300
rect 251824 46248 251876 46300
rect 62028 46180 62080 46232
rect 327724 46180 327776 46232
rect 338120 46180 338172 46232
rect 367100 46180 367152 46232
rect 367836 46180 367888 46232
rect 3424 45500 3476 45552
rect 14464 45500 14516 45552
rect 182824 45500 182876 45552
rect 296720 45500 296772 45552
rect 297640 45500 297692 45552
rect 48320 44820 48372 44872
rect 258724 44820 258776 44872
rect 298836 44820 298888 44872
rect 360844 44820 360896 44872
rect 113180 43460 113232 43512
rect 250536 43460 250588 43512
rect 89720 43392 89772 43444
rect 305828 43392 305880 43444
rect 317328 43392 317380 43444
rect 427820 43392 427872 43444
rect 313280 42712 313332 42764
rect 313924 42712 313976 42764
rect 429200 42712 429252 42764
rect 35992 42032 36044 42084
rect 285128 42032 285180 42084
rect 342352 41352 342404 41404
rect 430580 41352 430632 41404
rect 38568 40808 38620 40860
rect 132500 40808 132552 40860
rect 120080 40740 120132 40792
rect 253204 40740 253256 40792
rect 93952 40672 94004 40724
rect 302976 40672 303028 40724
rect 309140 40060 309192 40112
rect 342352 40060 342404 40112
rect 288348 39584 288400 39636
rect 336004 39584 336056 39636
rect 210424 39516 210476 39568
rect 302240 39516 302292 39568
rect 185584 39448 185636 39500
rect 300768 39448 300820 39500
rect 117320 39380 117372 39432
rect 287796 39380 287848 39432
rect 11152 39312 11204 39364
rect 272616 39312 272668 39364
rect 302240 39312 302292 39364
rect 433340 39312 433392 39364
rect 300768 38632 300820 38684
rect 307208 38632 307260 38684
rect 232504 38020 232556 38072
rect 299480 38020 299532 38072
rect 92480 37952 92532 38004
rect 300124 37952 300176 38004
rect 26240 37884 26292 37936
rect 264428 37884 264480 37936
rect 299480 37884 299532 37936
rect 434720 37884 434772 37936
rect 222844 37204 222896 37256
rect 287060 37204 287112 37256
rect 288348 37204 288400 37256
rect 211804 36592 211856 36644
rect 295340 36592 295392 36644
rect 2780 36524 2832 36576
rect 269764 36524 269816 36576
rect 436192 36524 436244 36576
rect 206284 35300 206336 35352
rect 293960 35300 294012 35352
rect 111800 35232 111852 35284
rect 301688 35232 301740 35284
rect 44088 35164 44140 35216
rect 264336 35164 264388 35216
rect 293960 35164 294012 35216
rect 436284 35164 436336 35216
rect 289084 34416 289136 34468
rect 437480 34416 437532 34468
rect 41420 33804 41472 33856
rect 273904 33804 273956 33856
rect 30380 33736 30432 33788
rect 290464 33736 290516 33788
rect 288440 33124 288492 33176
rect 289084 33124 289136 33176
rect 3516 33056 3568 33108
rect 21364 33056 21416 33108
rect 327724 33056 327776 33108
rect 425060 33056 425112 33108
rect 118792 32444 118844 32496
rect 304356 32444 304408 32496
rect 95240 32376 95292 32428
rect 280988 32376 281040 32428
rect 327080 31764 327132 31816
rect 327724 31764 327776 31816
rect 246304 31220 246356 31272
rect 284392 31220 284444 31272
rect 85580 31152 85632 31204
rect 255964 31152 256016 31204
rect 438860 31152 438912 31204
rect 100760 31084 100812 31136
rect 289268 31084 289320 31136
rect 19432 31016 19484 31068
rect 293224 31016 293276 31068
rect 277400 30268 277452 30320
rect 278228 30268 278280 30320
rect 441620 30268 441672 30320
rect 110512 29656 110564 29708
rect 250444 29656 250496 29708
rect 82820 29588 82872 29640
rect 279424 29588 279476 29640
rect 59268 28908 59320 28960
rect 298100 28908 298152 28960
rect 298836 28908 298888 28960
rect 213276 28296 213328 28348
rect 274640 28296 274692 28348
rect 443000 28296 443052 28348
rect 44180 28228 44232 28280
rect 276848 28228 276900 28280
rect 64512 27548 64564 27600
rect 307760 27548 307812 27600
rect 308404 27548 308456 27600
rect 198004 26936 198056 26988
rect 17960 26868 18012 26920
rect 265716 26868 265768 26920
rect 270500 26868 270552 26920
rect 444380 26868 444432 26920
rect 216036 25576 216088 25628
rect 271972 25576 272024 25628
rect 445852 25576 445904 25628
rect 20720 25508 20772 25560
rect 296076 25508 296128 25560
rect 264336 24760 264388 24812
rect 445944 24760 445996 24812
rect 96620 24216 96672 24268
rect 302884 24216 302936 24268
rect 63500 24148 63552 24200
rect 294604 24148 294656 24200
rect 2872 24080 2924 24132
rect 264244 24080 264296 24132
rect 263600 23468 263652 23520
rect 264336 23468 264388 23520
rect 77300 22856 77352 22908
rect 260104 22856 260156 22908
rect 209044 22788 209096 22840
rect 259552 22788 259604 22840
rect 447140 22788 447192 22840
rect 9680 22720 9732 22772
rect 275284 22720 275336 22772
rect 253296 22040 253348 22092
rect 449900 22040 449952 22092
rect 252560 21564 252612 21616
rect 253296 21564 253348 21616
rect 69020 21496 69072 21548
rect 257344 21496 257396 21548
rect 91100 21428 91152 21480
rect 298744 21428 298796 21480
rect 67548 21360 67600 21412
rect 329104 21360 329156 21412
rect 331956 21360 332008 21412
rect 3424 20612 3476 20664
rect 22744 20612 22796 20664
rect 507124 20612 507176 20664
rect 579988 20612 580040 20664
rect 232596 20000 232648 20052
rect 249800 20000 249852 20052
rect 451280 20000 451332 20052
rect 22100 19932 22152 19984
rect 307116 19932 307168 19984
rect 20 19252 72 19304
rect 1308 19252 1360 19304
rect 249156 19252 249208 19304
rect 104164 18708 104216 18760
rect 307024 18708 307076 18760
rect 60832 18640 60884 18692
rect 265624 18640 265676 18692
rect 246304 18572 246356 18624
rect 452660 18572 452712 18624
rect 75920 17416 75972 17468
rect 254584 17416 254636 17468
rect 244924 17348 244976 17400
rect 454132 17348 454184 17400
rect 69112 17280 69164 17332
rect 305736 17280 305788 17332
rect 13820 17212 13872 17264
rect 283564 17212 283616 17264
rect 282276 15988 282328 16040
rect 454040 15988 454092 16040
rect 85672 15920 85724 15972
rect 286416 15920 286468 15972
rect 79232 15852 79284 15904
rect 304264 15852 304316 15904
rect 337016 15104 337068 15156
rect 501052 15104 501104 15156
rect 39120 14560 39172 14612
rect 284944 14560 284996 14612
rect 17040 14492 17092 14544
rect 262864 14492 262916 14544
rect 164424 14424 164476 14476
rect 417424 14424 417476 14476
rect 314660 13744 314712 13796
rect 315304 13744 315356 13796
rect 467840 13744 467892 13796
rect 249248 13676 249300 13728
rect 358084 13676 358136 13728
rect 58440 13064 58492 13116
rect 276756 13064 276808 13116
rect 248420 12452 248472 12504
rect 249248 12452 249300 12504
rect 202144 11772 202196 11824
rect 255872 11772 255924 11824
rect 353944 11772 353996 11824
rect 34520 11704 34572 11756
rect 280896 11704 280948 11756
rect 283564 11704 283616 11756
rect 478880 11704 478932 11756
rect 63040 10344 63092 10396
rect 282368 10344 282420 10396
rect 305552 10344 305604 10396
rect 331864 10344 331916 10396
rect 226984 10276 227036 10328
rect 258264 10276 258316 10328
rect 486424 10276 486476 10328
rect 186964 9596 187016 9648
rect 324964 9596 325016 9648
rect 325608 9596 325660 9648
rect 369860 9596 369912 9648
rect 499764 9596 499816 9648
rect 332048 9528 332100 9580
rect 423680 9528 423732 9580
rect 331588 9256 331640 9308
rect 332048 9256 332100 9308
rect 3424 8984 3476 9036
rect 29644 8984 29696 9036
rect 65524 8984 65576 9036
rect 283656 8984 283708 9036
rect 13544 8916 13596 8968
rect 249064 8916 249116 8968
rect 319720 8916 319772 8968
rect 334624 8916 334676 8968
rect 340972 8916 341024 8968
rect 369860 8916 369912 8968
rect 181444 8236 181496 8288
rect 283564 8236 283616 8288
rect 339960 8236 340012 8288
rect 431960 8236 432012 8288
rect 280804 8168 280856 8220
rect 344284 8168 344336 8220
rect 215944 7624 215996 7676
rect 301780 7624 301832 7676
rect 8760 7556 8812 7608
rect 267004 7556 267056 7608
rect 306748 6876 306800 6928
rect 339960 6876 340012 6928
rect 174544 6808 174596 6860
rect 242164 6808 242216 6860
rect 281908 6808 281960 6860
rect 439504 6808 439556 6860
rect 543004 6808 543056 6860
rect 580172 6808 580224 6860
rect 301780 6740 301832 6792
rect 363604 6740 363656 6792
rect 308496 6672 308548 6724
rect 309876 6672 309928 6724
rect 35808 6264 35860 6316
rect 136456 6264 136508 6316
rect 104532 6196 104584 6248
rect 305644 6196 305696 6248
rect 28908 6128 28960 6180
rect 295984 6128 296036 6180
rect 63132 5448 63184 5500
rect 251180 5448 251232 5500
rect 257068 5448 257120 5500
rect 257436 5448 257488 5500
rect 448520 5448 448572 5500
rect 251180 4972 251232 5024
rect 251916 4972 251968 5024
rect 180064 4904 180116 4956
rect 239220 4904 239272 4956
rect 213184 4836 213236 4888
rect 294880 4836 294932 4888
rect 27712 4768 27764 4820
rect 291936 4768 291988 4820
rect 356796 4768 356848 4820
rect 191104 4088 191156 4140
rect 246396 4088 246448 4140
rect 300768 4088 300820 4140
rect 307208 4088 307260 4140
rect 332692 4088 332744 4140
rect 333244 4088 333296 4140
rect 352564 4088 352616 4140
rect 239220 4020 239272 4072
rect 282276 4020 282328 4072
rect 349804 4020 349856 4072
rect 350448 4020 350500 4072
rect 377404 4020 377456 4072
rect 347044 3952 347096 4004
rect 354036 3952 354088 4004
rect 351184 3884 351236 3936
rect 351644 3884 351696 3936
rect 495532 3884 495584 3936
rect 125876 3680 125928 3732
rect 164884 3680 164936 3732
rect 78588 3612 78640 3664
rect 104164 3612 104216 3664
rect 109316 3612 109368 3664
rect 171784 3612 171836 3664
rect 6460 3544 6512 3596
rect 79324 3544 79376 3596
rect 85580 3544 85632 3596
rect 86500 3544 86552 3596
rect 93860 3544 93912 3596
rect 94780 3544 94832 3596
rect 103336 3544 103388 3596
rect 195428 3544 195480 3596
rect 242992 3544 243044 3596
rect 244924 3544 244976 3596
rect 267740 3544 267792 3596
rect 271972 3544 272024 3596
rect 316132 3544 316184 3596
rect 317328 3544 317380 3596
rect 2780 3476 2832 3528
rect 3700 3476 3752 3528
rect 19340 3476 19392 3528
rect 20260 3476 20312 3528
rect 33048 3476 33100 3528
rect 150624 3476 150676 3528
rect 242900 3476 242952 3528
rect 244096 3476 244148 3528
rect 307760 3476 307812 3528
rect 309048 3476 309100 3528
rect 332600 3476 332652 3528
rect 333888 3476 333940 3528
rect 24216 3408 24268 3460
rect 188528 3408 188580 3460
rect 276020 3408 276072 3460
rect 276756 3408 276808 3460
rect 44180 3340 44232 3392
rect 45100 3340 45152 3392
rect 52460 3340 52512 3392
rect 53380 3340 53432 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 118700 3340 118752 3392
rect 119896 3340 119948 3392
rect 1676 3272 1728 3324
rect 7748 3272 7800 3324
rect 235816 3068 235868 3120
rect 238024 3068 238076 3120
rect 292580 3000 292632 3052
rect 293960 3000 294012 3052
rect 43076 2116 43128 2168
rect 301504 2116 301556 2168
rect 30104 2048 30156 2100
rect 301596 2048 301648 2100
<< metal2 >>
rect 6932 703582 7972 703610
rect 6932 686526 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 697610 24348 703520
rect 40512 700398 40540 703520
rect 72988 702778 73016 703520
rect 82084 703248 82136 703254
rect 82084 703190 82136 703196
rect 79324 703044 79376 703050
rect 79324 702986 79376 702992
rect 78588 702840 78640 702846
rect 78588 702782 78640 702788
rect 71780 702772 71832 702778
rect 71780 702714 71832 702720
rect 72976 702772 73028 702778
rect 72976 702714 73028 702720
rect 69204 702636 69256 702642
rect 69204 702578 69256 702584
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 62028 700324 62080 700330
rect 62028 700266 62080 700272
rect 24308 697604 24360 697610
rect 24308 697546 24360 697552
rect 6920 686520 6972 686526
rect 6920 686462 6972 686468
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 59268 681896 59320 681902
rect 59268 681838 59320 681844
rect 57796 681828 57848 681834
rect 57796 681770 57848 681776
rect 4804 681760 4856 681766
rect 4804 681702 4856 681708
rect 55128 681760 55180 681766
rect 55128 681702 55180 681708
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 2780 658232 2832 658238
rect 2778 658200 2780 658209
rect 2832 658200 2834 658209
rect 2778 658135 2834 658144
rect 3436 638246 3464 671191
rect 4816 658238 4844 681702
rect 53748 681012 53800 681018
rect 53748 680954 53800 680960
rect 33048 676252 33100 676258
rect 33048 676194 33100 676200
rect 4804 658232 4856 658238
rect 4804 658174 4856 658180
rect 3424 638240 3476 638246
rect 3424 638182 3476 638188
rect 4068 635520 4120 635526
rect 4068 635462 4120 635468
rect 3424 634092 3476 634098
rect 3424 634034 3476 634040
rect 3436 606121 3464 634034
rect 4080 632097 4108 635462
rect 4066 632088 4122 632097
rect 4066 632023 4122 632032
rect 3514 619168 3570 619177
rect 3514 619103 3570 619112
rect 3528 618662 3556 619103
rect 3516 618656 3568 618662
rect 3516 618598 3568 618604
rect 7564 618656 7616 618662
rect 7564 618598 7616 618604
rect 3422 606112 3478 606121
rect 3422 606047 3478 606056
rect 7576 589966 7604 618598
rect 7564 589960 7616 589966
rect 7564 589902 7616 589908
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3238 566944 3294 566953
rect 3238 566879 3294 566888
rect 3252 565894 3280 566879
rect 3240 565888 3292 565894
rect 3240 565830 3292 565836
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3436 538898 3464 579935
rect 32956 573368 33008 573374
rect 32956 573310 33008 573316
rect 30288 567248 30340 567254
rect 30288 567190 30340 567196
rect 25504 565888 25556 565894
rect 25504 565830 25556 565836
rect 25516 545086 25544 565830
rect 25504 545080 25556 545086
rect 25504 545022 25556 545028
rect 3424 538892 3476 538898
rect 3424 538834 3476 538840
rect 3148 528556 3200 528562
rect 3148 528498 3200 528504
rect 3160 527921 3188 528498
rect 3146 527912 3202 527921
rect 3146 527847 3202 527856
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 11704 514820 11756 514826
rect 3424 514762 3476 514768
rect 11704 514762 11756 514768
rect 3146 501800 3202 501809
rect 3146 501735 3202 501744
rect 3160 497486 3188 501735
rect 11716 498846 11744 514762
rect 11704 498840 11756 498846
rect 11704 498782 11756 498788
rect 3148 497480 3200 497486
rect 3148 497422 3200 497428
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 11704 474768 11756 474774
rect 11704 474710 11756 474716
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 4804 462596 4856 462602
rect 2780 462538 2832 462544
rect 4804 462538 4856 462544
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 4816 438870 4844 462538
rect 11716 439210 11744 474710
rect 30300 468489 30328 567190
rect 32968 475386 32996 573310
rect 32956 475380 33008 475386
rect 32956 475322 33008 475328
rect 30286 468480 30342 468489
rect 30286 468415 30342 468424
rect 32956 458856 33008 458862
rect 32956 458798 33008 458804
rect 30288 451308 30340 451314
rect 30288 451250 30340 451256
rect 11704 439204 11756 439210
rect 11704 439146 11756 439152
rect 4804 438864 4856 438870
rect 4804 438806 4856 438812
rect 3424 429888 3476 429894
rect 3424 429830 3476 429836
rect 3436 410553 3464 429830
rect 3514 423600 3570 423609
rect 3514 423535 3570 423544
rect 3528 422346 3556 423535
rect 3516 422340 3568 422346
rect 3516 422282 3568 422288
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3422 397488 3478 397497
rect 3422 397423 3478 397432
rect 3436 392630 3464 397423
rect 3424 392624 3476 392630
rect 3424 392566 3476 392572
rect 4804 387864 4856 387870
rect 4804 387806 4856 387812
rect 3424 378820 3476 378826
rect 3424 378762 3476 378768
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 2780 346316 2832 346322
rect 2780 346258 2832 346264
rect 2792 345409 2820 346258
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 3436 319297 3464 378762
rect 3516 372564 3568 372570
rect 3516 372506 3568 372512
rect 3528 371385 3556 372506
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 4816 346322 4844 387806
rect 15844 357468 15896 357474
rect 15844 357410 15896 357416
rect 15856 346390 15884 357410
rect 30300 352617 30328 451250
rect 32968 360874 32996 458798
rect 32956 360868 33008 360874
rect 32956 360810 33008 360816
rect 30286 352608 30342 352617
rect 30286 352543 30342 352552
rect 21364 351960 21416 351966
rect 21364 351902 21416 351908
rect 15844 346384 15896 346390
rect 15844 346326 15896 346332
rect 4804 346316 4856 346322
rect 4804 346258 4856 346264
rect 7564 331288 7616 331294
rect 7564 331230 7616 331236
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 313954 3464 319223
rect 3424 313948 3476 313954
rect 3424 313890 3476 313896
rect 3424 306332 3476 306338
rect 3424 306274 3476 306280
rect 3436 306241 3464 306274
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 7576 293894 7604 331230
rect 21376 306338 21404 351902
rect 21364 306332 21416 306338
rect 21364 306274 21416 306280
rect 22744 299600 22796 299606
rect 22744 299542 22796 299548
rect 17224 297424 17276 297430
rect 17224 297366 17276 297372
rect 3424 293888 3476 293894
rect 3424 293830 3476 293836
rect 7564 293888 7616 293894
rect 7564 293830 7616 293836
rect 3436 293185 3464 293830
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 8208 292596 8260 292602
rect 8208 292538 8260 292544
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 248414 3464 254079
rect 3436 248386 3556 248414
rect 3424 241460 3476 241466
rect 3424 241402 3476 241408
rect 3436 241097 3464 241402
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3528 240106 3556 248386
rect 3516 240100 3568 240106
rect 3516 240042 3568 240048
rect 4804 229764 4856 229770
rect 4804 229706 4856 229712
rect 3424 225616 3476 225622
rect 3424 225558 3476 225564
rect 1306 224224 1362 224233
rect 1306 224159 1362 224168
rect 1320 19310 1348 224159
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3436 201929 3464 225558
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 4816 97782 4844 229706
rect 2780 97776 2832 97782
rect 2780 97718 2832 97724
rect 4804 97776 4856 97782
rect 4804 97718 4856 97724
rect 2792 97617 2820 97718
rect 2778 97608 2834 97617
rect 2778 97543 2834 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 6920 58676 6972 58682
rect 6920 58618 6972 58624
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 4160 51740 4212 51746
rect 4160 51682 4212 51688
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2780 36576 2832 36582
rect 2780 36518 2832 36524
rect 20 19304 72 19310
rect 20 19246 72 19252
rect 1308 19304 1360 19310
rect 1308 19246 1360 19252
rect 32 16574 60 19246
rect 32 16546 152 16574
rect 124 354 152 16546
rect 2792 3534 2820 36518
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 2872 24132 2924 24138
rect 2872 24074 2924 24080
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 1676 3324 1728 3330
rect 1676 3266 1728 3272
rect 1688 480 1716 3266
rect 2884 480 2912 24074
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 4172 16574 4200 51682
rect 6932 16574 6960 58618
rect 8220 16574 8248 292538
rect 14464 264240 14516 264246
rect 14464 264182 14516 264188
rect 14476 215286 14504 264182
rect 15844 257372 15896 257378
rect 15844 257314 15896 257320
rect 14464 215280 14516 215286
rect 14464 215222 14516 215228
rect 11704 209092 11756 209098
rect 11704 209034 11756 209040
rect 11716 111790 11744 209034
rect 14464 177336 14516 177342
rect 14464 177278 14516 177284
rect 11704 111784 11756 111790
rect 11704 111726 11756 111732
rect 11058 76528 11114 76537
rect 11058 76463 11114 76472
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 4172 16546 5304 16574
rect 6932 16546 7512 16574
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3436 6497 3464 8978
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3712 354 3740 3470
rect 5276 480 5304 16546
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6472 480 6500 3538
rect 7484 3482 7512 16546
rect 7760 16561 8248 16574
rect 7760 16552 8262 16561
rect 7760 16546 8206 16552
rect 7484 3454 7696 3482
rect 7668 480 7696 3454
rect 7760 3330 7788 16546
rect 8206 16487 8262 16496
rect 8760 7608 8812 7614
rect 8760 7550 8812 7556
rect 7748 3324 7800 3330
rect 7748 3266 7800 3272
rect 8772 480 8800 7550
rect 4038 354 4150 480
rect 3712 326 4150 354
rect 4038 -960 4150 326
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 22714
rect 11072 6914 11100 76463
rect 14476 45558 14504 177278
rect 15856 137970 15884 257314
rect 15844 137964 15896 137970
rect 15844 137906 15896 137912
rect 17236 59362 17264 297366
rect 21364 268388 21416 268394
rect 21364 268330 21416 268336
rect 17224 59356 17276 59362
rect 17224 59298 17276 59304
rect 19340 55888 19392 55894
rect 19340 55830 19392 55836
rect 15200 46300 15252 46306
rect 15200 46242 15252 46248
rect 14464 45552 14516 45558
rect 14464 45494 14516 45500
rect 11152 39364 11204 39370
rect 11152 39306 11204 39312
rect 11164 16574 11192 39306
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 13832 16574 13860 17206
rect 15212 16574 15240 46242
rect 17960 26920 18012 26926
rect 17960 26862 18012 26868
rect 11164 16546 11928 16574
rect 13832 16546 14320 16574
rect 15212 16546 15976 16574
rect 11072 6886 11192 6914
rect 11164 480 11192 6886
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 11900 354 11928 16546
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13556 480 13584 8910
rect 12318 354 12430 480
rect 11900 326 12430 354
rect 12318 -960 12430 326
rect 13514 -960 13626 480
rect 14292 354 14320 16546
rect 15948 480 15976 16546
rect 17040 14544 17092 14550
rect 17040 14486 17092 14492
rect 17052 480 17080 14486
rect 14710 354 14822 480
rect 14292 326 14822 354
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 26862
rect 19352 3534 19380 55830
rect 21376 33114 21404 268330
rect 21364 33108 21416 33114
rect 21364 33050 21416 33056
rect 19432 31068 19484 31074
rect 19432 31010 19484 31016
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19444 480 19472 31010
rect 20720 25560 20772 25566
rect 20720 25502 20772 25508
rect 20732 16574 20760 25502
rect 22756 20670 22784 299542
rect 25504 290488 25556 290494
rect 25504 290430 25556 290436
rect 25516 150414 25544 290430
rect 29644 279472 29696 279478
rect 29644 279414 29696 279420
rect 25504 150408 25556 150414
rect 25504 150350 25556 150356
rect 24860 50380 24912 50386
rect 24860 50322 24912 50328
rect 22744 20664 22796 20670
rect 22744 20606 22796 20612
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22112 16574 22140 19926
rect 24872 16574 24900 50322
rect 26240 37936 26292 37942
rect 26240 37878 26292 37884
rect 20732 16546 21864 16574
rect 22112 16546 22600 16574
rect 24872 16546 25360 16574
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20272 354 20300 3470
rect 21836 480 21864 16546
rect 20598 354 20710 480
rect 20272 326 20710 354
rect 20598 -960 20710 326
rect 21794 -960 21906 480
rect 22572 354 22600 16546
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24228 480 24256 3402
rect 25332 480 25360 16546
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26252 354 26280 37878
rect 29656 9042 29684 279414
rect 32404 253224 32456 253230
rect 32404 253166 32456 253172
rect 32416 85542 32444 253166
rect 32404 85536 32456 85542
rect 32404 85478 32456 85484
rect 31760 53168 31812 53174
rect 31760 53110 31812 53116
rect 30380 33788 30432 33794
rect 30380 33730 30432 33736
rect 30392 16574 30420 33730
rect 31772 16574 31800 53110
rect 30392 16546 30880 16574
rect 31772 16546 31984 16574
rect 29644 9036 29696 9042
rect 29644 8978 29696 8984
rect 28908 6180 28960 6186
rect 28908 6122 28960 6128
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 27724 480 27752 4762
rect 28920 480 28948 6122
rect 30104 2100 30156 2106
rect 30104 2042 30156 2048
rect 30116 480 30144 2042
rect 26486 354 26598 480
rect 26252 326 26598 354
rect 26486 -960 26598 326
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 16546
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 33060 3534 33088 676194
rect 48136 673532 48188 673538
rect 48136 673474 48188 673480
rect 44088 665304 44140 665310
rect 44088 665246 44140 665252
rect 42708 665236 42760 665242
rect 42708 665178 42760 665184
rect 39948 658980 40000 658986
rect 39948 658922 40000 658928
rect 34428 650072 34480 650078
rect 34428 650014 34480 650020
rect 34152 640348 34204 640354
rect 34152 640290 34204 640296
rect 33782 549264 33838 549273
rect 33782 549199 33838 549208
rect 33796 451314 33824 549199
rect 34164 541686 34192 640290
rect 34336 585200 34388 585206
rect 34336 585142 34388 585148
rect 34244 556912 34296 556918
rect 34244 556854 34296 556860
rect 34152 541680 34204 541686
rect 34152 541622 34204 541628
rect 34256 457502 34284 556854
rect 34348 485790 34376 585142
rect 34440 549273 34468 650014
rect 37096 645924 37148 645930
rect 37096 645866 37148 645872
rect 35714 586392 35770 586401
rect 35714 586327 35770 586336
rect 35624 579692 35676 579698
rect 35624 579634 35676 579640
rect 34426 549264 34482 549273
rect 34426 549199 34482 549208
rect 34336 485784 34388 485790
rect 34336 485726 34388 485732
rect 35532 483676 35584 483682
rect 35532 483618 35584 483624
rect 34336 472660 34388 472666
rect 34336 472602 34388 472608
rect 34244 457496 34296 457502
rect 34244 457438 34296 457444
rect 33784 451308 33836 451314
rect 33784 451250 33836 451256
rect 34348 376718 34376 472602
rect 35544 400994 35572 483618
rect 35636 479534 35664 579634
rect 35728 483682 35756 586327
rect 37004 581120 37056 581126
rect 37004 581062 37056 581068
rect 35808 575544 35860 575550
rect 35808 575486 35860 575492
rect 35716 483676 35768 483682
rect 35716 483618 35768 483624
rect 35624 479528 35676 479534
rect 35624 479470 35676 479476
rect 35716 456068 35768 456074
rect 35716 456010 35768 456016
rect 35622 447808 35678 447817
rect 35622 447743 35678 447752
rect 35532 400988 35584 400994
rect 35532 400930 35584 400936
rect 34428 400920 34480 400926
rect 34428 400862 34480 400868
rect 34336 376712 34388 376718
rect 34336 376654 34388 376660
rect 33784 294024 33836 294030
rect 33784 293966 33836 293972
rect 33796 164218 33824 293966
rect 34440 258058 34468 400862
rect 35532 362976 35584 362982
rect 35532 362918 35584 362924
rect 34428 258052 34480 258058
rect 34428 257994 34480 258000
rect 34440 257378 34468 257994
rect 34428 257372 34480 257378
rect 34428 257314 34480 257320
rect 34612 241460 34664 241466
rect 34612 241402 34664 241408
rect 34624 240786 34652 241402
rect 35544 240786 35572 362918
rect 35636 349110 35664 447743
rect 35728 357406 35756 456010
rect 35716 357400 35768 357406
rect 35716 357342 35768 357348
rect 35624 349104 35676 349110
rect 35624 349046 35676 349052
rect 34612 240780 34664 240786
rect 34612 240722 34664 240728
rect 35532 240780 35584 240786
rect 35532 240722 35584 240728
rect 33784 164212 33836 164218
rect 33784 164154 33836 164160
rect 33140 62824 33192 62830
rect 33140 62766 33192 62772
rect 33152 16574 33180 62766
rect 33152 16546 33640 16574
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33612 480 33640 16546
rect 34520 11756 34572 11762
rect 34520 11698 34572 11704
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 11698
rect 35820 6322 35848 575486
rect 36636 485852 36688 485858
rect 36636 485794 36688 485800
rect 36544 457496 36596 457502
rect 36544 457438 36596 457444
rect 36556 359514 36584 457438
rect 36648 403646 36676 485794
rect 37016 483002 37044 581062
rect 37108 546417 37136 645866
rect 37188 641776 37240 641782
rect 37188 641718 37240 641724
rect 37094 546408 37150 546417
rect 37094 546343 37150 546352
rect 37096 540388 37148 540394
rect 37096 540330 37148 540336
rect 37004 482996 37056 483002
rect 37004 482938 37056 482944
rect 37004 442740 37056 442746
rect 37004 442682 37056 442688
rect 37016 442270 37044 442682
rect 37004 442264 37056 442270
rect 37004 442206 37056 442212
rect 36636 403640 36688 403646
rect 36636 403582 36688 403588
rect 36544 359508 36596 359514
rect 36544 359450 36596 359456
rect 37016 341562 37044 442206
rect 37108 434654 37136 540330
rect 37200 525745 37228 641718
rect 38568 638988 38620 638994
rect 38568 638930 38620 638936
rect 38384 545148 38436 545154
rect 38384 545090 38436 545096
rect 37186 525736 37242 525745
rect 37186 525671 37242 525680
rect 37200 442746 37228 525671
rect 38396 445641 38424 545090
rect 38580 540394 38608 638930
rect 39764 632732 39816 632738
rect 39764 632674 39816 632680
rect 39672 582480 39724 582486
rect 39672 582422 39724 582428
rect 38568 540388 38620 540394
rect 38568 540330 38620 540336
rect 38476 539776 38528 539782
rect 38476 539718 38528 539724
rect 38382 445632 38438 445641
rect 38382 445567 38438 445576
rect 37188 442740 37240 442746
rect 37188 442682 37240 442688
rect 37096 434648 37148 434654
rect 37096 434590 37148 434596
rect 38488 431934 38516 539718
rect 38580 539646 38608 540330
rect 38568 539640 38620 539646
rect 38568 539582 38620 539588
rect 39684 488510 39712 582422
rect 39776 535430 39804 632674
rect 39960 557462 39988 658922
rect 41236 655580 41288 655586
rect 41236 655522 41288 655528
rect 41052 582412 41104 582418
rect 41052 582354 41104 582360
rect 39948 557456 40000 557462
rect 39948 557398 40000 557404
rect 39856 556844 39908 556850
rect 39856 556786 39908 556792
rect 39764 535424 39816 535430
rect 39764 535366 39816 535372
rect 39672 488504 39724 488510
rect 39672 488446 39724 488452
rect 39672 479528 39724 479534
rect 39672 479470 39724 479476
rect 38568 476128 38620 476134
rect 38568 476070 38620 476076
rect 38476 431928 38528 431934
rect 38476 431870 38528 431876
rect 38476 387116 38528 387122
rect 38476 387058 38528 387064
rect 37188 369912 37240 369918
rect 37188 369854 37240 369860
rect 37004 341556 37056 341562
rect 37004 341498 37056 341504
rect 37096 331900 37148 331906
rect 37096 331842 37148 331848
rect 37108 331294 37136 331842
rect 37096 331288 37148 331294
rect 37096 331230 37148 331236
rect 37108 244254 37136 331230
rect 37096 244248 37148 244254
rect 37096 244190 37148 244196
rect 35900 66904 35952 66910
rect 35900 66846 35952 66852
rect 35912 6914 35940 66846
rect 37200 53106 37228 369854
rect 38488 291174 38516 387058
rect 38108 291168 38160 291174
rect 38108 291110 38160 291116
rect 38476 291168 38528 291174
rect 38476 291110 38528 291116
rect 38120 290494 38148 291110
rect 38108 290488 38160 290494
rect 38108 290430 38160 290436
rect 37188 53100 37240 53106
rect 37188 53042 37240 53048
rect 37280 49020 37332 49026
rect 37280 48962 37332 48968
rect 35992 42084 36044 42090
rect 35992 42026 36044 42032
rect 36004 16574 36032 42026
rect 37292 16574 37320 48962
rect 38580 40866 38608 476070
rect 39304 394800 39356 394806
rect 39304 394742 39356 394748
rect 39316 372570 39344 394742
rect 39684 385150 39712 479470
rect 39776 439006 39804 535366
rect 39868 457570 39896 556786
rect 40684 553444 40736 553450
rect 40684 553386 40736 553392
rect 40696 539578 40724 553386
rect 40684 539572 40736 539578
rect 40684 539514 40736 539520
rect 39948 490612 40000 490618
rect 39948 490554 40000 490560
rect 39856 457564 39908 457570
rect 39856 457506 39908 457512
rect 39764 439000 39816 439006
rect 39764 438942 39816 438948
rect 39960 387258 39988 490554
rect 41064 489938 41092 582354
rect 41248 554742 41276 655522
rect 42524 629944 42576 629950
rect 42524 629886 42576 629892
rect 41326 586800 41382 586809
rect 41326 586735 41382 586744
rect 41236 554736 41288 554742
rect 41236 554678 41288 554684
rect 41144 547936 41196 547942
rect 41144 547878 41196 547884
rect 41052 489932 41104 489938
rect 41052 489874 41104 489880
rect 40960 481704 41012 481710
rect 40960 481646 41012 481652
rect 40972 406434 41000 481646
rect 40960 406428 41012 406434
rect 40960 406370 41012 406376
rect 41064 399498 41092 489874
rect 41156 448497 41184 547878
rect 41236 491972 41288 491978
rect 41236 491914 41288 491920
rect 41142 448488 41198 448497
rect 41142 448423 41198 448432
rect 41156 447817 41184 448423
rect 41142 447808 41198 447817
rect 41142 447743 41198 447752
rect 41052 399492 41104 399498
rect 41052 399434 41104 399440
rect 41248 391950 41276 491914
rect 41340 485790 41368 586735
rect 42536 533390 42564 629886
rect 42720 564398 42748 665178
rect 43996 627224 44048 627230
rect 43996 627166 44048 627172
rect 43810 585440 43866 585449
rect 43810 585375 43866 585384
rect 43718 568576 43774 568585
rect 43718 568511 43774 568520
rect 43732 567866 43760 568511
rect 42800 567860 42852 567866
rect 42800 567802 42852 567808
rect 43720 567860 43772 567866
rect 43720 567802 43772 567808
rect 42812 567254 42840 567802
rect 42800 567248 42852 567254
rect 42800 567190 42852 567196
rect 42708 564392 42760 564398
rect 42708 564334 42760 564340
rect 42616 559564 42668 559570
rect 42616 559506 42668 559512
rect 42524 533384 42576 533390
rect 42524 533326 42576 533332
rect 41328 485784 41380 485790
rect 41328 485726 41380 485732
rect 42628 459513 42656 559506
rect 42708 539504 42760 539510
rect 42708 539446 42760 539452
rect 42614 459504 42670 459513
rect 42614 459439 42670 459448
rect 41328 443692 41380 443698
rect 41328 443634 41380 443640
rect 41236 391944 41288 391950
rect 41236 391886 41288 391892
rect 41236 389836 41288 389842
rect 41236 389778 41288 389784
rect 39948 387252 40000 387258
rect 39948 387194 40000 387200
rect 39672 385144 39724 385150
rect 39672 385086 39724 385092
rect 39684 383654 39712 385086
rect 39948 383716 40000 383722
rect 39948 383658 40000 383664
rect 39684 383626 39896 383654
rect 39304 372564 39356 372570
rect 39304 372506 39356 372512
rect 39868 249082 39896 383626
rect 39856 249076 39908 249082
rect 39856 249018 39908 249024
rect 39960 240106 39988 383658
rect 41052 359508 41104 359514
rect 41052 359450 41104 359456
rect 41064 306338 41092 359450
rect 41144 356108 41196 356114
rect 41144 356050 41196 356056
rect 41052 306332 41104 306338
rect 41052 306274 41104 306280
rect 41156 280158 41184 356050
rect 41248 335170 41276 389778
rect 41340 344350 41368 443634
rect 42064 430636 42116 430642
rect 42064 430578 42116 430584
rect 41420 352572 41472 352578
rect 41420 352514 41472 352520
rect 41432 351966 41460 352514
rect 41420 351960 41472 351966
rect 41420 351902 41472 351908
rect 41328 344344 41380 344350
rect 41328 344286 41380 344292
rect 42076 337890 42104 430578
rect 42628 397458 42656 459439
rect 42720 434722 42748 539446
rect 43824 491978 43852 585375
rect 43904 573436 43956 573442
rect 43904 573378 43956 573384
rect 43812 491972 43864 491978
rect 43812 491914 43864 491920
rect 42800 488504 42852 488510
rect 42800 488446 42852 488452
rect 42708 434716 42760 434722
rect 42708 434658 42760 434664
rect 42708 432608 42760 432614
rect 42708 432550 42760 432556
rect 42720 431934 42748 432550
rect 42708 431928 42760 431934
rect 42708 431870 42760 431876
rect 42720 430642 42748 431870
rect 42708 430636 42760 430642
rect 42708 430578 42760 430584
rect 42812 400926 42840 488446
rect 43916 475454 43944 573378
rect 44008 557534 44036 627166
rect 44100 565146 44128 665246
rect 48044 652792 48096 652798
rect 48044 652734 48096 652740
rect 46848 638920 46900 638926
rect 46848 638862 46900 638868
rect 45376 636948 45428 636954
rect 45376 636890 45428 636896
rect 45284 630012 45336 630018
rect 45284 629954 45336 629960
rect 45190 588160 45246 588169
rect 45190 588095 45246 588104
rect 44088 565140 44140 565146
rect 44088 565082 44140 565088
rect 44008 557506 44128 557534
rect 44100 537878 44128 557506
rect 44088 537872 44140 537878
rect 44088 537814 44140 537820
rect 43996 537600 44048 537606
rect 43996 537542 44048 537548
rect 43904 475448 43956 475454
rect 43904 475390 43956 475396
rect 43812 433288 43864 433294
rect 43812 433230 43864 433236
rect 42800 400920 42852 400926
rect 42800 400862 42852 400868
rect 42616 397452 42668 397458
rect 42616 397394 42668 397400
rect 42708 382288 42760 382294
rect 42708 382230 42760 382236
rect 42616 352572 42668 352578
rect 42616 352514 42668 352520
rect 42064 337884 42116 337890
rect 42064 337826 42116 337832
rect 41236 335164 41288 335170
rect 41236 335106 41288 335112
rect 42628 316742 42656 352514
rect 42616 316736 42668 316742
rect 42616 316678 42668 316684
rect 41236 294092 41288 294098
rect 41236 294034 41288 294040
rect 40868 280152 40920 280158
rect 40868 280094 40920 280100
rect 41144 280152 41196 280158
rect 41144 280094 41196 280100
rect 40880 279478 40908 280094
rect 40868 279472 40920 279478
rect 40868 279414 40920 279420
rect 39948 240100 40000 240106
rect 39948 240042 40000 240048
rect 39960 238814 39988 240042
rect 39948 238808 40000 238814
rect 39948 238750 40000 238756
rect 41248 214674 41276 294034
rect 41328 293276 41380 293282
rect 41328 293218 41380 293224
rect 41236 214668 41288 214674
rect 41236 214610 41288 214616
rect 41340 71738 41368 293218
rect 42720 77994 42748 382230
rect 42800 380180 42852 380186
rect 42800 380122 42852 380128
rect 42812 378826 42840 380122
rect 42800 378820 42852 378826
rect 42800 378762 42852 378768
rect 42800 360868 42852 360874
rect 42800 360810 42852 360816
rect 42812 360262 42840 360810
rect 42800 360256 42852 360262
rect 42800 360198 42852 360204
rect 43824 340202 43852 433230
rect 43916 380186 43944 475390
rect 44008 437238 44036 537542
rect 43996 437232 44048 437238
rect 43996 437174 44048 437180
rect 44100 433294 44128 537814
rect 45204 530602 45232 588095
rect 45296 539782 45324 629954
rect 45284 539776 45336 539782
rect 45284 539718 45336 539724
rect 45388 539510 45416 636890
rect 46756 627360 46808 627366
rect 46756 627302 46808 627308
rect 46570 586664 46626 586673
rect 46570 586599 46626 586608
rect 45468 554668 45520 554674
rect 45468 554610 45520 554616
rect 45376 539504 45428 539510
rect 45376 539446 45428 539452
rect 45376 537532 45428 537538
rect 45376 537474 45428 537480
rect 45284 533384 45336 533390
rect 45284 533326 45336 533332
rect 45192 530596 45244 530602
rect 45192 530538 45244 530544
rect 45192 438320 45244 438326
rect 45192 438262 45244 438268
rect 44088 433288 44140 433294
rect 44088 433230 44140 433236
rect 43996 392216 44048 392222
rect 43996 392158 44048 392164
rect 43904 380180 43956 380186
rect 43904 380122 43956 380128
rect 43904 364404 43956 364410
rect 43904 364346 43956 364352
rect 43812 340196 43864 340202
rect 43812 340138 43864 340144
rect 43812 284368 43864 284374
rect 43812 284310 43864 284316
rect 43824 229090 43852 284310
rect 43916 264246 43944 364346
rect 44008 282878 44036 392158
rect 44088 360256 44140 360262
rect 44088 360198 44140 360204
rect 43996 282872 44048 282878
rect 43996 282814 44048 282820
rect 43904 264240 43956 264246
rect 43904 264182 43956 264188
rect 43812 229084 43864 229090
rect 43812 229026 43864 229032
rect 42708 77988 42760 77994
rect 42708 77930 42760 77936
rect 41328 71732 41380 71738
rect 41328 71674 41380 71680
rect 40040 65544 40092 65550
rect 40040 65486 40092 65492
rect 38568 40860 38620 40866
rect 38568 40802 38620 40808
rect 40052 16574 40080 65486
rect 44100 35222 44128 360198
rect 45204 337958 45232 438262
rect 45296 436082 45324 533326
rect 45388 451274 45416 537474
rect 45480 451926 45508 554610
rect 46480 536920 46532 536926
rect 46480 536862 46532 536868
rect 45468 451920 45520 451926
rect 45468 451862 45520 451868
rect 45388 451246 45508 451274
rect 45480 438274 45508 451246
rect 45480 438258 45600 438274
rect 45480 438252 45612 438258
rect 45480 438246 45560 438252
rect 45560 438194 45612 438200
rect 46204 438252 46256 438258
rect 46204 438194 46256 438200
rect 45284 436076 45336 436082
rect 45284 436018 45336 436024
rect 45468 436076 45520 436082
rect 45468 436018 45520 436024
rect 45284 345092 45336 345098
rect 45284 345034 45336 345040
rect 45192 337952 45244 337958
rect 45192 337894 45244 337900
rect 45296 268462 45324 345034
rect 45480 333878 45508 436018
rect 46216 339318 46244 438194
rect 46492 437374 46520 536862
rect 46584 490618 46612 586599
rect 46664 534132 46716 534138
rect 46664 534074 46716 534080
rect 46572 490612 46624 490618
rect 46572 490554 46624 490560
rect 46676 438802 46704 534074
rect 46768 529922 46796 627302
rect 46860 536110 46888 638862
rect 47952 585812 48004 585818
rect 47952 585754 48004 585760
rect 47964 585585 47992 585754
rect 47950 585576 48006 585585
rect 47950 585511 48006 585520
rect 47952 585268 48004 585274
rect 47952 585210 48004 585216
rect 46848 536104 46900 536110
rect 46848 536046 46900 536052
rect 46756 529916 46808 529922
rect 46756 529858 46808 529864
rect 47964 492658 47992 585210
rect 48056 554674 48084 652734
rect 48148 574054 48176 673474
rect 52368 663808 52420 663814
rect 52368 663750 52420 663756
rect 50804 659728 50856 659734
rect 50804 659670 50856 659676
rect 49608 656940 49660 656946
rect 49608 656882 49660 656888
rect 48228 638308 48280 638314
rect 48228 638250 48280 638256
rect 48136 574048 48188 574054
rect 48136 573990 48188 573996
rect 48148 573374 48176 573990
rect 48136 573368 48188 573374
rect 48136 573310 48188 573316
rect 48136 561672 48188 561678
rect 48136 561614 48188 561620
rect 48044 554668 48096 554674
rect 48044 554610 48096 554616
rect 48044 540252 48096 540258
rect 48044 540194 48096 540200
rect 47952 492652 48004 492658
rect 47952 492594 48004 492600
rect 47860 492108 47912 492114
rect 47860 492050 47912 492056
rect 47676 459604 47728 459610
rect 47676 459546 47728 459552
rect 46756 451920 46808 451926
rect 46756 451862 46808 451868
rect 46664 438796 46716 438802
rect 46664 438738 46716 438744
rect 46480 437368 46532 437374
rect 46480 437310 46532 437316
rect 46768 396030 46796 451862
rect 47584 434648 47636 434654
rect 47584 434590 47636 434596
rect 46848 396772 46900 396778
rect 46848 396714 46900 396720
rect 46756 396024 46808 396030
rect 46756 395966 46808 395972
rect 46756 392692 46808 392698
rect 46756 392634 46808 392640
rect 46664 339448 46716 339454
rect 46664 339390 46716 339396
rect 46204 339312 46256 339318
rect 46204 339254 46256 339260
rect 45468 333872 45520 333878
rect 45468 333814 45520 333820
rect 45376 311160 45428 311166
rect 45376 311102 45428 311108
rect 45284 268456 45336 268462
rect 45284 268398 45336 268404
rect 45388 244186 45416 311102
rect 45468 280220 45520 280226
rect 45468 280162 45520 280168
rect 45376 244180 45428 244186
rect 45376 244122 45428 244128
rect 45480 202298 45508 280162
rect 46676 245546 46704 339390
rect 46768 332586 46796 392634
rect 46860 336734 46888 396714
rect 46848 336728 46900 336734
rect 46848 336670 46900 336676
rect 47596 336394 47624 434590
rect 47688 364410 47716 459546
rect 47872 393990 47900 492050
rect 48056 440298 48084 540194
rect 48148 460222 48176 561614
rect 48240 535294 48268 638250
rect 49332 627292 49384 627298
rect 49332 627234 49384 627240
rect 48228 535288 48280 535294
rect 48228 535230 48280 535236
rect 48240 534138 48268 535230
rect 49344 535226 49372 627234
rect 49424 583772 49476 583778
rect 49424 583714 49476 583720
rect 49332 535220 49384 535226
rect 49332 535162 49384 535168
rect 49344 534177 49372 535162
rect 49330 534168 49386 534177
rect 48228 534132 48280 534138
rect 49330 534103 49386 534112
rect 48228 534074 48280 534080
rect 48228 492652 48280 492658
rect 48228 492594 48280 492600
rect 48240 491502 48268 492594
rect 49436 492114 49464 583714
rect 49516 563100 49568 563106
rect 49516 563042 49568 563048
rect 49424 492108 49476 492114
rect 49424 492050 49476 492056
rect 48228 491496 48280 491502
rect 48228 491438 48280 491444
rect 48136 460216 48188 460222
rect 48136 460158 48188 460164
rect 48148 459610 48176 460158
rect 48136 459604 48188 459610
rect 48136 459546 48188 459552
rect 48044 440292 48096 440298
rect 48044 440234 48096 440240
rect 48136 435396 48188 435402
rect 48136 435338 48188 435344
rect 48148 434654 48176 435338
rect 48136 434648 48188 434654
rect 48136 434590 48188 434596
rect 47860 393984 47912 393990
rect 47860 393926 47912 393932
rect 48240 386510 48268 491438
rect 48964 490000 49016 490006
rect 48964 489942 49016 489948
rect 48976 489841 49004 489942
rect 48962 489832 49018 489841
rect 48962 489767 49018 489776
rect 48976 402257 49004 489767
rect 49528 464370 49556 563042
rect 49620 557530 49648 656882
rect 50712 635588 50764 635594
rect 50712 635530 50764 635536
rect 50344 557592 50396 557598
rect 50344 557534 50396 557540
rect 49608 557524 49660 557530
rect 49608 557466 49660 557472
rect 49620 556918 49648 557466
rect 49608 556912 49660 556918
rect 49608 556854 49660 556860
rect 49608 536852 49660 536858
rect 49608 536794 49660 536800
rect 49516 464364 49568 464370
rect 49516 464306 49568 464312
rect 48962 402248 49018 402257
rect 48962 402183 49018 402192
rect 49424 399628 49476 399634
rect 49424 399570 49476 399576
rect 48228 386504 48280 386510
rect 48228 386446 48280 386452
rect 48136 385076 48188 385082
rect 48136 385018 48188 385024
rect 47676 364404 47728 364410
rect 47676 364346 47728 364352
rect 47584 336388 47636 336394
rect 47584 336330 47636 336336
rect 48044 334008 48096 334014
rect 48044 333950 48096 333956
rect 46756 332580 46808 332586
rect 46756 332522 46808 332528
rect 46756 287088 46808 287094
rect 46756 287030 46808 287036
rect 46664 245540 46716 245546
rect 46664 245482 46716 245488
rect 46768 207670 46796 287030
rect 47952 277432 48004 277438
rect 47952 277374 48004 277380
rect 46756 207664 46808 207670
rect 46756 207606 46808 207612
rect 45468 202292 45520 202298
rect 45468 202234 45520 202240
rect 47964 188358 47992 277374
rect 48056 238678 48084 333950
rect 48148 267714 48176 385018
rect 48136 267708 48188 267714
rect 48136 267650 48188 267656
rect 48044 238672 48096 238678
rect 48044 238614 48096 238620
rect 48240 235958 48268 386446
rect 49436 338026 49464 399570
rect 49528 368558 49556 464306
rect 49620 438870 49648 536794
rect 50356 458182 50384 557534
rect 50724 538150 50752 635530
rect 50816 561678 50844 659670
rect 52276 637016 52328 637022
rect 52276 636958 52328 636964
rect 50988 636880 51040 636886
rect 50988 636822 51040 636828
rect 50896 578944 50948 578950
rect 50896 578886 50948 578892
rect 50804 561672 50856 561678
rect 50804 561614 50856 561620
rect 50712 538144 50764 538150
rect 50712 538086 50764 538092
rect 50724 536926 50752 538086
rect 50712 536920 50764 536926
rect 50712 536862 50764 536868
rect 50620 536716 50672 536722
rect 50620 536658 50672 536664
rect 50344 458176 50396 458182
rect 50344 458118 50396 458124
rect 50528 457564 50580 457570
rect 50528 457506 50580 457512
rect 50540 456822 50568 457506
rect 50528 456816 50580 456822
rect 50528 456758 50580 456764
rect 49608 438864 49660 438870
rect 49608 438806 49660 438812
rect 49620 438190 49648 438806
rect 49608 438184 49660 438190
rect 49608 438126 49660 438132
rect 50632 437306 50660 536658
rect 50908 478990 50936 578886
rect 51000 534070 51028 636822
rect 52092 632800 52144 632806
rect 52092 632742 52144 632748
rect 52104 538966 52132 632742
rect 52182 583944 52238 583953
rect 52182 583879 52238 583888
rect 52092 538960 52144 538966
rect 52092 538902 52144 538908
rect 51724 536104 51776 536110
rect 51724 536046 51776 536052
rect 50988 534064 51040 534070
rect 50988 534006 51040 534012
rect 50896 478984 50948 478990
rect 50896 478926 50948 478932
rect 50896 456816 50948 456822
rect 50896 456758 50948 456764
rect 50802 438832 50858 438841
rect 50802 438767 50858 438776
rect 50712 438184 50764 438190
rect 50712 438126 50764 438132
rect 50620 437300 50672 437306
rect 50620 437242 50672 437248
rect 49608 389224 49660 389230
rect 49608 389166 49660 389172
rect 49516 368552 49568 368558
rect 49516 368494 49568 368500
rect 49424 338020 49476 338026
rect 49424 337962 49476 337968
rect 48320 306332 48372 306338
rect 48320 306274 48372 306280
rect 48332 253910 48360 306274
rect 49620 298897 49648 389166
rect 50724 337754 50752 438126
rect 50712 337748 50764 337754
rect 50712 337690 50764 337696
rect 50816 336462 50844 438767
rect 50908 359582 50936 456758
rect 50988 440292 51040 440298
rect 50988 440234 51040 440240
rect 51000 438841 51028 440234
rect 50986 438832 51042 438841
rect 50986 438767 51042 438776
rect 51736 438666 51764 536046
rect 52196 499574 52224 583879
rect 52288 538014 52316 636958
rect 52380 564330 52408 663750
rect 53656 661700 53708 661706
rect 53656 661642 53708 661648
rect 53564 584452 53616 584458
rect 53564 584394 53616 584400
rect 53576 583817 53604 584394
rect 53562 583808 53618 583817
rect 53562 583743 53618 583752
rect 53472 582548 53524 582554
rect 53472 582490 53524 582496
rect 52368 564324 52420 564330
rect 52368 564266 52420 564272
rect 52380 563106 52408 564266
rect 52368 563100 52420 563106
rect 52368 563042 52420 563048
rect 52366 539472 52422 539481
rect 52366 539407 52368 539416
rect 52420 539407 52422 539416
rect 52368 539378 52420 539384
rect 52276 538008 52328 538014
rect 52276 537950 52328 537956
rect 52288 537606 52316 537950
rect 52276 537600 52328 537606
rect 52276 537542 52328 537548
rect 52196 499546 52408 499574
rect 52276 491428 52328 491434
rect 52276 491370 52328 491376
rect 52182 488608 52238 488617
rect 52182 488543 52238 488552
rect 52196 488510 52224 488543
rect 52184 488504 52236 488510
rect 52184 488446 52236 488452
rect 52184 478984 52236 478990
rect 52184 478926 52236 478932
rect 51724 438660 51776 438666
rect 51724 438602 51776 438608
rect 51736 438326 51764 438602
rect 51724 438320 51776 438326
rect 51724 438262 51776 438268
rect 52000 398132 52052 398138
rect 52000 398074 52052 398080
rect 50986 390824 51042 390833
rect 50986 390759 51042 390768
rect 51000 390726 51028 390759
rect 50988 390720 51040 390726
rect 50988 390662 51040 390668
rect 50896 359576 50948 359582
rect 50896 359518 50948 359524
rect 50804 336456 50856 336462
rect 50804 336398 50856 336404
rect 50804 322380 50856 322386
rect 50804 322322 50856 322328
rect 49606 298888 49662 298897
rect 49606 298823 49662 298832
rect 49608 294160 49660 294166
rect 49608 294102 49660 294108
rect 48320 253904 48372 253910
rect 48320 253846 48372 253852
rect 48964 253904 49016 253910
rect 48964 253846 49016 253852
rect 48976 253230 49004 253846
rect 48964 253224 49016 253230
rect 48964 253166 49016 253172
rect 48228 235952 48280 235958
rect 48228 235894 48280 235900
rect 49620 210361 49648 294102
rect 50816 245614 50844 322322
rect 50804 245608 50856 245614
rect 50804 245550 50856 245556
rect 50908 234530 50936 359518
rect 51000 255270 51028 390662
rect 52012 333946 52040 398074
rect 52092 394120 52144 394126
rect 52092 394062 52144 394068
rect 52104 339250 52132 394062
rect 52196 393314 52224 478926
rect 52288 399566 52316 491370
rect 52380 487830 52408 499546
rect 53484 492658 53512 582490
rect 53564 581052 53616 581058
rect 53564 580994 53616 581000
rect 53472 492652 53524 492658
rect 53472 492594 53524 492600
rect 52368 487824 52420 487830
rect 52368 487766 52420 487772
rect 52276 399560 52328 399566
rect 52276 399502 52328 399508
rect 52196 393286 52316 393314
rect 52288 388006 52316 393286
rect 52380 388482 52408 487766
rect 53576 485110 53604 580994
rect 53668 562358 53696 661642
rect 53760 638926 53788 680954
rect 55036 674960 55088 674966
rect 55036 674902 55088 674908
rect 53748 638920 53800 638926
rect 53748 638862 53800 638868
rect 54760 638376 54812 638382
rect 54760 638318 54812 638324
rect 53748 634160 53800 634166
rect 53748 634102 53800 634108
rect 53656 562352 53708 562358
rect 53656 562294 53708 562300
rect 53760 535362 53788 634102
rect 53840 574796 53892 574802
rect 53840 574738 53892 574744
rect 53852 573442 53880 574738
rect 53840 573436 53892 573442
rect 53840 573378 53892 573384
rect 54484 562352 54536 562358
rect 54484 562294 54536 562300
rect 53748 535356 53800 535362
rect 53748 535298 53800 535304
rect 53656 492652 53708 492658
rect 53656 492594 53708 492600
rect 53668 491366 53696 492594
rect 53656 491360 53708 491366
rect 53656 491302 53708 491308
rect 53564 485104 53616 485110
rect 53564 485046 53616 485052
rect 53472 398200 53524 398206
rect 53472 398142 53524 398148
rect 52460 392624 52512 392630
rect 52460 392566 52512 392572
rect 52472 392018 52500 392566
rect 52460 392012 52512 392018
rect 52460 391954 52512 391960
rect 52368 388476 52420 388482
rect 52368 388418 52420 388424
rect 52276 388000 52328 388006
rect 52276 387942 52328 387948
rect 52184 387184 52236 387190
rect 52184 387126 52236 387132
rect 52196 339454 52224 387126
rect 52184 339448 52236 339454
rect 52184 339390 52236 339396
rect 52092 339244 52144 339250
rect 52092 339186 52144 339192
rect 52184 336592 52236 336598
rect 52184 336534 52236 336540
rect 52000 333940 52052 333946
rect 52000 333882 52052 333888
rect 52092 324964 52144 324970
rect 52092 324906 52144 324912
rect 52104 274650 52132 324906
rect 52092 274644 52144 274650
rect 52092 274586 52144 274592
rect 52092 268456 52144 268462
rect 52092 268398 52144 268404
rect 52104 267034 52132 268398
rect 52092 267028 52144 267034
rect 52092 266970 52144 266976
rect 50988 255264 51040 255270
rect 50988 255206 51040 255212
rect 50896 234524 50948 234530
rect 50896 234466 50948 234472
rect 52104 224942 52132 266970
rect 52196 255202 52224 336534
rect 52288 279478 52316 387942
rect 53484 335238 53512 398142
rect 53576 391270 53604 485046
rect 53668 402974 53696 491302
rect 53760 439550 53788 535298
rect 53840 485920 53892 485926
rect 53840 485862 53892 485868
rect 53852 485790 53880 485862
rect 53840 485784 53892 485790
rect 53840 485726 53892 485732
rect 53748 439544 53800 439550
rect 53748 439486 53800 439492
rect 53668 402946 53788 402974
rect 53656 392012 53708 392018
rect 53656 391954 53708 391960
rect 53564 391264 53616 391270
rect 53564 391206 53616 391212
rect 53564 385688 53616 385694
rect 53564 385630 53616 385636
rect 53576 335306 53604 385630
rect 53668 383654 53696 391954
rect 53760 388090 53788 402946
rect 53852 389230 53880 485726
rect 54496 463010 54524 562294
rect 54772 536722 54800 638318
rect 54944 632936 54996 632942
rect 54944 632878 54996 632884
rect 54850 585304 54906 585313
rect 54850 585239 54906 585248
rect 54760 536716 54812 536722
rect 54760 536658 54812 536664
rect 54864 492794 54892 585239
rect 54956 538082 54984 632878
rect 55048 574802 55076 674902
rect 55140 635662 55168 681702
rect 56508 657008 56560 657014
rect 56508 656950 56560 656956
rect 56324 635724 56376 635730
rect 56324 635666 56376 635672
rect 55128 635656 55180 635662
rect 55128 635598 55180 635604
rect 56232 582616 56284 582622
rect 56232 582558 56284 582564
rect 55036 574796 55088 574802
rect 55036 574738 55088 574744
rect 54944 538076 54996 538082
rect 54944 538018 54996 538024
rect 54956 536858 54984 538018
rect 54944 536852 54996 536858
rect 54944 536794 54996 536800
rect 55036 534064 55088 534070
rect 55036 534006 55088 534012
rect 55048 533633 55076 534006
rect 55034 533624 55090 533633
rect 55034 533559 55090 533568
rect 56244 533458 56272 582558
rect 56336 537946 56364 635666
rect 56416 583840 56468 583846
rect 56416 583782 56468 583788
rect 56428 558890 56456 583782
rect 56416 558884 56468 558890
rect 56416 558826 56468 558832
rect 56520 557462 56548 656950
rect 57808 643754 57836 681770
rect 59084 659796 59136 659802
rect 59084 659738 59136 659744
rect 58624 654832 58676 654838
rect 58624 654774 58676 654780
rect 57888 652860 57940 652866
rect 57888 652802 57940 652808
rect 57796 643748 57848 643754
rect 57796 643690 57848 643696
rect 57796 638444 57848 638450
rect 57796 638386 57848 638392
rect 57704 632868 57756 632874
rect 57704 632810 57756 632816
rect 57612 581664 57664 581670
rect 57612 581606 57664 581612
rect 56508 557456 56560 557462
rect 56508 557398 56560 557404
rect 56520 556850 56548 557398
rect 56508 556844 56560 556850
rect 56508 556786 56560 556792
rect 56508 556232 56560 556238
rect 56508 556174 56560 556180
rect 56414 543008 56470 543017
rect 56414 542943 56470 542952
rect 56324 537940 56376 537946
rect 56324 537882 56376 537888
rect 56336 537538 56364 537882
rect 56324 537532 56376 537538
rect 56324 537474 56376 537480
rect 56232 533452 56284 533458
rect 56232 533394 56284 533400
rect 56324 494760 56376 494766
rect 56324 494702 56376 494708
rect 54852 492788 54904 492794
rect 54852 492730 54904 492736
rect 55128 492788 55180 492794
rect 55128 492730 55180 492736
rect 54944 465724 54996 465730
rect 54944 465666 54996 465672
rect 54484 463004 54536 463010
rect 54484 462946 54536 462952
rect 54760 394052 54812 394058
rect 54760 393994 54812 394000
rect 53840 389224 53892 389230
rect 53840 389166 53892 389172
rect 53852 388618 53880 389166
rect 53840 388612 53892 388618
rect 53840 388554 53892 388560
rect 53760 388062 53880 388090
rect 53746 387968 53802 387977
rect 53746 387903 53748 387912
rect 53800 387903 53802 387912
rect 53748 387874 53800 387880
rect 53852 387818 53880 388062
rect 53760 387790 53880 387818
rect 53760 385082 53788 387790
rect 53748 385076 53800 385082
rect 53748 385018 53800 385024
rect 53668 383626 53788 383654
rect 53656 368552 53708 368558
rect 53656 368494 53708 368500
rect 53564 335300 53616 335306
rect 53564 335242 53616 335248
rect 53472 335232 53524 335238
rect 53472 335174 53524 335180
rect 53576 334014 53604 335242
rect 53564 334008 53616 334014
rect 53564 333950 53616 333956
rect 52368 302932 52420 302938
rect 52368 302874 52420 302880
rect 52276 279472 52328 279478
rect 52276 279414 52328 279420
rect 52276 273284 52328 273290
rect 52276 273226 52328 273232
rect 52184 255196 52236 255202
rect 52184 255138 52236 255144
rect 52092 224936 52144 224942
rect 52092 224878 52144 224884
rect 49606 210352 49662 210361
rect 49606 210287 49662 210296
rect 52288 189854 52316 273226
rect 52276 189848 52328 189854
rect 52276 189790 52328 189796
rect 47952 188352 48004 188358
rect 47952 188294 48004 188300
rect 52380 68338 52408 302874
rect 53668 301510 53696 368494
rect 53656 301504 53708 301510
rect 53656 301446 53708 301452
rect 53562 300112 53618 300121
rect 53562 300047 53618 300056
rect 53104 292732 53156 292738
rect 53104 292674 53156 292680
rect 52460 269068 52512 269074
rect 52460 269010 52512 269016
rect 52472 268394 52500 269010
rect 52460 268388 52512 268394
rect 52460 268330 52512 268336
rect 53116 189038 53144 292674
rect 53576 269074 53604 300047
rect 53656 274712 53708 274718
rect 53656 274654 53708 274660
rect 53564 269068 53616 269074
rect 53564 269010 53616 269016
rect 53564 255332 53616 255338
rect 53564 255274 53616 255280
rect 53576 233102 53604 255274
rect 53564 233096 53616 233102
rect 53564 233038 53616 233044
rect 53668 199510 53696 274654
rect 53760 238746 53788 383626
rect 54772 336598 54800 393994
rect 54852 385756 54904 385762
rect 54852 385698 54904 385704
rect 54864 339522 54892 385698
rect 54956 370530 54984 465666
rect 55140 393314 55168 492730
rect 55864 458244 55916 458250
rect 55864 458186 55916 458192
rect 55680 444372 55732 444378
rect 55680 444314 55732 444320
rect 55692 443698 55720 444314
rect 55680 443692 55732 443698
rect 55680 443634 55732 443640
rect 55876 394738 55904 458186
rect 56336 436014 56364 494702
rect 56428 444378 56456 542943
rect 56520 455394 56548 556174
rect 57624 553489 57652 581606
rect 57610 553480 57666 553489
rect 57610 553415 57666 553424
rect 57612 553376 57664 553382
rect 57612 553318 57664 553324
rect 57244 552696 57296 552702
rect 57244 552638 57296 552644
rect 56508 455388 56560 455394
rect 56508 455330 56560 455336
rect 57256 454442 57284 552638
rect 57336 530664 57388 530670
rect 57336 530606 57388 530612
rect 57348 529922 57376 530606
rect 57336 529916 57388 529922
rect 57336 529858 57388 529864
rect 56508 454436 56560 454442
rect 56508 454378 56560 454384
rect 57244 454436 57296 454442
rect 57244 454378 57296 454384
rect 56520 453354 56548 454378
rect 56508 453348 56560 453354
rect 56508 453290 56560 453296
rect 56416 444372 56468 444378
rect 56416 444314 56468 444320
rect 56324 436008 56376 436014
rect 56324 435950 56376 435956
rect 55956 396092 56008 396098
rect 55956 396034 56008 396040
rect 55864 394732 55916 394738
rect 55864 394674 55916 394680
rect 55048 393286 55168 393314
rect 55048 389230 55076 393286
rect 55036 389224 55088 389230
rect 55036 389166 55088 389172
rect 54944 370524 54996 370530
rect 54944 370466 54996 370472
rect 54852 339516 54904 339522
rect 54852 339458 54904 339464
rect 54760 336592 54812 336598
rect 54760 336534 54812 336540
rect 54852 334620 54904 334626
rect 54852 334562 54904 334568
rect 54760 295996 54812 296002
rect 54760 295938 54812 295944
rect 54484 266416 54536 266422
rect 54484 266358 54536 266364
rect 53748 238740 53800 238746
rect 53748 238682 53800 238688
rect 54496 235890 54524 266358
rect 54484 235884 54536 235890
rect 54484 235826 54536 235832
rect 53656 199504 53708 199510
rect 53656 199446 53708 199452
rect 53104 189032 53156 189038
rect 53104 188974 53156 188980
rect 53840 75200 53892 75206
rect 53840 75142 53892 75148
rect 52368 68332 52420 68338
rect 52368 68274 52420 68280
rect 45558 61568 45614 61577
rect 45558 61503 45614 61512
rect 44088 35216 44140 35222
rect 44088 35158 44140 35164
rect 41420 33856 41472 33862
rect 41420 33798 41472 33804
rect 41432 16574 41460 33798
rect 44180 28280 44232 28286
rect 44180 28222 44232 28228
rect 36004 16546 36768 16574
rect 37292 16546 38424 16574
rect 40052 16546 40264 16574
rect 41432 16546 41920 16574
rect 35912 6886 36032 6914
rect 35808 6316 35860 6322
rect 35808 6258 35860 6264
rect 36004 480 36032 6886
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 16546
rect 38396 480 38424 16546
rect 39120 14612 39172 14618
rect 39120 14554 39172 14560
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 14554
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 16546
rect 41892 480 41920 16546
rect 44192 3398 44220 28222
rect 45572 16574 45600 61503
rect 52460 60104 52512 60110
rect 52460 60046 52512 60052
rect 49700 58744 49752 58750
rect 49700 58686 49752 58692
rect 46940 55956 46992 55962
rect 46940 55898 46992 55904
rect 46952 16574 46980 55898
rect 48320 44872 48372 44878
rect 48320 44814 48372 44820
rect 48332 16574 48360 44814
rect 49712 16574 49740 58686
rect 51080 54664 51132 54670
rect 51080 54606 51132 54612
rect 45572 16546 46704 16574
rect 46952 16546 47440 16574
rect 48332 16546 48544 16574
rect 49712 16546 50200 16574
rect 44270 13016 44326 13025
rect 44270 12951 44326 12960
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 43076 2168 43128 2174
rect 43076 2110 43128 2116
rect 43088 480 43116 2110
rect 44284 480 44312 12951
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45112 354 45140 3334
rect 46676 480 46704 16546
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47412 354 47440 16546
rect 47830 354 47942 480
rect 47412 326 47942 354
rect 48516 354 48544 16546
rect 50172 480 50200 16546
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 47830 -960 47942 326
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51092 354 51120 54606
rect 52472 3398 52500 60046
rect 52552 57248 52604 57254
rect 52552 57190 52604 57196
rect 52460 3392 52512 3398
rect 52460 3334 52512 3340
rect 52564 480 52592 57190
rect 53852 16574 53880 75142
rect 54772 69766 54800 295938
rect 54864 266354 54892 334562
rect 54956 322318 54984 370466
rect 54944 322312 54996 322318
rect 54944 322254 54996 322260
rect 54852 266348 54904 266354
rect 54852 266290 54904 266296
rect 54944 264988 54996 264994
rect 54944 264930 54996 264936
rect 54956 231742 54984 264930
rect 55048 240106 55076 389166
rect 55968 355366 55996 396034
rect 56416 392624 56468 392630
rect 56416 392566 56468 392572
rect 55956 355360 56008 355366
rect 55956 355302 56008 355308
rect 55968 354674 55996 355302
rect 55968 354646 56272 354674
rect 55128 329180 55180 329186
rect 55128 329122 55180 329128
rect 55140 287026 55168 329122
rect 56244 308417 56272 354646
rect 56428 336666 56456 392566
rect 56520 355434 56548 453290
rect 57348 435946 57376 529858
rect 57624 454034 57652 553318
rect 57716 536654 57744 632810
rect 57808 538121 57836 638386
rect 57900 552702 57928 652802
rect 58636 556238 58664 654774
rect 58992 561604 59044 561610
rect 58992 561546 59044 561552
rect 58716 558884 58768 558890
rect 58716 558826 58768 558832
rect 58624 556232 58676 556238
rect 58624 556174 58676 556180
rect 57888 552696 57940 552702
rect 57888 552638 57940 552644
rect 57794 538112 57850 538121
rect 57794 538047 57850 538056
rect 57704 536648 57756 536654
rect 57704 536590 57756 536596
rect 57704 455388 57756 455394
rect 57704 455330 57756 455336
rect 57716 454102 57744 455330
rect 57704 454096 57756 454102
rect 57704 454038 57756 454044
rect 57612 454028 57664 454034
rect 57612 453970 57664 453976
rect 57336 435940 57388 435946
rect 57336 435882 57388 435888
rect 57716 390522 57744 454038
rect 57808 441614 57836 538047
rect 57888 533996 57940 534002
rect 57888 533938 57940 533944
rect 57900 533905 57928 533938
rect 57886 533896 57942 533905
rect 57886 533831 57942 533840
rect 58728 492658 58756 558826
rect 58716 492652 58768 492658
rect 58716 492594 58768 492600
rect 59004 462233 59032 561546
rect 59096 560250 59124 659738
rect 59176 638240 59228 638246
rect 59176 638182 59228 638188
rect 59084 560244 59136 560250
rect 59084 560186 59136 560192
rect 59188 536790 59216 638182
rect 59280 579630 59308 681838
rect 61936 666596 61988 666602
rect 61936 666538 61988 666544
rect 61844 663876 61896 663882
rect 61844 663818 61896 663824
rect 60648 661088 60700 661094
rect 60648 661030 60700 661036
rect 60372 635792 60424 635798
rect 60372 635734 60424 635740
rect 59268 579624 59320 579630
rect 59268 579566 59320 579572
rect 59280 578950 59308 579566
rect 59268 578944 59320 578950
rect 59268 578886 59320 578892
rect 60280 563236 60332 563242
rect 60280 563178 60332 563184
rect 60292 561610 60320 563178
rect 60280 561604 60332 561610
rect 60280 561546 60332 561552
rect 59268 560244 59320 560250
rect 59268 560186 59320 560192
rect 59280 559570 59308 560186
rect 59268 559564 59320 559570
rect 59268 559506 59320 559512
rect 59268 550588 59320 550594
rect 59268 550530 59320 550536
rect 59176 536784 59228 536790
rect 59176 536726 59228 536732
rect 59176 492652 59228 492658
rect 59176 492594 59228 492600
rect 59188 491570 59216 492594
rect 59176 491564 59228 491570
rect 59176 491506 59228 491512
rect 59084 463004 59136 463010
rect 59084 462946 59136 462952
rect 59096 462398 59124 462946
rect 59084 462392 59136 462398
rect 59084 462334 59136 462340
rect 58990 462224 59046 462233
rect 58990 462159 59046 462168
rect 58992 451308 59044 451314
rect 58992 451250 59044 451256
rect 58624 448588 58676 448594
rect 58624 448530 58676 448536
rect 57808 441586 57928 441614
rect 57900 438734 57928 441586
rect 57888 438728 57940 438734
rect 57888 438670 57940 438676
rect 57796 396840 57848 396846
rect 57796 396782 57848 396788
rect 57704 390516 57756 390522
rect 57704 390458 57756 390464
rect 57244 387252 57296 387258
rect 57244 387194 57296 387200
rect 57256 386578 57284 387194
rect 57244 386572 57296 386578
rect 57244 386514 57296 386520
rect 56508 355428 56560 355434
rect 56508 355370 56560 355376
rect 56416 336660 56468 336666
rect 56416 336602 56468 336608
rect 56520 329798 56548 355370
rect 56508 329792 56560 329798
rect 56508 329734 56560 329740
rect 56508 326528 56560 326534
rect 56508 326470 56560 326476
rect 56324 309188 56376 309194
rect 56324 309130 56376 309136
rect 56230 308408 56286 308417
rect 56230 308343 56286 308352
rect 55128 287020 55180 287026
rect 55128 286962 55180 286968
rect 56336 270502 56364 309130
rect 56416 303748 56468 303754
rect 56416 303690 56468 303696
rect 56324 270496 56376 270502
rect 56324 270438 56376 270444
rect 55864 264240 55916 264246
rect 55864 264182 55916 264188
rect 55876 263634 55904 264182
rect 56232 263696 56284 263702
rect 56232 263638 56284 263644
rect 55864 263628 55916 263634
rect 55864 263570 55916 263576
rect 55864 245540 55916 245546
rect 55864 245482 55916 245488
rect 55036 240100 55088 240106
rect 55036 240042 55088 240048
rect 54944 231736 54996 231742
rect 54944 231678 54996 231684
rect 55876 224874 55904 245482
rect 56244 235249 56272 263638
rect 56324 263628 56376 263634
rect 56324 263570 56376 263576
rect 56230 235240 56286 235249
rect 56230 235175 56286 235184
rect 56336 233238 56364 263570
rect 56428 260846 56456 303690
rect 56520 263566 56548 326470
rect 57256 297498 57284 386514
rect 57716 358086 57744 390458
rect 57808 387802 57836 396782
rect 57796 387796 57848 387802
rect 57796 387738 57848 387744
rect 57796 387252 57848 387258
rect 57796 387194 57848 387200
rect 57704 358080 57756 358086
rect 57704 358022 57756 358028
rect 57244 297492 57296 297498
rect 57244 297434 57296 297440
rect 57520 285728 57572 285734
rect 57520 285670 57572 285676
rect 56508 263560 56560 263566
rect 56508 263502 56560 263508
rect 56508 262268 56560 262274
rect 56508 262210 56560 262216
rect 56416 260840 56468 260846
rect 56416 260782 56468 260788
rect 56416 245676 56468 245682
rect 56416 245618 56468 245624
rect 56428 245546 56456 245618
rect 56416 245540 56468 245546
rect 56416 245482 56468 245488
rect 56324 233232 56376 233238
rect 56324 233174 56376 233180
rect 55864 224868 55916 224874
rect 55864 224810 55916 224816
rect 56520 213314 56548 262210
rect 56508 213308 56560 213314
rect 56508 213250 56560 213256
rect 57532 192545 57560 285670
rect 57716 271862 57744 358022
rect 57808 339425 57836 387194
rect 57794 339416 57850 339425
rect 57794 339351 57850 339360
rect 57900 337822 57928 438670
rect 58636 438462 58664 448530
rect 58624 438456 58676 438462
rect 58624 438398 58676 438404
rect 58624 387796 58676 387802
rect 58624 387738 58676 387744
rect 58636 340270 58664 387738
rect 59004 386374 59032 451250
rect 59096 391882 59124 462334
rect 59188 410582 59216 491506
rect 59280 448594 59308 550530
rect 60384 540258 60412 635734
rect 60554 584080 60610 584089
rect 60554 584015 60610 584024
rect 60464 567248 60516 567254
rect 60464 567190 60516 567196
rect 60096 540252 60148 540258
rect 60096 540194 60148 540200
rect 60372 540252 60424 540258
rect 60372 540194 60424 540200
rect 60108 539714 60136 540194
rect 60096 539708 60148 539714
rect 60096 539650 60148 539656
rect 60476 468518 60504 567190
rect 60568 563174 60596 584015
rect 60660 563242 60688 661030
rect 61752 641844 61804 641850
rect 61752 641786 61804 641792
rect 60648 563236 60700 563242
rect 60648 563178 60700 563184
rect 60556 563168 60608 563174
rect 60556 563110 60608 563116
rect 61384 563168 61436 563174
rect 61384 563110 61436 563116
rect 60648 563100 60700 563106
rect 60648 563042 60700 563048
rect 60660 547874 60688 563042
rect 60568 547846 60688 547874
rect 60464 468512 60516 468518
rect 60464 468454 60516 468460
rect 59268 448588 59320 448594
rect 59268 448530 59320 448536
rect 59176 410576 59228 410582
rect 59176 410518 59228 410524
rect 59084 391876 59136 391882
rect 59084 391818 59136 391824
rect 58992 386368 59044 386374
rect 58992 386310 59044 386316
rect 59096 367062 59124 391818
rect 60004 386368 60056 386374
rect 60004 386310 60056 386316
rect 59358 379536 59414 379545
rect 59280 379494 59358 379522
rect 59280 373994 59308 379494
rect 59358 379471 59414 379480
rect 59188 373966 59308 373994
rect 59084 367056 59136 367062
rect 59084 366998 59136 367004
rect 59084 344344 59136 344350
rect 59084 344286 59136 344292
rect 59096 343670 59124 344286
rect 59084 343664 59136 343670
rect 59084 343606 59136 343612
rect 58624 340264 58676 340270
rect 58624 340206 58676 340212
rect 57888 337816 57940 337822
rect 57888 337758 57940 337764
rect 57796 327820 57848 327826
rect 57796 327762 57848 327768
rect 57808 285666 57836 327762
rect 57796 285660 57848 285666
rect 57796 285602 57848 285608
rect 57796 279472 57848 279478
rect 57796 279414 57848 279420
rect 57808 278905 57836 279414
rect 57794 278896 57850 278905
rect 57794 278831 57850 278840
rect 57704 271856 57756 271862
rect 57704 271798 57756 271804
rect 57704 269816 57756 269822
rect 57704 269758 57756 269764
rect 57612 249076 57664 249082
rect 57612 249018 57664 249024
rect 57624 248538 57652 249018
rect 57612 248532 57664 248538
rect 57612 248474 57664 248480
rect 57624 216578 57652 248474
rect 57612 216572 57664 216578
rect 57612 216514 57664 216520
rect 57518 192536 57574 192545
rect 57518 192471 57574 192480
rect 57716 182850 57744 269758
rect 57900 237386 57928 337758
rect 59096 336054 59124 343606
rect 59084 336048 59136 336054
rect 59084 335990 59136 335996
rect 59084 289876 59136 289882
rect 59084 289818 59136 289824
rect 58900 240780 58952 240786
rect 58900 240722 58952 240728
rect 57888 237380 57940 237386
rect 57888 237322 57940 237328
rect 58912 235754 58940 240722
rect 58900 235748 58952 235754
rect 58900 235690 58952 235696
rect 59096 228478 59124 289818
rect 59084 228472 59136 228478
rect 59084 228414 59136 228420
rect 57704 182844 57756 182850
rect 57704 182786 57756 182792
rect 57796 127016 57848 127022
rect 57796 126958 57848 126964
rect 56508 122868 56560 122874
rect 56508 122810 56560 122816
rect 56520 91050 56548 122810
rect 57808 93809 57836 126958
rect 57888 120148 57940 120154
rect 57888 120090 57940 120096
rect 57794 93800 57850 93809
rect 57794 93735 57850 93744
rect 56508 91044 56560 91050
rect 56508 90986 56560 90992
rect 57900 74526 57928 120090
rect 57888 74520 57940 74526
rect 57888 74462 57940 74468
rect 54760 69760 54812 69766
rect 54760 69702 54812 69708
rect 55220 69692 55272 69698
rect 55220 69634 55272 69640
rect 55232 16574 55260 69634
rect 59188 64258 59216 373966
rect 59268 372632 59320 372638
rect 59268 372574 59320 372580
rect 59176 64252 59228 64258
rect 59176 64194 59228 64200
rect 56600 60036 56652 60042
rect 56600 59978 56652 59984
rect 56612 16574 56640 59978
rect 59280 28966 59308 372574
rect 60016 353258 60044 386310
rect 60476 373998 60504 468454
rect 60568 464438 60596 547846
rect 60740 546508 60792 546514
rect 60740 546450 60792 546456
rect 60752 546417 60780 546450
rect 60738 546408 60794 546417
rect 60738 546343 60794 546352
rect 60648 543720 60700 543726
rect 60648 543662 60700 543668
rect 60556 464432 60608 464438
rect 60556 464374 60608 464380
rect 60464 373992 60516 373998
rect 60464 373934 60516 373940
rect 60476 372638 60504 373934
rect 60464 372632 60516 372638
rect 60464 372574 60516 372580
rect 60372 369164 60424 369170
rect 60372 369106 60424 369112
rect 60004 353252 60056 353258
rect 60004 353194 60056 353200
rect 60384 339386 60412 369106
rect 60568 367169 60596 464374
rect 60660 442950 60688 543662
rect 60740 543040 60792 543046
rect 60738 543008 60740 543017
rect 60792 543008 60794 543017
rect 60738 542943 60794 542952
rect 61396 538801 61424 563110
rect 61764 543726 61792 641786
rect 61856 564262 61884 663818
rect 61948 566506 61976 666538
rect 62040 663066 62068 700266
rect 68928 690668 68980 690674
rect 68928 690610 68980 690616
rect 68652 687948 68704 687954
rect 68652 687890 68704 687896
rect 67546 679144 67602 679153
rect 67546 679079 67602 679088
rect 64696 677612 64748 677618
rect 64696 677554 64748 677560
rect 63224 670744 63276 670750
rect 63224 670686 63276 670692
rect 62028 663060 62080 663066
rect 62028 663002 62080 663008
rect 62040 661706 62068 663002
rect 62028 661700 62080 661706
rect 62028 661642 62080 661648
rect 63132 647352 63184 647358
rect 63132 647294 63184 647300
rect 62028 647284 62080 647290
rect 62028 647226 62080 647232
rect 61936 566500 61988 566506
rect 61936 566442 61988 566448
rect 61844 564256 61896 564262
rect 61844 564198 61896 564204
rect 61856 563106 61884 564198
rect 61844 563100 61896 563106
rect 61844 563042 61896 563048
rect 61752 543720 61804 543726
rect 61752 543662 61804 543668
rect 61382 538792 61438 538801
rect 61382 538727 61438 538736
rect 61844 480208 61896 480214
rect 61844 480150 61896 480156
rect 61752 477556 61804 477562
rect 61752 477498 61804 477504
rect 61382 463584 61438 463593
rect 61382 463519 61438 463528
rect 61396 462369 61424 463519
rect 61382 462360 61438 462369
rect 61382 462295 61438 462304
rect 60648 442944 60700 442950
rect 60648 442886 60700 442892
rect 60648 384532 60700 384538
rect 60648 384474 60700 384480
rect 60554 367160 60610 367169
rect 60554 367095 60610 367104
rect 60462 356688 60518 356697
rect 60462 356623 60518 356632
rect 60372 339380 60424 339386
rect 60372 339322 60424 339328
rect 60476 333810 60504 356623
rect 60464 333804 60516 333810
rect 60464 333746 60516 333752
rect 60556 330540 60608 330546
rect 60556 330482 60608 330488
rect 60372 288448 60424 288454
rect 60372 288390 60424 288396
rect 60384 238134 60412 288390
rect 60568 286958 60596 330482
rect 60556 286952 60608 286958
rect 60556 286894 60608 286900
rect 60464 247104 60516 247110
rect 60464 247046 60516 247052
rect 60372 238128 60424 238134
rect 60372 238070 60424 238076
rect 60476 222902 60504 247046
rect 60464 222896 60516 222902
rect 60464 222838 60516 222844
rect 60660 69018 60688 384474
rect 61396 367033 61424 462295
rect 61764 385014 61792 477498
rect 61856 447273 61884 480150
rect 61948 467838 61976 566442
rect 62040 546650 62068 647226
rect 62120 554736 62172 554742
rect 62120 554678 62172 554684
rect 62028 546644 62080 546650
rect 62028 546586 62080 546592
rect 62028 540932 62080 540938
rect 62028 540874 62080 540880
rect 61936 467832 61988 467838
rect 61936 467774 61988 467780
rect 61936 448520 61988 448526
rect 61936 448462 61988 448468
rect 61842 447264 61898 447273
rect 61842 447199 61898 447208
rect 61844 440292 61896 440298
rect 61844 440234 61896 440240
rect 61752 385008 61804 385014
rect 61752 384950 61804 384956
rect 61764 384538 61792 384950
rect 61752 384532 61804 384538
rect 61752 384474 61804 384480
rect 61382 367024 61438 367033
rect 61382 366959 61438 366968
rect 61660 351892 61712 351898
rect 61660 351834 61712 351840
rect 60740 72480 60792 72486
rect 60740 72422 60792 72428
rect 60648 69012 60700 69018
rect 60648 68954 60700 68960
rect 59358 57216 59414 57225
rect 59358 57151 59414 57160
rect 59268 28960 59320 28966
rect 59268 28902 59320 28908
rect 53852 16546 54984 16574
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 53380 3392 53432 3398
rect 53380 3334 53432 3340
rect 51326 354 51438 480
rect 51092 326 51438 354
rect 51326 -960 51438 326
rect 52522 -960 52634 480
rect 53392 354 53420 3334
rect 54956 480 54984 16546
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58440 13116 58492 13122
rect 58440 13058 58492 13064
rect 58452 480 58480 13058
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 57151
rect 60752 6914 60780 72422
rect 61672 65618 61700 351834
rect 61856 339590 61884 440234
rect 61948 349178 61976 448462
rect 62040 440910 62068 540874
rect 62132 456754 62160 554678
rect 63144 549234 63172 647294
rect 63236 571266 63264 670686
rect 64512 669384 64564 669390
rect 64512 669326 64564 669332
rect 63408 658300 63460 658306
rect 63408 658242 63460 658248
rect 63316 640416 63368 640422
rect 63316 640358 63368 640364
rect 63224 571260 63276 571266
rect 63224 571202 63276 571208
rect 63224 568676 63276 568682
rect 63224 568618 63276 568624
rect 63132 549228 63184 549234
rect 63132 549170 63184 549176
rect 63236 480254 63264 568618
rect 63328 540938 63356 640358
rect 63420 558890 63448 658242
rect 64524 571334 64552 669326
rect 64604 648644 64656 648650
rect 64604 648586 64656 648592
rect 64512 571328 64564 571334
rect 64512 571270 64564 571276
rect 63500 564392 63552 564398
rect 63500 564334 63552 564340
rect 63408 558884 63460 558890
rect 63408 558826 63460 558832
rect 63408 549228 63460 549234
rect 63408 549170 63460 549176
rect 63420 548622 63448 549170
rect 63408 548616 63460 548622
rect 63408 548558 63460 548564
rect 63316 540932 63368 540938
rect 63316 540874 63368 540880
rect 63236 480226 63356 480254
rect 63038 477592 63094 477601
rect 63038 477527 63040 477536
rect 63092 477527 63094 477536
rect 63040 477498 63092 477504
rect 63328 470218 63356 480226
rect 63316 470212 63368 470218
rect 63316 470154 63368 470160
rect 62764 466404 62816 466410
rect 62764 466346 62816 466352
rect 62120 456748 62172 456754
rect 62120 456690 62172 456696
rect 62132 456074 62160 456690
rect 62120 456068 62172 456074
rect 62120 456010 62172 456016
rect 62028 440904 62080 440910
rect 62028 440846 62080 440852
rect 62040 440298 62068 440846
rect 62028 440292 62080 440298
rect 62028 440234 62080 440240
rect 62028 375420 62080 375426
rect 62028 375362 62080 375368
rect 61936 349172 61988 349178
rect 61936 349114 61988 349120
rect 61844 339584 61896 339590
rect 61844 339526 61896 339532
rect 61844 291848 61896 291854
rect 61844 291790 61896 291796
rect 61856 276690 61884 291790
rect 61844 276684 61896 276690
rect 61844 276626 61896 276632
rect 61844 258120 61896 258126
rect 61844 258062 61896 258068
rect 61752 251252 61804 251258
rect 61752 251194 61804 251200
rect 61764 234598 61792 251194
rect 61752 234592 61804 234598
rect 61752 234534 61804 234540
rect 61856 229906 61884 258062
rect 61844 229900 61896 229906
rect 61844 229842 61896 229848
rect 61660 65612 61712 65618
rect 61660 65554 61712 65560
rect 62040 46238 62068 375362
rect 62776 369850 62804 466346
rect 63130 446040 63186 446049
rect 63130 445975 63186 445984
rect 63144 445806 63172 445975
rect 63132 445800 63184 445806
rect 63132 445742 63184 445748
rect 63144 441614 63172 445742
rect 63144 441586 63264 441614
rect 62764 369844 62816 369850
rect 62764 369786 62816 369792
rect 63132 349036 63184 349042
rect 63132 348978 63184 348984
rect 62028 46232 62080 46238
rect 62028 46174 62080 46180
rect 60832 18692 60884 18698
rect 60832 18634 60884 18640
rect 60844 16574 60872 18634
rect 60844 16546 61608 16574
rect 60752 6886 60872 6914
rect 60844 480 60872 6886
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61580 354 61608 16546
rect 63040 10396 63092 10402
rect 63040 10338 63092 10344
rect 63052 3482 63080 10338
rect 63144 5506 63172 348978
rect 63236 347750 63264 441586
rect 63328 374678 63356 470154
rect 63420 448526 63448 548558
rect 63512 466410 63540 564334
rect 64144 558884 64196 558890
rect 64144 558826 64196 558832
rect 64156 557666 64184 558826
rect 64144 557660 64196 557666
rect 64144 557602 64196 557608
rect 63500 466404 63552 466410
rect 63500 466346 63552 466352
rect 64156 459542 64184 557602
rect 64616 550594 64644 648586
rect 64708 578241 64736 677554
rect 67454 675744 67510 675753
rect 67454 675679 67510 675688
rect 66076 673736 66128 673742
rect 66076 673678 66128 673684
rect 65892 670812 65944 670818
rect 65892 670754 65944 670760
rect 64788 651432 64840 651438
rect 64788 651374 64840 651380
rect 64694 578232 64750 578241
rect 64694 578167 64750 578176
rect 64800 552022 64828 651374
rect 65904 571810 65932 670754
rect 65984 666664 66036 666670
rect 65984 666606 66036 666612
rect 65892 571804 65944 571810
rect 65892 571746 65944 571752
rect 65892 571328 65944 571334
rect 65892 571270 65944 571276
rect 64788 552016 64840 552022
rect 64788 551958 64840 551964
rect 65616 552016 65668 552022
rect 65616 551958 65668 551964
rect 64604 550588 64656 550594
rect 64604 550530 64656 550536
rect 64788 546644 64840 546650
rect 64788 546586 64840 546592
rect 64696 484424 64748 484430
rect 64696 484366 64748 484372
rect 64234 468480 64290 468489
rect 64234 468415 64290 468424
rect 64248 467974 64276 468415
rect 64236 467968 64288 467974
rect 64234 467936 64236 467945
rect 64288 467936 64290 467945
rect 64234 467871 64290 467880
rect 63500 459536 63552 459542
rect 63500 459478 63552 459484
rect 64144 459536 64196 459542
rect 64144 459478 64196 459484
rect 63512 458862 63540 459478
rect 63500 458856 63552 458862
rect 63500 458798 63552 458804
rect 64144 448588 64196 448594
rect 64144 448530 64196 448536
rect 63408 448520 63460 448526
rect 63408 448462 63460 448468
rect 63408 441584 63460 441590
rect 63408 441526 63460 441532
rect 63316 374672 63368 374678
rect 63316 374614 63368 374620
rect 63224 347744 63276 347750
rect 63224 347686 63276 347692
rect 63224 270564 63276 270570
rect 63224 270506 63276 270512
rect 63236 237289 63264 270506
rect 63222 237280 63278 237289
rect 63222 237215 63278 237224
rect 63328 206378 63356 374614
rect 63420 340950 63448 441526
rect 64156 351898 64184 448530
rect 64604 442944 64656 442950
rect 64604 442886 64656 442892
rect 64616 441658 64644 442886
rect 64604 441652 64656 441658
rect 64604 441594 64656 441600
rect 64510 364440 64566 364449
rect 64510 364375 64566 364384
rect 64144 351892 64196 351898
rect 64144 351834 64196 351840
rect 63408 340944 63460 340950
rect 63408 340886 63460 340892
rect 63316 206372 63368 206378
rect 63316 206314 63368 206320
rect 64524 27606 64552 364375
rect 64616 342310 64644 441594
rect 64708 439618 64736 484366
rect 64800 447166 64828 546586
rect 65524 541680 65576 541686
rect 65524 541622 65576 541628
rect 64788 447160 64840 447166
rect 64788 447102 64840 447108
rect 65536 441522 65564 541622
rect 65628 452606 65656 551958
rect 65904 471102 65932 571270
rect 65996 568274 66024 666606
rect 66088 574025 66116 673678
rect 66168 669452 66220 669458
rect 66168 669394 66220 669400
rect 66074 574016 66130 574025
rect 66074 573951 66130 573960
rect 66076 571804 66128 571810
rect 66076 571746 66128 571752
rect 65984 568268 66036 568274
rect 65984 568210 66036 568216
rect 65996 567254 66024 568210
rect 65984 567248 66036 567254
rect 65984 567190 66036 567196
rect 65982 546136 66038 546145
rect 65982 546071 66038 546080
rect 65996 545154 66024 546071
rect 65984 545148 66036 545154
rect 65984 545090 66036 545096
rect 66088 473346 66116 571746
rect 66180 569906 66208 669394
rect 67364 667956 67416 667962
rect 67364 667898 67416 667904
rect 66168 569900 66220 569906
rect 66168 569842 66220 569848
rect 66996 569900 67048 569906
rect 66996 569842 67048 569848
rect 67008 568954 67036 569842
rect 66996 568948 67048 568954
rect 66996 568890 67048 568896
rect 66904 565140 66956 565146
rect 66904 565082 66956 565088
rect 66260 480888 66312 480894
rect 66260 480830 66312 480836
rect 66272 479534 66300 480830
rect 66260 479528 66312 479534
rect 66260 479470 66312 479476
rect 66076 473340 66128 473346
rect 66076 473282 66128 473288
rect 66088 472666 66116 473282
rect 66076 472660 66128 472666
rect 66076 472602 66128 472608
rect 65892 471096 65944 471102
rect 65892 471038 65944 471044
rect 66168 470484 66220 470490
rect 66168 470426 66220 470432
rect 65616 452600 65668 452606
rect 65616 452542 65668 452548
rect 65628 451314 65656 452542
rect 65616 451308 65668 451314
rect 65616 451250 65668 451256
rect 65616 447160 65668 447166
rect 65616 447102 65668 447108
rect 65524 441516 65576 441522
rect 65524 441458 65576 441464
rect 64696 439612 64748 439618
rect 64696 439554 64748 439560
rect 64786 401704 64842 401713
rect 64786 401639 64788 401648
rect 64840 401639 64842 401648
rect 64788 401610 64840 401616
rect 64696 394732 64748 394738
rect 64696 394674 64748 394680
rect 64708 362914 64736 394674
rect 64800 373318 64828 401610
rect 65524 376780 65576 376786
rect 65524 376722 65576 376728
rect 64788 373312 64840 373318
rect 64788 373254 64840 373260
rect 64696 362908 64748 362914
rect 64696 362850 64748 362856
rect 64696 349172 64748 349178
rect 64696 349114 64748 349120
rect 64604 342304 64656 342310
rect 64604 342246 64656 342252
rect 64604 339584 64656 339590
rect 64604 339526 64656 339532
rect 64616 73166 64644 339526
rect 64604 73160 64656 73166
rect 64604 73102 64656 73108
rect 64708 49706 64736 349114
rect 65536 299470 65564 376722
rect 65628 349042 65656 447102
rect 66180 404433 66208 470426
rect 66916 465730 66944 565082
rect 67008 470490 67036 568890
rect 67376 568682 67404 667898
rect 67468 575249 67496 675679
rect 67560 577810 67588 679079
rect 67638 678192 67694 678201
rect 67638 678127 67694 678136
rect 67652 677618 67680 678127
rect 67640 677612 67692 677618
rect 67640 677554 67692 677560
rect 67638 676424 67694 676433
rect 67638 676359 67694 676368
rect 67652 676258 67680 676359
rect 67640 676252 67692 676258
rect 67640 676194 67692 676200
rect 67638 675200 67694 675209
rect 67638 675135 67694 675144
rect 67652 674966 67680 675135
rect 67640 674960 67692 674966
rect 67640 674902 67692 674908
rect 67638 674384 67694 674393
rect 67638 674319 67694 674328
rect 67652 673538 67680 674319
rect 67730 673840 67786 673849
rect 67730 673775 67786 673784
rect 67744 673742 67772 673775
rect 67732 673736 67784 673742
rect 67732 673678 67784 673684
rect 67640 673532 67692 673538
rect 67640 673474 67692 673480
rect 68664 671809 68692 687890
rect 68836 685160 68888 685166
rect 68836 685102 68888 685108
rect 68742 677104 68798 677113
rect 68742 677039 68798 677048
rect 68650 671800 68706 671809
rect 68650 671735 68706 671744
rect 67638 670984 67694 670993
rect 67638 670919 67694 670928
rect 67652 670750 67680 670919
rect 68664 670818 68692 671735
rect 68652 670812 68704 670818
rect 68652 670754 68704 670760
rect 67640 670744 67692 670750
rect 67640 670686 67692 670692
rect 67638 670304 67694 670313
rect 67638 670239 67694 670248
rect 67652 669390 67680 670239
rect 67730 669624 67786 669633
rect 67730 669559 67786 669568
rect 67640 669384 67692 669390
rect 67640 669326 67692 669332
rect 67744 667962 67772 669559
rect 67824 669452 67876 669458
rect 67824 669394 67876 669400
rect 67836 669361 67864 669394
rect 67822 669352 67878 669361
rect 67822 669287 67878 669296
rect 67822 668264 67878 668273
rect 67822 668199 67878 668208
rect 67732 667956 67784 667962
rect 67732 667898 67784 667904
rect 67638 666904 67694 666913
rect 67638 666839 67694 666848
rect 67652 666602 67680 666839
rect 67836 666670 67864 668199
rect 67824 666664 67876 666670
rect 67824 666606 67876 666612
rect 67640 666596 67692 666602
rect 67640 666538 67692 666544
rect 68560 666596 68612 666602
rect 68560 666538 68612 666544
rect 67730 665544 67786 665553
rect 67730 665479 67786 665488
rect 67744 665310 67772 665479
rect 67732 665304 67784 665310
rect 67638 665272 67694 665281
rect 67732 665246 67784 665252
rect 67638 665207 67640 665216
rect 67692 665207 67694 665216
rect 67640 665178 67692 665184
rect 67730 664184 67786 664193
rect 67730 664119 67786 664128
rect 67638 663912 67694 663921
rect 67638 663847 67640 663856
rect 67692 663847 67694 663856
rect 67640 663818 67692 663824
rect 67744 663814 67772 664119
rect 67732 663808 67784 663814
rect 67732 663750 67784 663756
rect 67640 663060 67692 663066
rect 67640 663002 67692 663008
rect 67652 662969 67680 663002
rect 67638 662960 67694 662969
rect 67638 662895 67694 662904
rect 67638 661464 67694 661473
rect 67638 661399 67694 661408
rect 67652 661094 67680 661399
rect 67640 661088 67692 661094
rect 67640 661030 67692 661036
rect 67730 660104 67786 660113
rect 67730 660039 67786 660048
rect 67640 659796 67692 659802
rect 67640 659738 67692 659744
rect 67652 659705 67680 659738
rect 67744 659734 67772 660039
rect 67732 659728 67784 659734
rect 67638 659696 67694 659705
rect 67732 659670 67784 659676
rect 67638 659631 67694 659640
rect 68572 658986 68600 666538
rect 68560 658980 68612 658986
rect 68560 658922 68612 658928
rect 68572 658889 68600 658922
rect 68558 658880 68614 658889
rect 68558 658815 68614 658824
rect 67638 658744 67694 658753
rect 67638 658679 67694 658688
rect 67652 658306 67680 658679
rect 67640 658300 67692 658306
rect 67640 658242 67692 658248
rect 67730 657384 67786 657393
rect 67730 657319 67786 657328
rect 67744 656946 67772 657319
rect 68192 657008 68244 657014
rect 68192 656950 68244 656956
rect 67732 656940 67784 656946
rect 67732 656882 67784 656888
rect 68204 656713 68232 656950
rect 68190 656704 68246 656713
rect 68190 656639 68246 656648
rect 67638 656024 67694 656033
rect 67638 655959 67694 655968
rect 67652 655586 67680 655959
rect 67640 655580 67692 655586
rect 67640 655522 67692 655528
rect 67640 654832 67692 654838
rect 67638 654800 67640 654809
rect 67692 654800 67694 654809
rect 67638 654735 67694 654744
rect 67730 653304 67786 653313
rect 67730 653239 67786 653248
rect 67744 652798 67772 653239
rect 67916 652860 67968 652866
rect 67916 652802 67968 652808
rect 67732 652792 67784 652798
rect 67928 652769 67956 652802
rect 67732 652734 67784 652740
rect 67914 652760 67970 652769
rect 67914 652695 67970 652704
rect 67638 651944 67694 651953
rect 67638 651879 67694 651888
rect 67652 651438 67680 651879
rect 67640 651432 67692 651438
rect 67640 651374 67692 651380
rect 67640 650072 67692 650078
rect 67638 650040 67640 650049
rect 67692 650040 67694 650049
rect 67638 649975 67694 649984
rect 67638 649224 67694 649233
rect 67638 649159 67694 649168
rect 67652 648650 67680 649159
rect 67640 648644 67692 648650
rect 67640 648586 67692 648592
rect 67730 647864 67786 647873
rect 67730 647799 67786 647808
rect 67744 647358 67772 647799
rect 67732 647352 67784 647358
rect 67638 647320 67694 647329
rect 67732 647294 67784 647300
rect 67638 647255 67640 647264
rect 67692 647255 67694 647264
rect 67640 647226 67692 647232
rect 67638 646504 67694 646513
rect 67638 646439 67694 646448
rect 67652 645930 67680 646439
rect 67640 645924 67692 645930
rect 67640 645866 67692 645872
rect 68558 643784 68614 643793
rect 68558 643719 68614 643728
rect 67730 642424 67786 642433
rect 67730 642359 67786 642368
rect 67638 641880 67694 641889
rect 67744 641850 67772 642359
rect 67638 641815 67694 641824
rect 67732 641844 67784 641850
rect 67652 641782 67680 641815
rect 67732 641786 67784 641792
rect 67640 641776 67692 641782
rect 67640 641718 67692 641724
rect 67730 641064 67786 641073
rect 67730 640999 67786 641008
rect 67638 640520 67694 640529
rect 67638 640455 67694 640464
rect 67652 640422 67680 640455
rect 67640 640416 67692 640422
rect 67640 640358 67692 640364
rect 67744 640354 67772 640999
rect 67732 640348 67784 640354
rect 67732 640290 67784 640296
rect 67640 579624 67692 579630
rect 67640 579566 67692 579572
rect 67652 579329 67680 579566
rect 67638 579320 67694 579329
rect 67638 579255 67694 579264
rect 67730 578232 67786 578241
rect 67730 578167 67786 578176
rect 67638 577824 67694 577833
rect 67560 577782 67638 577810
rect 67454 575240 67510 575249
rect 67454 575175 67510 575184
rect 67364 568676 67416 568682
rect 67364 568618 67416 568624
rect 67560 480214 67588 577782
rect 67638 577759 67694 577768
rect 67744 577289 67772 578167
rect 67730 577280 67786 577289
rect 67730 577215 67786 577224
rect 67638 575784 67694 575793
rect 67638 575719 67694 575728
rect 67652 575550 67680 575719
rect 67640 575544 67692 575550
rect 67640 575486 67692 575492
rect 67640 574796 67692 574802
rect 67640 574738 67692 574744
rect 67652 574569 67680 574738
rect 67638 574560 67694 574569
rect 67638 574495 67694 574504
rect 67640 574048 67692 574054
rect 67640 573990 67692 573996
rect 67730 574016 67786 574025
rect 67652 573889 67680 573990
rect 67730 573951 67786 573960
rect 67638 573880 67694 573889
rect 67638 573815 67694 573824
rect 67744 573345 67772 573951
rect 67730 573336 67786 573345
rect 67730 573271 67786 573280
rect 67640 571804 67692 571810
rect 67640 571746 67692 571752
rect 67652 571713 67680 571746
rect 67638 571704 67694 571713
rect 67638 571639 67694 571648
rect 67732 571328 67784 571334
rect 67732 571270 67784 571276
rect 67640 571260 67692 571266
rect 67640 571202 67692 571208
rect 67652 571033 67680 571202
rect 67638 571024 67694 571033
rect 67638 570959 67694 570968
rect 67744 570353 67772 571270
rect 67730 570344 67786 570353
rect 67730 570279 67786 570288
rect 67638 569120 67694 569129
rect 67638 569055 67694 569064
rect 67652 568682 67680 569055
rect 67822 568984 67878 568993
rect 67822 568919 67824 568928
rect 67876 568919 67878 568928
rect 67824 568890 67876 568896
rect 67640 568676 67692 568682
rect 67640 568618 67692 568624
rect 67638 568304 67694 568313
rect 67638 568239 67640 568248
rect 67692 568239 67694 568248
rect 67640 568210 67692 568216
rect 67640 567860 67692 567866
rect 67640 567802 67692 567808
rect 67652 567769 67680 567802
rect 67638 567760 67694 567769
rect 67638 567695 67694 567704
rect 67640 566500 67692 566506
rect 67640 566442 67692 566448
rect 67652 566409 67680 566442
rect 67638 566400 67694 566409
rect 67638 566335 67694 566344
rect 67640 565140 67692 565146
rect 67640 565082 67692 565088
rect 67652 565049 67680 565082
rect 67638 565040 67694 565049
rect 67638 564975 67694 564984
rect 67638 564904 67694 564913
rect 67638 564839 67694 564848
rect 67652 564466 67680 564839
rect 67640 564460 67692 564466
rect 67640 564402 67692 564408
rect 67640 564324 67692 564330
rect 67640 564266 67692 564272
rect 67652 564233 67680 564266
rect 67732 564256 67784 564262
rect 67638 564224 67694 564233
rect 67732 564198 67784 564204
rect 67638 564159 67694 564168
rect 67744 563689 67772 564198
rect 67730 563680 67786 563689
rect 67730 563615 67786 563624
rect 67640 562352 67692 562358
rect 67638 562320 67640 562329
rect 67692 562320 67694 562329
rect 67638 562255 67694 562264
rect 67732 561672 67784 561678
rect 67732 561614 67784 561620
rect 67640 561604 67692 561610
rect 67640 561546 67692 561552
rect 67652 561513 67680 561546
rect 67638 561504 67694 561513
rect 67638 561439 67694 561448
rect 67744 560969 67772 561614
rect 67730 560960 67786 560969
rect 67730 560895 67786 560904
rect 67640 560244 67692 560250
rect 67640 560186 67692 560192
rect 67652 559609 67680 560186
rect 67638 559600 67694 559609
rect 67638 559535 67694 559544
rect 67730 558104 67786 558113
rect 67730 558039 67786 558048
rect 67640 557660 67692 557666
rect 67640 557602 67692 557608
rect 67652 557569 67680 557602
rect 67744 557598 67772 558039
rect 67732 557592 67784 557598
rect 67638 557560 67694 557569
rect 67732 557534 67784 557540
rect 67638 557495 67694 557504
rect 67824 557524 67876 557530
rect 67824 557466 67876 557472
rect 67640 557456 67692 557462
rect 67836 557433 67864 557466
rect 67640 557398 67692 557404
rect 67822 557424 67878 557433
rect 67652 556889 67680 557398
rect 67822 557359 67878 557368
rect 67638 556880 67694 556889
rect 67638 556815 67694 556824
rect 67732 556164 67784 556170
rect 67732 556106 67784 556112
rect 67638 555384 67694 555393
rect 67638 555319 67694 555328
rect 67652 554810 67680 555319
rect 67744 554849 67772 556106
rect 67730 554840 67786 554849
rect 67640 554804 67692 554810
rect 67730 554775 67786 554784
rect 67640 554746 67692 554752
rect 67914 554704 67970 554713
rect 67640 554668 67692 554674
rect 67914 554639 67970 554648
rect 67640 554610 67692 554616
rect 67652 554169 67680 554610
rect 67638 554160 67694 554169
rect 67638 554095 67694 554104
rect 67928 553450 67956 554639
rect 67916 553444 67968 553450
rect 67916 553386 67968 553392
rect 67640 552696 67692 552702
rect 67638 552664 67640 552673
rect 67692 552664 67694 552673
rect 67638 552599 67694 552608
rect 67640 552016 67692 552022
rect 67638 551984 67640 551993
rect 67692 551984 67694 551993
rect 67638 551919 67694 551928
rect 67640 550588 67692 550594
rect 67640 550530 67692 550536
rect 67652 549409 67680 550530
rect 67638 549400 67694 549409
rect 67638 549335 67694 549344
rect 67730 549264 67786 549273
rect 67730 549199 67786 549208
rect 67640 548616 67692 548622
rect 67638 548584 67640 548593
rect 67692 548584 67694 548593
rect 67638 548519 67694 548528
rect 67744 547942 67772 549199
rect 67732 547936 67784 547942
rect 67732 547878 67784 547884
rect 67638 547224 67694 547233
rect 67638 547159 67694 547168
rect 67652 546650 67680 547159
rect 67640 546644 67692 546650
rect 67640 546586 67692 546592
rect 67638 546544 67694 546553
rect 67638 546479 67640 546488
rect 67692 546479 67694 546488
rect 67640 546450 67692 546456
rect 67638 545184 67694 545193
rect 67638 545119 67640 545128
rect 67692 545119 67694 545128
rect 67640 545090 67692 545096
rect 68572 545086 68600 643719
rect 68756 576854 68784 677039
rect 68848 666602 68876 685102
rect 68836 666596 68888 666602
rect 68836 666538 68888 666544
rect 68940 654809 68968 690610
rect 69112 680400 69164 680406
rect 69112 680342 69164 680348
rect 68926 654800 68982 654809
rect 68926 654735 68982 654744
rect 68834 651400 68890 651409
rect 68834 651335 68890 651344
rect 68664 576826 68784 576854
rect 68664 576609 68692 576826
rect 68650 576600 68706 576609
rect 68650 576535 68706 576544
rect 68560 545080 68612 545086
rect 68560 545022 68612 545028
rect 68572 543833 68600 545022
rect 68190 543824 68246 543833
rect 68190 543759 68246 543768
rect 68558 543824 68614 543833
rect 68558 543759 68614 543768
rect 67732 543720 67784 543726
rect 67732 543662 67784 543668
rect 67638 543280 67694 543289
rect 67638 543215 67694 543224
rect 67652 543046 67680 543215
rect 67744 543153 67772 543662
rect 67730 543144 67786 543153
rect 67730 543079 67786 543088
rect 67640 543040 67692 543046
rect 67640 542982 67692 542988
rect 67640 541680 67692 541686
rect 67640 541622 67692 541628
rect 67652 541249 67680 541622
rect 67638 541240 67694 541249
rect 67638 541175 67694 541184
rect 67640 540932 67692 540938
rect 67640 540874 67692 540880
rect 67652 540569 67680 540874
rect 67638 540560 67694 540569
rect 67638 540495 67694 540504
rect 67730 489152 67786 489161
rect 67730 489087 67786 489096
rect 67744 488578 67772 489087
rect 67732 488572 67784 488578
rect 67732 488514 67784 488520
rect 67640 488504 67692 488510
rect 67640 488446 67692 488452
rect 67652 488073 67680 488446
rect 67638 488064 67694 488073
rect 67638 487999 67694 488008
rect 67638 487928 67694 487937
rect 67638 487863 67694 487872
rect 67652 487830 67680 487863
rect 67640 487824 67692 487830
rect 67640 487766 67692 487772
rect 67730 486568 67786 486577
rect 67730 486503 67786 486512
rect 67744 485926 67772 486503
rect 67732 485920 67784 485926
rect 67638 485888 67694 485897
rect 67732 485862 67784 485868
rect 67638 485823 67640 485832
rect 67692 485823 67694 485832
rect 67640 485794 67692 485800
rect 67638 485208 67694 485217
rect 67638 485143 67694 485152
rect 67652 485110 67680 485143
rect 67640 485104 67692 485110
rect 67640 485046 67692 485052
rect 67638 483984 67694 483993
rect 67638 483919 67694 483928
rect 67652 483682 67680 483919
rect 67640 483676 67692 483682
rect 67640 483618 67692 483624
rect 68008 482996 68060 483002
rect 68008 482938 68060 482944
rect 68020 482497 68048 482938
rect 68006 482488 68062 482497
rect 68006 482423 68062 482432
rect 68098 481536 68154 481545
rect 68098 481471 68154 481480
rect 67638 481128 67694 481137
rect 67638 481063 67694 481072
rect 67652 480894 67680 481063
rect 67640 480888 67692 480894
rect 67640 480830 67692 480836
rect 68112 480593 68140 481471
rect 68098 480584 68154 480593
rect 68098 480519 68154 480528
rect 67548 480208 67600 480214
rect 67548 480150 67600 480156
rect 67560 479233 67588 480150
rect 67638 479768 67694 479777
rect 67638 479703 67694 479712
rect 67546 479224 67602 479233
rect 67546 479159 67602 479168
rect 67652 478922 67680 479703
rect 67640 478916 67692 478922
rect 67640 478858 67692 478864
rect 67638 478272 67694 478281
rect 67638 478207 67694 478216
rect 67652 477562 67680 478207
rect 67640 477556 67692 477562
rect 67640 477498 67692 477504
rect 67638 476504 67694 476513
rect 67638 476439 67694 476448
rect 67652 476134 67680 476439
rect 67640 476128 67692 476134
rect 67640 476070 67692 476076
rect 67638 475688 67694 475697
rect 67638 475623 67694 475632
rect 67652 475454 67680 475623
rect 67640 475448 67692 475454
rect 67640 475390 67692 475396
rect 67732 475380 67784 475386
rect 67732 475322 67784 475328
rect 67744 475017 67772 475322
rect 67730 475008 67786 475017
rect 67560 474966 67730 474994
rect 67088 471096 67140 471102
rect 67088 471038 67140 471044
rect 66996 470484 67048 470490
rect 66996 470426 67048 470432
rect 66904 465724 66956 465730
rect 66904 465666 66956 465672
rect 66166 404424 66222 404433
rect 66166 404359 66222 404368
rect 66180 376718 66208 404359
rect 66168 376712 66220 376718
rect 66168 376654 66220 376660
rect 67100 375426 67128 471038
rect 67456 467832 67508 467838
rect 67456 467774 67508 467780
rect 67468 466857 67496 467774
rect 67454 466848 67510 466857
rect 67454 466783 67510 466792
rect 67362 453384 67418 453393
rect 67362 453319 67418 453328
rect 67376 451926 67404 453319
rect 67364 451920 67416 451926
rect 67364 451862 67416 451868
rect 67468 403034 67496 466783
rect 67456 403028 67508 403034
rect 67456 402970 67508 402976
rect 67364 392080 67416 392086
rect 67364 392022 67416 392028
rect 67376 391882 67404 392022
rect 67364 391876 67416 391882
rect 67364 391818 67416 391824
rect 67088 375420 67140 375426
rect 67088 375362 67140 375368
rect 67468 371793 67496 402970
rect 67560 380361 67588 474966
rect 67730 474943 67786 474952
rect 67640 473340 67692 473346
rect 67640 473282 67692 473288
rect 67652 472705 67680 473282
rect 67638 472696 67694 472705
rect 67638 472631 67694 472640
rect 67732 471096 67784 471102
rect 67730 471064 67732 471073
rect 67784 471064 67786 471073
rect 67730 470999 67786 471008
rect 67732 470484 67784 470490
rect 67732 470426 67784 470432
rect 67638 470248 67694 470257
rect 67638 470183 67640 470192
rect 67692 470183 67694 470192
rect 67640 470154 67692 470160
rect 67744 469713 67772 470426
rect 67730 469704 67786 469713
rect 67730 469639 67786 469648
rect 67638 468888 67694 468897
rect 67638 468823 67694 468832
rect 67652 468518 67680 468823
rect 67640 468512 67692 468518
rect 67640 468454 67692 468460
rect 67638 468208 67694 468217
rect 67638 468143 67694 468152
rect 67652 467974 67680 468143
rect 67640 467968 67692 467974
rect 67640 467910 67692 467916
rect 67640 466404 67692 466410
rect 67640 466346 67692 466352
rect 67652 465633 67680 466346
rect 67730 466168 67786 466177
rect 67730 466103 67786 466112
rect 67744 465730 67772 466103
rect 67732 465724 67784 465730
rect 67732 465666 67784 465672
rect 67638 465624 67694 465633
rect 67638 465559 67694 465568
rect 67638 464808 67694 464817
rect 67638 464743 67694 464752
rect 67652 464370 67680 464743
rect 67732 464432 67784 464438
rect 67732 464374 67784 464380
rect 67640 464364 67692 464370
rect 67640 464306 67692 464312
rect 67744 464273 67772 464374
rect 67730 464264 67786 464273
rect 67730 464199 67786 464208
rect 67638 462768 67694 462777
rect 67638 462703 67694 462712
rect 67652 462398 67680 462703
rect 67640 462392 67692 462398
rect 67640 462334 67692 462340
rect 67640 460216 67692 460222
rect 67638 460184 67640 460193
rect 67692 460184 67694 460193
rect 67638 460119 67694 460128
rect 67640 459536 67692 459542
rect 67640 459478 67692 459484
rect 67652 458833 67680 459478
rect 67730 459368 67786 459377
rect 67730 459303 67786 459312
rect 67638 458824 67694 458833
rect 67638 458759 67694 458768
rect 67744 458250 67772 459303
rect 67732 458244 67784 458250
rect 67732 458186 67784 458192
rect 67640 457496 67692 457502
rect 67638 457464 67640 457473
rect 67692 457464 67694 457473
rect 67638 457399 67694 457408
rect 67638 457328 67694 457337
rect 67638 457263 67694 457272
rect 67652 456822 67680 457263
rect 67640 456816 67692 456822
rect 67640 456758 67692 456764
rect 67732 456748 67784 456754
rect 67732 456690 67784 456696
rect 67744 456249 67772 456690
rect 67730 456240 67786 456249
rect 67730 456175 67786 456184
rect 67638 454608 67694 454617
rect 67638 454543 67694 454552
rect 67652 454102 67680 454543
rect 67640 454096 67692 454102
rect 67640 454038 67692 454044
rect 68006 454064 68062 454073
rect 68006 453999 68008 454008
rect 68060 453999 68062 454008
rect 68008 453970 68060 453976
rect 67640 453348 67692 453354
rect 67640 453290 67692 453296
rect 67652 453257 67680 453290
rect 67638 453248 67694 453257
rect 67638 453183 67694 453192
rect 67640 452600 67692 452606
rect 67638 452568 67640 452577
rect 67692 452568 67694 452577
rect 67638 452503 67694 452512
rect 67640 451240 67692 451246
rect 67640 451182 67692 451188
rect 67652 450809 67680 451182
rect 67638 450800 67694 450809
rect 67638 450735 67694 450744
rect 67730 449168 67786 449177
rect 67730 449103 67786 449112
rect 67744 448594 67772 449103
rect 67732 448588 67784 448594
rect 67732 448530 67784 448536
rect 67640 448520 67692 448526
rect 67638 448488 67640 448497
rect 67692 448488 67694 448497
rect 67638 448423 67694 448432
rect 67638 447264 67694 447273
rect 67638 447199 67694 447208
rect 67652 447166 67680 447199
rect 67640 447160 67692 447166
rect 67640 447102 67692 447108
rect 67638 446448 67694 446457
rect 67638 446383 67694 446392
rect 67652 445806 67680 446383
rect 67640 445800 67692 445806
rect 67640 445742 67692 445748
rect 67640 444372 67692 444378
rect 67640 444314 67692 444320
rect 67652 443873 67680 444314
rect 68204 444281 68232 543759
rect 68466 484664 68522 484673
rect 68466 484599 68522 484608
rect 68480 484430 68508 484599
rect 68468 484424 68520 484430
rect 68468 484366 68520 484372
rect 68664 477057 68692 576535
rect 68848 551449 68876 651335
rect 68926 644600 68982 644609
rect 68926 644535 68982 644544
rect 68834 551440 68890 551449
rect 68756 551398 68834 551426
rect 68650 477048 68706 477057
rect 68650 476983 68706 476992
rect 68190 444272 68246 444281
rect 68190 444207 68246 444216
rect 67638 443864 67694 443873
rect 67638 443799 67694 443808
rect 67730 442504 67786 442513
rect 67730 442439 67786 442448
rect 67638 442368 67694 442377
rect 67638 442303 67694 442312
rect 67652 442270 67680 442303
rect 67640 442264 67692 442270
rect 67640 442206 67692 442212
rect 67744 441658 67772 442439
rect 67732 441652 67784 441658
rect 67732 441594 67784 441600
rect 68204 441614 68232 444207
rect 68204 441586 68324 441614
rect 67640 441516 67692 441522
rect 67640 441458 67692 441464
rect 67652 441153 67680 441458
rect 67638 441144 67694 441153
rect 67638 441079 67694 441088
rect 67638 441008 67694 441017
rect 67638 440943 67694 440952
rect 67652 440910 67680 440943
rect 67640 440904 67692 440910
rect 67640 440846 67692 440852
rect 67640 385008 67692 385014
rect 67640 384950 67692 384956
rect 67652 384849 67680 384950
rect 67638 384840 67694 384849
rect 67638 384775 67694 384784
rect 67638 382528 67694 382537
rect 67638 382463 67694 382472
rect 67652 382294 67680 382463
rect 67640 382288 67692 382294
rect 67640 382230 67692 382236
rect 67638 380896 67694 380905
rect 67638 380831 67694 380840
rect 67546 380352 67602 380361
rect 67546 380287 67602 380296
rect 67652 379953 67680 380831
rect 67914 380760 67970 380769
rect 67914 380695 67970 380704
rect 67928 380186 67956 380695
rect 67916 380180 67968 380186
rect 67916 380122 67968 380128
rect 67638 379944 67694 379953
rect 67638 379879 67694 379888
rect 67638 377088 67694 377097
rect 67638 377023 67694 377032
rect 67652 376786 67680 377023
rect 67640 376780 67692 376786
rect 67640 376722 67692 376728
rect 67732 376712 67784 376718
rect 67732 376654 67784 376660
rect 67638 375592 67694 375601
rect 67638 375527 67694 375536
rect 67652 375426 67680 375527
rect 67640 375420 67692 375426
rect 67640 375362 67692 375368
rect 67640 374672 67692 374678
rect 67638 374640 67640 374649
rect 67692 374640 67694 374649
rect 67638 374575 67694 374584
rect 67744 374513 67772 376654
rect 67730 374504 67786 374513
rect 67730 374439 67786 374448
rect 67732 373992 67784 373998
rect 67732 373934 67784 373940
rect 67640 373312 67692 373318
rect 67744 373289 67772 373934
rect 67640 373254 67692 373260
rect 67730 373280 67786 373289
rect 67652 372473 67680 373254
rect 67730 373215 67786 373224
rect 67638 372464 67694 372473
rect 67638 372399 67694 372408
rect 67454 371784 67510 371793
rect 67454 371719 67510 371728
rect 67640 370524 67692 370530
rect 67640 370466 67692 370472
rect 67652 370433 67680 370466
rect 67638 370424 67694 370433
rect 67638 370359 67694 370368
rect 67640 369844 67692 369850
rect 67640 369786 67692 369792
rect 67652 369753 67680 369786
rect 67638 369744 67694 369753
rect 67638 369679 67694 369688
rect 67640 368552 67692 368558
rect 67638 368520 67640 368529
rect 67692 368520 67694 368529
rect 67638 368455 67694 368464
rect 67640 367056 67692 367062
rect 67638 367024 67640 367033
rect 67692 367024 67694 367033
rect 67638 366959 67694 366968
rect 67640 364336 67692 364342
rect 67638 364304 67640 364313
rect 68296 364334 68324 441586
rect 68664 398954 68692 476983
rect 68756 451897 68784 551398
rect 68834 551375 68890 551384
rect 68940 547874 68968 644535
rect 69124 581942 69152 680342
rect 69216 643249 69244 702578
rect 71044 692096 71096 692102
rect 71044 692038 71096 692044
rect 70032 681896 70084 681902
rect 70032 681838 70084 681844
rect 70044 679932 70072 681838
rect 70398 679824 70454 679833
rect 70454 679782 70702 679810
rect 70398 679759 70454 679768
rect 71056 679402 71084 692038
rect 71792 681018 71820 702714
rect 75184 700392 75236 700398
rect 75184 700334 75236 700340
rect 75196 685846 75224 700334
rect 75184 685840 75236 685846
rect 75184 685782 75236 685788
rect 77116 685840 77168 685846
rect 77116 685782 77168 685788
rect 75184 683188 75236 683194
rect 75184 683130 75236 683136
rect 74538 681864 74594 681873
rect 74538 681799 74594 681808
rect 71780 681012 71832 681018
rect 71780 680954 71832 680960
rect 72608 680400 72660 680406
rect 72608 680342 72660 680348
rect 72620 679932 72648 680342
rect 74552 679932 74580 681799
rect 75196 680513 75224 683130
rect 75182 680504 75238 680513
rect 75182 680439 75238 680448
rect 75196 679932 75224 680439
rect 77128 680377 77156 685782
rect 78600 683114 78628 702782
rect 78140 683086 78628 683114
rect 77114 680368 77170 680377
rect 77114 680303 77170 680312
rect 77128 679932 77156 680303
rect 78140 679425 78168 683086
rect 79336 680513 79364 702986
rect 80704 702500 80756 702506
rect 80704 702442 80756 702448
rect 80716 681834 80744 702442
rect 80704 681828 80756 681834
rect 80704 681770 80756 681776
rect 79322 680504 79378 680513
rect 79322 680439 79378 680448
rect 79336 679946 79364 680439
rect 80716 679946 80744 681770
rect 82096 680377 82124 703190
rect 89180 699825 89208 703520
rect 99288 703180 99340 703186
rect 99288 703122 99340 703128
rect 89166 699816 89222 699825
rect 89166 699751 89222 699760
rect 89720 686520 89772 686526
rect 89720 686462 89772 686468
rect 89074 680640 89130 680649
rect 89074 680575 89130 680584
rect 84842 680504 84898 680513
rect 84842 680439 84898 680448
rect 84856 680406 84884 680439
rect 84844 680400 84896 680406
rect 81622 680368 81678 680377
rect 81622 680303 81678 680312
rect 82082 680368 82138 680377
rect 84844 680342 84896 680348
rect 85486 680368 85542 680377
rect 82082 680303 82138 680312
rect 79336 679918 79718 679946
rect 80716 679918 81006 679946
rect 81636 679932 81664 680303
rect 84856 679932 84884 680342
rect 85486 680303 85542 680312
rect 85500 679932 85528 680303
rect 89088 679946 89116 680575
rect 89732 680513 89760 686462
rect 90640 681964 90692 681970
rect 90640 681906 90692 681912
rect 89718 680504 89774 680513
rect 89718 680439 89774 680448
rect 89732 679946 89760 680439
rect 89088 679918 89378 679946
rect 89732 679918 90022 679946
rect 90652 679932 90680 681906
rect 99300 681873 99328 703122
rect 102232 683800 102284 683806
rect 102232 683742 102284 683748
rect 98550 681864 98606 681873
rect 98550 681799 98606 681808
rect 99286 681864 99342 681873
rect 99286 681799 99342 681808
rect 91926 680368 91982 680377
rect 91926 680303 91982 680312
rect 91940 679932 91968 680303
rect 94870 679688 94926 679697
rect 96802 679688 96858 679697
rect 94926 679646 95174 679674
rect 94870 679623 94926 679632
rect 96858 679646 97106 679674
rect 96802 679623 96858 679632
rect 81898 679552 81954 679561
rect 85762 679552 85818 679561
rect 81954 679510 82294 679538
rect 81898 679487 81954 679496
rect 92938 679552 92994 679561
rect 85818 679510 86158 679538
rect 85762 679487 85818 679496
rect 96158 679552 96214 679561
rect 92994 679510 93242 679538
rect 92938 679487 92994 679496
rect 96214 679510 96462 679538
rect 96158 679487 96214 679496
rect 98564 679425 98592 681799
rect 102244 679946 102272 683742
rect 104912 681018 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 115204 703112 115256 703118
rect 115204 703054 115256 703060
rect 107568 702976 107620 702982
rect 107568 702918 107620 702924
rect 107580 681873 107608 702918
rect 113824 702772 113876 702778
rect 113824 702714 113876 702720
rect 113088 702568 113140 702574
rect 113088 702510 113140 702516
rect 110604 697604 110656 697610
rect 110604 697546 110656 697552
rect 106922 681864 106978 681873
rect 106922 681799 106978 681808
rect 107566 681864 107622 681873
rect 107566 681799 107622 681808
rect 104900 681012 104952 681018
rect 104900 680954 104952 680960
rect 102506 680504 102562 680513
rect 102506 680439 102562 680448
rect 102520 679946 102548 680439
rect 104806 680368 104862 680377
rect 104806 680303 104862 680312
rect 102244 679932 102364 679946
rect 102258 679918 102364 679932
rect 102520 679918 102902 679946
rect 104820 679932 104848 680303
rect 100666 679688 100722 679697
rect 100722 679646 100970 679674
rect 100666 679623 100722 679632
rect 99378 679552 99434 679561
rect 99434 679510 99682 679538
rect 99378 679487 99434 679496
rect 71778 679416 71834 679425
rect 71056 679386 71346 679402
rect 69296 679380 69348 679386
rect 69296 679322 69348 679328
rect 71044 679380 71346 679386
rect 71096 679374 71346 679380
rect 73618 679416 73674 679425
rect 71834 679374 71990 679402
rect 71778 679351 71834 679360
rect 75458 679416 75514 679425
rect 73674 679374 73922 679402
rect 73618 679351 73674 679360
rect 76194 679416 76250 679425
rect 75514 679374 75854 679402
rect 75458 679351 75514 679360
rect 78126 679416 78182 679425
rect 76250 679374 76498 679402
rect 77786 679374 78126 679402
rect 76194 679351 76250 679360
rect 78126 679351 78182 679360
rect 78862 679416 78918 679425
rect 80150 679416 80206 679425
rect 78918 679374 79074 679402
rect 78862 679351 78918 679360
rect 82726 679416 82782 679425
rect 80206 679374 80362 679402
rect 80150 679351 80206 679360
rect 84474 679416 84530 679425
rect 82782 679374 82938 679402
rect 84226 679374 84474 679402
rect 82726 679351 82782 679360
rect 84474 679351 84530 679360
rect 86498 679416 86554 679425
rect 87142 679416 87198 679425
rect 86554 679374 86802 679402
rect 86498 679351 86554 679360
rect 87786 679416 87842 679425
rect 87198 679374 87446 679402
rect 87142 679351 87198 679360
rect 91466 679416 91522 679425
rect 87842 679374 88090 679402
rect 91310 679374 91466 679402
rect 87786 679351 87842 679360
rect 92754 679416 92810 679425
rect 92598 679374 92754 679402
rect 91466 679351 91522 679360
rect 92754 679351 92810 679360
rect 94226 679416 94282 679425
rect 96158 679416 96214 679425
rect 94282 679374 94530 679402
rect 95818 679374 96158 679402
rect 94226 679351 94282 679360
rect 96158 679351 96214 679360
rect 97354 679416 97410 679425
rect 98550 679416 98606 679425
rect 97410 679374 97750 679402
rect 98394 679374 98550 679402
rect 97354 679351 97410 679360
rect 98550 679351 98606 679360
rect 100022 679416 100078 679425
rect 101310 679416 101366 679425
rect 100078 679374 100326 679402
rect 100022 679351 100078 679360
rect 102336 679402 102364 679918
rect 103334 679824 103390 679833
rect 103334 679759 103390 679768
rect 103348 679674 103376 679759
rect 103348 679646 103546 679674
rect 106936 679561 106964 681799
rect 109316 681760 109368 681766
rect 109316 681702 109368 681708
rect 107658 680504 107714 680513
rect 107658 680439 107714 680448
rect 107672 679946 107700 680439
rect 107672 679918 108054 679946
rect 109328 679932 109356 681702
rect 108394 679688 108450 679697
rect 108450 679646 108698 679674
rect 108394 679623 108450 679632
rect 105818 679552 105874 679561
rect 106922 679552 106978 679561
rect 105874 679510 106122 679538
rect 106766 679510 106922 679538
rect 105818 679487 105874 679496
rect 106922 679487 106978 679496
rect 102598 679416 102654 679425
rect 101366 679374 101614 679402
rect 102258 679374 102598 679402
rect 101310 679351 101366 679360
rect 105634 679416 105690 679425
rect 105478 679374 105634 679402
rect 102598 679351 102654 679360
rect 105634 679351 105690 679360
rect 107106 679416 107162 679425
rect 107162 679374 107410 679402
rect 107106 679351 107162 679360
rect 71044 679322 71096 679328
rect 69202 643240 69258 643249
rect 69202 643175 69258 643184
rect 69204 637220 69256 637226
rect 69204 637162 69256 637168
rect 69112 581936 69164 581942
rect 69112 581878 69164 581884
rect 68848 547846 68968 547874
rect 68848 544513 68876 547846
rect 68834 544504 68890 544513
rect 68834 544439 68890 544448
rect 68848 460934 68876 544439
rect 69124 482633 69152 581878
rect 69216 557534 69244 637162
rect 69308 580689 69336 679322
rect 110418 672616 110474 672625
rect 110418 672551 110474 672560
rect 109040 658436 109092 658442
rect 109040 658378 109092 658384
rect 69664 643748 69716 643754
rect 69664 643690 69716 643696
rect 69676 584390 69704 643690
rect 69768 640070 70058 640098
rect 69768 637226 69796 640070
rect 69756 637220 69808 637226
rect 69756 637162 69808 637168
rect 70688 630018 70716 640098
rect 71332 638994 71360 640098
rect 71320 638988 71372 638994
rect 71320 638930 71372 638936
rect 71976 635798 72004 640098
rect 71964 635792 72016 635798
rect 71964 635734 72016 635740
rect 72620 635610 72648 640098
rect 72700 638512 72752 638518
rect 72700 638454 72752 638460
rect 71792 635582 72648 635610
rect 71792 632738 71820 635582
rect 71780 632732 71832 632738
rect 71780 632674 71832 632680
rect 70676 630012 70728 630018
rect 70676 629954 70728 629960
rect 72712 625154 72740 638454
rect 73264 635730 73292 640098
rect 73908 638926 73936 640098
rect 73896 638920 73948 638926
rect 73896 638862 73948 638868
rect 74552 637650 74580 640098
rect 75823 640070 75868 640098
rect 74448 637628 74500 637634
rect 74552 637622 74672 637650
rect 74448 637574 74500 637576
rect 74448 637570 74580 637574
rect 74460 637546 74580 637570
rect 74552 636954 74580 637546
rect 74540 636948 74592 636954
rect 74540 636890 74592 636896
rect 73252 635724 73304 635730
rect 73252 635666 73304 635672
rect 73804 635724 73856 635730
rect 73804 635666 73856 635672
rect 72436 625126 72740 625154
rect 70766 586392 70822 586401
rect 70766 586327 70822 586336
rect 70398 585168 70454 585177
rect 70398 585103 70454 585112
rect 69664 584384 69716 584390
rect 69664 584326 69716 584332
rect 70308 584384 70360 584390
rect 70308 584326 70360 584332
rect 70320 583914 70348 584326
rect 70308 583908 70360 583914
rect 70308 583850 70360 583856
rect 69756 581936 69808 581942
rect 69808 581884 70058 581890
rect 69756 581878 70058 581884
rect 69768 581862 70058 581878
rect 70216 581732 70268 581738
rect 70216 581674 70268 581680
rect 70228 581233 70256 581674
rect 70214 581224 70270 581233
rect 70214 581159 70270 581168
rect 69294 580680 69350 580689
rect 69294 580615 69350 580624
rect 69662 580680 69718 580689
rect 69662 580615 69718 580624
rect 69676 579698 69704 580615
rect 69664 579692 69716 579698
rect 69664 579634 69716 579640
rect 69216 557506 69704 557534
rect 69676 540682 69704 557506
rect 69846 544368 69902 544377
rect 69846 544303 69902 544312
rect 69860 544218 69888 544303
rect 69860 544190 70164 544218
rect 69676 540654 70058 540682
rect 69676 528554 69704 540654
rect 70136 538218 70164 544190
rect 70320 540954 70348 583850
rect 70412 581233 70440 585103
rect 70492 581868 70544 581874
rect 70492 581810 70544 581816
rect 70398 581224 70454 581233
rect 70398 581159 70454 581168
rect 70412 581126 70440 581159
rect 70400 581120 70452 581126
rect 70400 581062 70452 581068
rect 70504 581058 70532 581810
rect 70780 581754 70808 586327
rect 71962 585576 72018 585585
rect 71962 585511 72018 585520
rect 71976 585206 72004 585511
rect 71964 585200 72016 585206
rect 71964 585142 72016 585148
rect 70950 584080 71006 584089
rect 70950 584015 71006 584024
rect 72238 584080 72294 584089
rect 72238 584015 72294 584024
rect 70964 581890 70992 584015
rect 72252 581890 72280 584015
rect 70964 581862 71300 581890
rect 71792 581874 72280 581890
rect 71780 581868 72280 581874
rect 71832 581862 72280 581868
rect 71780 581810 71832 581816
rect 72436 581806 72464 625126
rect 73342 586800 73398 586809
rect 73342 586735 73398 586744
rect 73356 586401 73384 586735
rect 73342 586392 73398 586401
rect 73342 586327 73398 586336
rect 72698 585576 72754 585585
rect 72698 585511 72754 585520
rect 72712 581890 72740 585511
rect 73356 581890 73384 586327
rect 72634 581862 72740 581890
rect 73278 581862 73384 581890
rect 70702 581726 70808 581754
rect 72424 581800 72476 581806
rect 72424 581742 72476 581748
rect 73816 581738 73844 635666
rect 74644 627230 74672 637622
rect 75840 637566 75868 640070
rect 75828 637560 75880 637566
rect 75828 637502 75880 637508
rect 75920 637492 75972 637498
rect 75920 637434 75972 637440
rect 75932 627366 75960 637434
rect 76484 629950 76512 640098
rect 77128 637498 77156 640098
rect 77390 638888 77446 638897
rect 77390 638823 77446 638832
rect 77116 637492 77168 637498
rect 77116 637434 77168 637440
rect 76472 629944 76524 629950
rect 76472 629886 76524 629892
rect 75920 627360 75972 627366
rect 75920 627302 75972 627308
rect 74632 627224 74684 627230
rect 74632 627166 74684 627172
rect 75734 589248 75790 589257
rect 75734 589183 75790 589192
rect 75644 585200 75696 585206
rect 75644 585142 75696 585148
rect 74630 583944 74686 583953
rect 74630 583879 74686 583888
rect 74644 581890 74672 583879
rect 75656 583817 75684 585142
rect 75274 583808 75330 583817
rect 75274 583743 75330 583752
rect 75642 583808 75698 583817
rect 75642 583743 75698 583752
rect 75288 581890 75316 583743
rect 75748 582486 75776 589183
rect 76746 587888 76802 587897
rect 76746 587823 76802 587832
rect 76010 585440 76066 585449
rect 76010 585375 76066 585384
rect 76024 585274 76052 585375
rect 76012 585268 76064 585274
rect 76012 585210 76064 585216
rect 75736 582480 75788 582486
rect 75736 582422 75788 582428
rect 75748 582162 75776 582422
rect 74566 581862 74672 581890
rect 75210 581862 75316 581890
rect 75656 582134 75776 582162
rect 75656 581754 75684 582134
rect 76024 581890 76052 585210
rect 76760 583778 76788 587823
rect 77404 585206 77432 638823
rect 77772 625154 77800 640098
rect 78416 637022 78444 640098
rect 79060 638314 79088 640098
rect 79048 638308 79100 638314
rect 79048 638250 79100 638256
rect 78404 637016 78456 637022
rect 78404 636958 78456 636964
rect 79704 627298 79732 640098
rect 80975 640070 81020 640098
rect 80992 639849 81020 640070
rect 80978 639840 81034 639849
rect 80978 639775 81034 639784
rect 80704 635656 80756 635662
rect 80704 635598 80756 635604
rect 79692 627292 79744 627298
rect 79692 627234 79744 627240
rect 77496 625126 77800 625154
rect 77496 624481 77524 625126
rect 77482 624472 77538 624481
rect 77482 624407 77538 624416
rect 79966 589248 80022 589257
rect 79966 589183 80022 589192
rect 78678 587752 78734 587761
rect 78678 587687 78734 587696
rect 78692 586673 78720 587687
rect 78678 586664 78734 586673
rect 78678 586599 78734 586608
rect 77392 585200 77444 585206
rect 77392 585142 77444 585148
rect 78218 585168 78274 585177
rect 78218 585103 78274 585112
rect 77392 583908 77444 583914
rect 77392 583850 77444 583856
rect 76748 583772 76800 583778
rect 76748 583714 76800 583720
rect 76760 581890 76788 583714
rect 77404 581890 77432 583850
rect 76024 581862 76452 581890
rect 76760 581862 77096 581890
rect 77404 581862 77740 581890
rect 78232 581754 78260 585103
rect 78692 581890 78720 586599
rect 79980 582418 80008 589183
rect 80716 583030 80744 635598
rect 80992 635594 81020 639775
rect 81438 638888 81494 638897
rect 81438 638823 81494 638832
rect 80980 635588 81032 635594
rect 80980 635530 81032 635536
rect 80796 591932 80848 591938
rect 80796 591874 80848 591880
rect 80808 585818 80836 591874
rect 80796 585812 80848 585818
rect 80796 585754 80848 585760
rect 80704 583024 80756 583030
rect 80704 582966 80756 582972
rect 79968 582412 80020 582418
rect 79968 582354 80020 582360
rect 79980 581890 80008 582354
rect 78692 581862 79028 581890
rect 79718 581862 80008 581890
rect 80808 581890 80836 585754
rect 81452 584458 81480 638823
rect 81636 632806 81664 640098
rect 82280 638450 82308 640098
rect 82268 638444 82320 638450
rect 82268 638386 82320 638392
rect 82924 638382 82952 640098
rect 82912 638376 82964 638382
rect 82912 638318 82964 638324
rect 83568 632942 83596 640098
rect 84212 638518 84240 640098
rect 84290 638888 84346 638897
rect 84290 638823 84346 638832
rect 84200 638512 84252 638518
rect 84200 638454 84252 638460
rect 83556 632936 83608 632942
rect 83556 632878 83608 632884
rect 81624 632800 81676 632806
rect 81624 632742 81676 632748
rect 84304 591938 84332 638823
rect 84856 636886 84884 640098
rect 86127 640070 86172 640098
rect 85580 637492 85632 637498
rect 85580 637434 85632 637440
rect 84844 636880 84896 636886
rect 84844 636822 84896 636828
rect 85592 629921 85620 637434
rect 86144 632874 86172 640070
rect 86788 637498 86816 640098
rect 86776 637492 86828 637498
rect 86776 637434 86828 637440
rect 86960 637492 87012 637498
rect 86960 637434 87012 637440
rect 86132 632868 86184 632874
rect 86132 632810 86184 632816
rect 86972 629921 87000 637434
rect 87432 634166 87460 640098
rect 88076 637498 88104 640098
rect 88064 637492 88116 637498
rect 88064 637434 88116 637440
rect 88720 636954 88748 640098
rect 88708 636948 88760 636954
rect 88708 636890 88760 636896
rect 87420 634160 87472 634166
rect 87420 634102 87472 634108
rect 85578 629912 85634 629921
rect 85578 629847 85634 629856
rect 86958 629912 87014 629921
rect 86958 629847 87014 629856
rect 89364 627201 89392 640098
rect 90008 632874 90036 640098
rect 91279 640070 91324 640098
rect 91296 635594 91324 640070
rect 91940 638246 91968 640098
rect 92386 638888 92442 638897
rect 92386 638823 92442 638832
rect 91928 638240 91980 638246
rect 91928 638182 91980 638188
rect 91284 635588 91336 635594
rect 91284 635530 91336 635536
rect 89996 632868 90048 632874
rect 89996 632810 90048 632816
rect 89350 627192 89406 627201
rect 89350 627127 89406 627136
rect 89626 593464 89682 593473
rect 89626 593399 89682 593408
rect 84292 591932 84344 591938
rect 84292 591874 84344 591880
rect 88246 588568 88302 588577
rect 88246 588503 88302 588512
rect 84290 588296 84346 588305
rect 84290 588231 84346 588240
rect 84106 586528 84162 586537
rect 84106 586463 84162 586472
rect 81440 584452 81492 584458
rect 81440 584394 81492 584400
rect 81452 581890 81480 584394
rect 84120 583846 84148 586463
rect 83372 583840 83424 583846
rect 84108 583840 84160 583846
rect 83372 583782 83424 583788
rect 84014 583808 84070 583817
rect 83278 582448 83334 582457
rect 83278 582383 83334 582392
rect 81898 582040 81954 582049
rect 81898 581975 81954 581984
rect 81912 581890 81940 581975
rect 83292 581890 83320 582383
rect 80808 581862 80960 581890
rect 81452 581862 81604 581890
rect 81912 581862 82248 581890
rect 82938 581862 83320 581890
rect 83384 581890 83412 583782
rect 84108 583782 84160 583788
rect 84014 583743 84070 583752
rect 84028 582457 84056 583743
rect 84014 582448 84070 582457
rect 84014 582383 84070 582392
rect 84304 581890 84332 588231
rect 85394 585440 85450 585449
rect 85394 585375 85450 585384
rect 85408 585274 85436 585375
rect 85396 585268 85448 585274
rect 85396 585210 85448 585216
rect 85118 585168 85174 585177
rect 85118 585103 85174 585112
rect 85132 582622 85160 585103
rect 85120 582616 85172 582622
rect 85120 582558 85172 582564
rect 85132 581890 85160 582558
rect 85408 582162 85436 585210
rect 86222 583808 86278 583817
rect 86222 583743 86278 583752
rect 86236 582554 86264 583743
rect 87696 583024 87748 583030
rect 87696 582966 87748 582972
rect 86224 582548 86276 582554
rect 86224 582490 86276 582496
rect 83384 581862 83536 581890
rect 84226 581862 84332 581890
rect 84870 581862 85160 581890
rect 85316 582134 85436 582162
rect 85316 581754 85344 582134
rect 86236 581890 86264 582490
rect 87708 582486 87736 582966
rect 87696 582480 87748 582486
rect 87696 582422 87748 582428
rect 87708 581890 87736 582422
rect 88260 581890 88288 588503
rect 88890 585168 88946 585177
rect 88890 585103 88946 585112
rect 88904 581890 88932 585103
rect 89640 584050 89668 593399
rect 91006 593328 91062 593337
rect 91006 593263 91062 593272
rect 90270 585168 90326 585177
rect 90270 585103 90326 585112
rect 89628 584044 89680 584050
rect 89628 583986 89680 583992
rect 89640 581890 89668 583986
rect 90284 581890 90312 585103
rect 91020 582554 91048 593263
rect 92400 589393 92428 638823
rect 92584 635730 92612 640098
rect 92572 635724 92624 635730
rect 92572 635666 92624 635672
rect 93228 635662 93256 640098
rect 93872 637634 93900 640098
rect 93860 637628 93912 637634
rect 93860 637570 93912 637576
rect 94516 635730 94544 640098
rect 95160 638761 95188 640098
rect 96431 640070 96476 640098
rect 95882 639704 95938 639713
rect 95882 639639 95938 639648
rect 95146 638752 95202 638761
rect 95146 638687 95202 638696
rect 95160 638518 95188 638687
rect 95148 638512 95200 638518
rect 95148 638454 95200 638460
rect 94504 635724 94556 635730
rect 94504 635666 94556 635672
rect 93216 635656 93268 635662
rect 93216 635598 93268 635604
rect 95896 596174 95924 639639
rect 96448 638246 96476 640070
rect 96436 638240 96488 638246
rect 96436 638182 96488 638188
rect 96528 638036 96580 638042
rect 96528 637978 96580 637984
rect 96540 635526 96568 637978
rect 96620 637492 96672 637498
rect 96620 637434 96672 637440
rect 96528 635520 96580 635526
rect 96528 635462 96580 635468
rect 96632 632738 96660 637434
rect 97092 632806 97120 640098
rect 97736 637498 97764 640098
rect 97724 637492 97776 637498
rect 97724 637434 97776 637440
rect 97080 632800 97132 632806
rect 97080 632742 97132 632748
rect 96620 632732 96672 632738
rect 96620 632674 96672 632680
rect 98380 629950 98408 640098
rect 99024 638450 99052 640098
rect 99012 638444 99064 638450
rect 99012 638386 99064 638392
rect 99668 638382 99696 640098
rect 100312 639010 100340 640098
rect 101583 640070 101628 640098
rect 99944 638982 100340 639010
rect 99656 638376 99708 638382
rect 99656 638318 99708 638324
rect 99668 638042 99696 638318
rect 99656 638036 99708 638042
rect 99656 637978 99708 637984
rect 99944 634166 99972 638982
rect 100298 638888 100354 638897
rect 100298 638823 100354 638832
rect 99932 634160 99984 634166
rect 99932 634102 99984 634108
rect 98368 629944 98420 629950
rect 98368 629886 98420 629892
rect 95896 596146 96108 596174
rect 91098 589384 91154 589393
rect 91098 589319 91154 589328
rect 92386 589384 92442 589393
rect 92386 589319 92442 589328
rect 91008 582548 91060 582554
rect 91008 582490 91060 582496
rect 91020 581890 91048 582490
rect 86158 581862 86264 581890
rect 87446 581862 87736 581890
rect 88090 581862 88288 581890
rect 88734 581862 88932 581890
rect 89378 581862 89668 581890
rect 90022 581862 90312 581890
rect 90666 581862 91048 581890
rect 91112 581890 91140 589319
rect 96080 588606 96108 596146
rect 96434 590064 96490 590073
rect 96434 589999 96490 590008
rect 96448 589966 96476 589999
rect 96160 589960 96212 589966
rect 96160 589902 96212 589908
rect 96436 589960 96488 589966
rect 96436 589902 96488 589908
rect 97262 589928 97318 589937
rect 96068 588600 96120 588606
rect 96068 588542 96120 588548
rect 96080 587926 96108 588542
rect 92296 587920 92348 587926
rect 92296 587862 92348 587868
rect 96068 587920 96120 587926
rect 96068 587862 96120 587868
rect 92308 581890 92336 587862
rect 94962 587208 95018 587217
rect 94962 587143 95018 587152
rect 94872 584248 94924 584254
rect 94872 584190 94924 584196
rect 93766 583808 93822 583817
rect 93766 583743 93822 583752
rect 93780 582418 93808 583743
rect 94134 582584 94190 582593
rect 94134 582519 94190 582528
rect 92848 582412 92900 582418
rect 92848 582354 92900 582360
rect 93768 582412 93820 582418
rect 93768 582354 93820 582360
rect 92860 581890 92888 582354
rect 94148 581890 94176 582519
rect 94884 581890 94912 584190
rect 91112 581862 91264 581890
rect 91954 581862 92336 581890
rect 92598 581862 92888 581890
rect 93886 581862 94176 581890
rect 94530 581862 94912 581890
rect 94976 581754 95004 587143
rect 96172 583846 96200 589902
rect 97262 589863 97318 589872
rect 96526 589248 96582 589257
rect 96526 589183 96582 589192
rect 96540 583914 96568 589183
rect 97170 587888 97226 587897
rect 97170 587823 97226 587832
rect 97184 586634 97212 587823
rect 97172 586628 97224 586634
rect 97172 586570 97224 586576
rect 97078 585168 97134 585177
rect 97078 585103 97134 585112
rect 97092 584066 97120 585103
rect 97184 584254 97212 586570
rect 97172 584248 97224 584254
rect 97172 584190 97224 584196
rect 97092 584038 97212 584066
rect 96528 583908 96580 583914
rect 96528 583850 96580 583856
rect 96160 583840 96212 583846
rect 96160 583782 96212 583788
rect 96172 581890 96200 583782
rect 96540 581890 96568 583850
rect 97184 581890 97212 584038
rect 95818 581862 96200 581890
rect 96462 581862 96568 581890
rect 97106 581862 97212 581890
rect 97276 581890 97304 589863
rect 100312 586514 100340 638823
rect 101404 637628 101456 637634
rect 101404 637570 101456 637576
rect 100128 586486 100340 586514
rect 98734 586392 98790 586401
rect 98734 586327 98790 586336
rect 98748 581890 98776 586327
rect 99102 584080 99158 584089
rect 99102 584015 99158 584024
rect 99116 583817 99144 584015
rect 99102 583808 99158 583817
rect 99102 583743 99158 583752
rect 99116 581890 99144 583743
rect 97276 581862 97704 581890
rect 98394 581862 98776 581890
rect 99038 581862 99144 581890
rect 100128 581754 100156 586486
rect 101310 585576 101366 585585
rect 101310 585511 101366 585520
rect 100574 581904 100630 581913
rect 101324 581890 101352 585511
rect 100970 581862 101352 581890
rect 100574 581839 100630 581848
rect 100588 581754 100616 581839
rect 101416 581806 101444 637570
rect 101600 637022 101628 640070
rect 101588 637016 101640 637022
rect 101588 636958 101640 636964
rect 102244 635526 102272 640098
rect 102888 638314 102916 640098
rect 103426 638888 103482 638897
rect 103426 638823 103482 638832
rect 102876 638308 102928 638314
rect 102876 638250 102928 638256
rect 102232 635520 102284 635526
rect 102232 635462 102284 635468
rect 103150 587480 103206 587489
rect 103150 587415 103206 587424
rect 101864 585132 101916 585138
rect 101864 585074 101916 585080
rect 101876 581890 101904 585074
rect 102600 583772 102652 583778
rect 102600 583714 102652 583720
rect 102612 581890 102640 583714
rect 103164 581890 103192 587415
rect 103440 583778 103468 638823
rect 103532 636886 103560 640098
rect 104176 638926 104204 640098
rect 104164 638920 104216 638926
rect 104164 638862 104216 638868
rect 104820 637498 104848 640098
rect 105464 637673 105492 640098
rect 106735 640070 106780 640098
rect 105544 638512 105596 638518
rect 105544 638454 105596 638460
rect 105450 637664 105506 637673
rect 105450 637599 105506 637608
rect 103612 637492 103664 637498
rect 103612 637434 103664 637440
rect 104808 637492 104860 637498
rect 104808 637434 104860 637440
rect 103520 636880 103572 636886
rect 103520 636822 103572 636828
rect 103624 596174 103652 637434
rect 105556 596174 105584 638454
rect 106752 625154 106780 640070
rect 107396 638625 107424 640098
rect 107382 638616 107438 638625
rect 107382 638551 107438 638560
rect 108040 634098 108068 640098
rect 108698 640070 108988 640098
rect 108856 639668 108908 639674
rect 108856 639610 108908 639616
rect 108868 634814 108896 639610
rect 108960 638518 108988 640070
rect 108948 638512 109000 638518
rect 108948 638454 109000 638460
rect 108868 634786 108988 634814
rect 108028 634092 108080 634098
rect 108028 634034 108080 634040
rect 107568 633004 107620 633010
rect 107568 632946 107620 632952
rect 106292 625126 106780 625154
rect 103624 596146 103744 596174
rect 105556 596146 105860 596174
rect 103428 583772 103480 583778
rect 103428 583714 103480 583720
rect 103716 582010 103744 596146
rect 105542 585576 105598 585585
rect 105542 585511 105598 585520
rect 105556 585138 105584 585511
rect 105544 585132 105596 585138
rect 105544 585074 105596 585080
rect 103888 584520 103940 584526
rect 103888 584462 103940 584468
rect 103704 582004 103756 582010
rect 103704 581946 103756 581952
rect 103900 581890 103928 584462
rect 104622 584080 104678 584089
rect 104622 584015 104678 584024
rect 104438 583944 104494 583953
rect 104438 583879 104494 583888
rect 101614 581862 101904 581890
rect 102258 581862 102640 581890
rect 102902 581862 103192 581890
rect 103546 581862 103928 581890
rect 73804 581732 73856 581738
rect 75656 581726 75808 581754
rect 78232 581726 78384 581754
rect 85316 581726 85468 581754
rect 94976 581726 95128 581754
rect 100128 581726 100616 581754
rect 101404 581800 101456 581806
rect 104452 581754 104480 583879
rect 101404 581742 101456 581748
rect 104190 581738 104480 581754
rect 104636 581754 104664 584015
rect 105728 583976 105780 583982
rect 105728 583918 105780 583924
rect 105740 581890 105768 583918
rect 105478 581862 105768 581890
rect 104190 581732 104492 581738
rect 104190 581726 104440 581732
rect 73804 581674 73856 581680
rect 104636 581726 104788 581754
rect 105636 581732 105688 581738
rect 104440 581674 104492 581680
rect 105636 581674 105688 581680
rect 105648 581058 105676 581674
rect 70492 581052 70544 581058
rect 70492 580994 70544 581000
rect 105636 581052 105688 581058
rect 105636 580994 105688 581000
rect 105832 580310 105860 596146
rect 105820 580304 105872 580310
rect 105820 580246 105872 580252
rect 106094 578232 106150 578241
rect 106094 578167 106150 578176
rect 105636 574524 105688 574530
rect 105636 574466 105688 574472
rect 105648 574433 105676 574466
rect 105634 574424 105690 574433
rect 105634 574359 105690 574368
rect 105648 567194 105676 574359
rect 106108 567194 106136 578167
rect 105556 567166 105676 567194
rect 105740 567166 106136 567194
rect 105556 557534 105584 567166
rect 105556 557506 105676 557534
rect 105648 555150 105676 557506
rect 105636 555144 105688 555150
rect 105636 555086 105688 555092
rect 70320 540926 70440 540954
rect 70124 538212 70176 538218
rect 70412 538214 70440 540926
rect 105478 540382 105676 540410
rect 70504 540110 70702 540138
rect 70504 539782 70532 540110
rect 70492 539776 70544 539782
rect 70492 539718 70544 539724
rect 71332 539646 71360 540138
rect 71976 539714 72004 540138
rect 71964 539708 72016 539714
rect 71964 539650 72016 539656
rect 71320 539640 71372 539646
rect 71320 539582 71372 539588
rect 70412 538186 70532 538214
rect 70124 538154 70176 538160
rect 69308 528526 69704 528554
rect 68926 482624 68982 482633
rect 68926 482559 68982 482568
rect 69110 482624 69166 482633
rect 69110 482559 69166 482568
rect 68940 481710 68968 482559
rect 69018 482488 69074 482497
rect 69018 482423 69074 482432
rect 68928 481704 68980 481710
rect 68928 481646 68980 481652
rect 69032 480254 69060 482423
rect 69202 480584 69258 480593
rect 69202 480519 69258 480528
rect 69032 480226 69152 480254
rect 68926 473784 68982 473793
rect 68926 473719 68982 473728
rect 68940 473385 68968 473719
rect 68926 473376 68982 473385
rect 68926 473311 68982 473320
rect 68848 460906 68968 460934
rect 68742 451888 68798 451897
rect 68742 451823 68798 451832
rect 68756 451274 68784 451823
rect 68756 451246 68876 451274
rect 68848 446434 68876 451246
rect 68756 446406 68876 446434
rect 68652 398948 68704 398954
rect 68652 398890 68704 398896
rect 68664 386866 68692 398890
rect 68756 394670 68784 446406
rect 68940 445505 68968 460906
rect 68926 445496 68982 445505
rect 68848 445454 68926 445482
rect 68744 394664 68796 394670
rect 68744 394606 68796 394612
rect 68664 386838 68784 386866
rect 68756 383722 68784 386838
rect 68744 383716 68796 383722
rect 68744 383658 68796 383664
rect 68756 383489 68784 383658
rect 68742 383480 68798 383489
rect 68742 383415 68798 383424
rect 67692 364304 67694 364313
rect 68296 364306 68692 364334
rect 67638 364239 67694 364248
rect 67640 362908 67692 362914
rect 67640 362850 67692 362856
rect 67652 362681 67680 362850
rect 67638 362672 67694 362681
rect 67638 362607 67694 362616
rect 67638 360768 67694 360777
rect 67638 360703 67694 360712
rect 67652 360262 67680 360703
rect 67640 360256 67692 360262
rect 67640 360198 67692 360204
rect 67730 360224 67786 360233
rect 67730 360159 67786 360168
rect 67638 359680 67694 359689
rect 67638 359615 67694 359624
rect 67652 359582 67680 359615
rect 67640 359576 67692 359582
rect 67640 359518 67692 359524
rect 67744 359514 67772 360159
rect 67732 359508 67784 359514
rect 67732 359450 67784 359456
rect 67546 358184 67602 358193
rect 67546 358119 67602 358128
rect 67560 357406 67588 358119
rect 67640 358080 67692 358086
rect 67638 358048 67640 358057
rect 67692 358048 67694 358057
rect 67638 357983 67694 357992
rect 66904 357400 66956 357406
rect 66904 357342 66956 357348
rect 67548 357400 67600 357406
rect 67548 357342 67600 357348
rect 65616 349036 65668 349042
rect 65616 348978 65668 348984
rect 66168 347744 66220 347750
rect 66166 347712 66168 347721
rect 66220 347712 66222 347721
rect 66166 347647 66222 347656
rect 66168 340944 66220 340950
rect 66168 340886 66220 340892
rect 66180 330614 66208 340886
rect 66168 330608 66220 330614
rect 66168 330550 66220 330556
rect 66916 327894 66944 357342
rect 68006 356960 68062 356969
rect 68006 356895 68062 356904
rect 68020 356114 68048 356895
rect 68008 356108 68060 356114
rect 68008 356050 68060 356056
rect 67730 355600 67786 355609
rect 67730 355535 67786 355544
rect 67640 355428 67692 355434
rect 67640 355370 67692 355376
rect 67652 355201 67680 355370
rect 67744 355366 67772 355535
rect 67732 355360 67784 355366
rect 67732 355302 67784 355308
rect 67638 355192 67694 355201
rect 67638 355127 67694 355136
rect 67546 353832 67602 353841
rect 67546 353767 67602 353776
rect 67560 353258 67588 353767
rect 66996 353252 67048 353258
rect 66996 353194 67048 353200
rect 67548 353252 67600 353258
rect 67548 353194 67600 353200
rect 67008 338774 67036 353194
rect 67640 351892 67692 351898
rect 67640 351834 67692 351840
rect 67652 351801 67680 351834
rect 67638 351792 67694 351801
rect 67638 351727 67694 351736
rect 67638 349208 67694 349217
rect 67638 349143 67640 349152
rect 67692 349143 67694 349152
rect 67640 349114 67692 349120
rect 67638 349072 67694 349081
rect 67638 349007 67640 349016
rect 67692 349007 67694 349016
rect 67640 348978 67692 348984
rect 67640 347744 67692 347750
rect 67638 347712 67640 347721
rect 67692 347712 67694 347721
rect 67638 347647 67694 347656
rect 68664 345098 68692 364306
rect 68848 346390 68876 445454
rect 68926 445431 68982 445440
rect 69124 439278 69152 480226
rect 69112 439272 69164 439278
rect 69112 439214 69164 439220
rect 69216 439113 69244 480519
rect 69308 460934 69336 528526
rect 70504 499574 70532 538186
rect 72620 535430 72648 540138
rect 73264 537946 73292 540138
rect 73344 538960 73396 538966
rect 73344 538902 73396 538908
rect 73356 537946 73384 538902
rect 73252 537940 73304 537946
rect 73252 537882 73304 537888
rect 73344 537940 73396 537946
rect 73344 537882 73396 537888
rect 73356 536858 73384 537882
rect 73344 536852 73396 536858
rect 73344 536794 73396 536800
rect 73804 536852 73856 536858
rect 73804 536794 73856 536800
rect 72608 535424 72660 535430
rect 72608 535366 72660 535372
rect 70504 499546 70900 499574
rect 70872 492833 70900 499546
rect 73816 494766 73844 536794
rect 73908 536110 73936 540138
rect 74552 537878 74580 540138
rect 75196 539510 75224 540138
rect 76467 540110 76512 540138
rect 75184 539504 75236 539510
rect 75184 539446 75236 539452
rect 74540 537872 74592 537878
rect 74540 537814 74592 537820
rect 74538 537432 74594 537441
rect 74538 537367 74594 537376
rect 73896 536104 73948 536110
rect 73896 536046 73948 536052
rect 73804 494760 73856 494766
rect 73804 494702 73856 494708
rect 70858 492824 70914 492833
rect 70858 492759 70914 492768
rect 70400 492040 70452 492046
rect 70400 491982 70452 491988
rect 70032 491496 70084 491502
rect 70032 491438 70084 491444
rect 70044 489940 70072 491438
rect 70412 489954 70440 491982
rect 70872 489954 70900 492759
rect 71780 491972 71832 491978
rect 71780 491914 71832 491920
rect 71792 489954 71820 491914
rect 74552 491434 74580 537367
rect 76484 533390 76512 540110
rect 76472 533384 76524 533390
rect 76472 533326 76524 533332
rect 77128 530670 77156 540138
rect 77772 539442 77800 540138
rect 77760 539436 77812 539442
rect 77760 539378 77812 539384
rect 78416 538014 78444 540138
rect 78404 538008 78456 538014
rect 78404 537950 78456 537956
rect 79060 535294 79088 540138
rect 79048 535288 79100 535294
rect 79048 535230 79100 535236
rect 79704 535226 79732 540138
rect 80348 538150 80376 540138
rect 80336 538144 80388 538150
rect 80336 538086 80388 538092
rect 80992 537946 81020 540138
rect 81636 538121 81664 540138
rect 82907 540110 82952 540138
rect 81622 538112 81678 538121
rect 81622 538047 81678 538056
rect 80980 537940 81032 537946
rect 80980 537882 81032 537888
rect 82820 536852 82872 536858
rect 82820 536794 82872 536800
rect 82832 536654 82860 536794
rect 82924 536722 82952 540110
rect 83568 538082 83596 540138
rect 83556 538076 83608 538082
rect 83556 538018 83608 538024
rect 83464 536852 83516 536858
rect 83464 536794 83516 536800
rect 82912 536716 82964 536722
rect 82912 536658 82964 536664
rect 82820 536648 82872 536654
rect 82820 536590 82872 536596
rect 79692 535220 79744 535226
rect 79692 535162 79744 535168
rect 77116 530664 77168 530670
rect 77116 530606 77168 530612
rect 79324 530596 79376 530602
rect 79324 530538 79376 530544
rect 76470 494728 76526 494737
rect 76470 494663 76526 494672
rect 74998 492824 75054 492833
rect 74998 492759 75054 492768
rect 74540 491428 74592 491434
rect 74540 491370 74592 491376
rect 72240 490612 72292 490618
rect 72240 490554 72292 490560
rect 72252 489954 72280 490554
rect 74356 490000 74408 490006
rect 70412 489926 70656 489954
rect 70872 489926 71300 489954
rect 71792 489926 71944 489954
rect 72252 489926 72588 489954
rect 73080 489938 73232 489954
rect 75012 489954 75040 492759
rect 75460 491428 75512 491434
rect 75460 491370 75512 491376
rect 75472 489954 75500 491370
rect 74408 489948 74520 489954
rect 74356 489942 74520 489948
rect 73068 489932 73232 489938
rect 73120 489926 73232 489932
rect 74368 489926 74520 489942
rect 75012 489926 75164 489954
rect 75472 489926 75808 489954
rect 76484 489940 76512 494663
rect 79336 492726 79364 530538
rect 82912 497480 82964 497486
rect 82912 497422 82964 497428
rect 82820 495576 82872 495582
rect 82820 495518 82872 495524
rect 80980 493400 81032 493406
rect 80980 493342 81032 493348
rect 79690 492824 79746 492833
rect 79690 492759 79746 492768
rect 79324 492720 79376 492726
rect 79324 492662 79376 492668
rect 77760 492652 77812 492658
rect 77760 492594 77812 492600
rect 78404 492652 78456 492658
rect 78404 492594 78456 492600
rect 76748 491564 76800 491570
rect 76748 491506 76800 491512
rect 76760 489954 76788 491506
rect 76760 489926 77096 489954
rect 77772 489940 77800 492594
rect 78416 489940 78444 492594
rect 79704 489940 79732 492759
rect 80060 491360 80112 491366
rect 80060 491302 80112 491308
rect 80072 489954 80100 491302
rect 80072 489926 80316 489954
rect 80992 489940 81020 493342
rect 81900 492788 81952 492794
rect 81900 492730 81952 492736
rect 81624 492108 81676 492114
rect 81624 492050 81676 492056
rect 81636 489940 81664 492050
rect 81912 489954 81940 492730
rect 82832 492658 82860 495518
rect 82924 494018 82952 497422
rect 83476 496097 83504 536794
rect 84212 534002 84240 540138
rect 84856 534070 84884 540138
rect 85500 536858 85528 540138
rect 86144 538218 86172 540138
rect 86132 538214 86184 538218
rect 86132 538212 86264 538214
rect 86184 538186 86264 538212
rect 86132 538154 86184 538160
rect 85488 536852 85540 536858
rect 85488 536794 85540 536800
rect 84844 534064 84896 534070
rect 84844 534006 84896 534012
rect 84200 533996 84252 534002
rect 84200 533938 84252 533944
rect 83556 533452 83608 533458
rect 83556 533394 83608 533400
rect 83462 496088 83518 496097
rect 83462 496023 83518 496032
rect 83568 495582 83596 533394
rect 86236 498817 86264 538186
rect 86788 535362 86816 540138
rect 87432 537538 87460 540138
rect 87420 537532 87472 537538
rect 87420 537474 87472 537480
rect 88076 536722 88104 540138
rect 89347 540110 89392 540138
rect 89364 537606 89392 540110
rect 89352 537600 89404 537606
rect 89352 537542 89404 537548
rect 88064 536716 88116 536722
rect 88064 536658 88116 536664
rect 86776 535356 86828 535362
rect 86776 535298 86828 535304
rect 90008 534818 90036 540138
rect 89996 534812 90048 534818
rect 89996 534754 90048 534760
rect 89628 533520 89680 533526
rect 89628 533462 89680 533468
rect 86958 531992 87014 532001
rect 86958 531927 87014 531936
rect 86222 498808 86278 498817
rect 86222 498743 86278 498752
rect 86132 498228 86184 498234
rect 86132 498170 86184 498176
rect 84842 497448 84898 497457
rect 84842 497383 84898 497392
rect 83556 495576 83608 495582
rect 83556 495518 83608 495524
rect 82912 494012 82964 494018
rect 82912 493954 82964 493960
rect 83556 494012 83608 494018
rect 83556 493954 83608 493960
rect 82912 493332 82964 493338
rect 82912 493274 82964 493280
rect 82820 492652 82872 492658
rect 82820 492594 82872 492600
rect 81912 489926 82248 489954
rect 82924 489940 82952 493274
rect 83568 489940 83596 493954
rect 84856 489940 84884 497383
rect 85488 495440 85540 495446
rect 85488 495382 85540 495388
rect 85500 489940 85528 495382
rect 86144 489940 86172 498170
rect 86776 491360 86828 491366
rect 86776 491302 86828 491308
rect 86788 489940 86816 491302
rect 86972 489954 87000 531927
rect 89640 493882 89668 533462
rect 90652 533390 90680 540138
rect 91296 538214 91324 540138
rect 91020 538186 91324 538214
rect 91020 536790 91048 538186
rect 91008 536784 91060 536790
rect 91940 536761 91968 540138
rect 91008 536726 91060 536732
rect 91926 536752 91982 536761
rect 90640 533384 90692 533390
rect 90640 533326 90692 533332
rect 91020 530738 91048 536726
rect 91926 536687 91982 536696
rect 91940 530738 91968 536687
rect 92584 535430 92612 540138
rect 93228 537878 93256 540138
rect 93872 539186 93900 540138
rect 93872 539158 93992 539186
rect 93860 538892 93912 538898
rect 93860 538834 93912 538840
rect 93872 538218 93900 538834
rect 93860 538212 93912 538218
rect 93860 538154 93912 538160
rect 93216 537872 93268 537878
rect 93216 537814 93268 537820
rect 93768 537872 93820 537878
rect 93768 537814 93820 537820
rect 92572 535424 92624 535430
rect 92572 535366 92624 535372
rect 93674 532128 93730 532137
rect 93674 532063 93730 532072
rect 91008 530732 91060 530738
rect 91008 530674 91060 530680
rect 91928 530732 91980 530738
rect 91928 530674 91980 530680
rect 91008 530596 91060 530602
rect 91008 530538 91060 530544
rect 90640 494828 90692 494834
rect 90640 494770 90692 494776
rect 89996 494284 90048 494290
rect 89996 494226 90048 494232
rect 88708 493876 88760 493882
rect 88708 493818 88760 493824
rect 89628 493876 89680 493882
rect 89628 493818 89680 493824
rect 88720 492794 88748 493818
rect 88708 492788 88760 492794
rect 88708 492730 88760 492736
rect 88064 492040 88116 492046
rect 88064 491982 88116 491988
rect 87372 490104 87428 490113
rect 87372 490039 87428 490048
rect 87386 489954 87414 490039
rect 86972 489940 87414 489954
rect 88076 489940 88104 491982
rect 88720 489940 88748 492730
rect 90008 489940 90036 494226
rect 90652 489940 90680 494770
rect 91020 491366 91048 530538
rect 91100 498840 91152 498846
rect 91100 498782 91152 498788
rect 91112 492250 91140 498782
rect 93688 494086 93716 532063
rect 92480 494080 92532 494086
rect 92480 494022 92532 494028
rect 93676 494080 93728 494086
rect 93676 494022 93728 494028
rect 91100 492244 91152 492250
rect 91100 492186 91152 492192
rect 91008 491360 91060 491366
rect 91008 491302 91060 491308
rect 91112 489954 91140 492186
rect 92492 492114 92520 494022
rect 92480 492108 92532 492114
rect 92480 492050 92532 492056
rect 92572 491632 92624 491638
rect 92572 491574 92624 491580
rect 91928 491496 91980 491502
rect 91928 491438 91980 491444
rect 91744 491360 91796 491366
rect 91744 491302 91796 491308
rect 91756 490686 91784 491302
rect 91744 490680 91796 490686
rect 91744 490622 91796 490628
rect 86972 489926 87400 489940
rect 91112 489926 91264 489954
rect 91940 489940 91968 491438
rect 92584 489940 92612 491574
rect 93216 491564 93268 491570
rect 93216 491506 93268 491512
rect 93228 489940 93256 491506
rect 93780 490618 93808 537814
rect 93964 536654 93992 539158
rect 94042 538792 94098 538801
rect 94042 538727 94098 538736
rect 93952 536648 94004 536654
rect 93952 536590 94004 536596
rect 94056 528554 94084 538727
rect 94516 538082 94544 540138
rect 95787 540110 95832 540138
rect 94504 538076 94556 538082
rect 94504 538018 94556 538024
rect 95804 536518 95832 540110
rect 95792 536512 95844 536518
rect 95792 536454 95844 536460
rect 96448 534750 96476 540138
rect 97092 536858 97120 540138
rect 97736 539510 97764 540138
rect 97724 539504 97776 539510
rect 97724 539446 97776 539452
rect 98380 538218 98408 540138
rect 98368 538212 98420 538218
rect 98368 538154 98420 538160
rect 97908 537600 97960 537606
rect 97908 537542 97960 537548
rect 97080 536852 97132 536858
rect 97080 536794 97132 536800
rect 96436 534744 96488 534750
rect 96436 534686 96488 534692
rect 95148 533452 95200 533458
rect 95148 533394 95200 533400
rect 93872 528526 94084 528554
rect 93768 490612 93820 490618
rect 93768 490554 93820 490560
rect 93872 489954 93900 528526
rect 95160 499574 95188 533394
rect 97814 533352 97870 533361
rect 97814 533287 97870 533296
rect 95068 499546 95188 499574
rect 95068 491502 95096 499546
rect 96528 496120 96580 496126
rect 96528 496062 96580 496068
rect 95148 494760 95200 494766
rect 95148 494702 95200 494708
rect 95056 491496 95108 491502
rect 95054 491464 95056 491473
rect 95108 491464 95110 491473
rect 95054 491399 95110 491408
rect 94134 489968 94190 489977
rect 93872 489940 94134 489954
rect 93886 489926 94134 489940
rect 95160 489940 95188 494702
rect 96540 494290 96568 496062
rect 96528 494284 96580 494290
rect 96528 494226 96580 494232
rect 95790 493368 95846 493377
rect 95790 493303 95846 493312
rect 95804 489940 95832 493303
rect 97828 492658 97856 533287
rect 97816 492652 97868 492658
rect 97816 492594 97868 492600
rect 97724 491428 97776 491434
rect 97724 491370 97776 491376
rect 96436 491360 96488 491366
rect 96436 491302 96488 491308
rect 97078 491328 97134 491337
rect 96448 489940 96476 491302
rect 97078 491263 97134 491272
rect 97092 489940 97120 491263
rect 97736 489940 97764 491370
rect 97920 491298 97948 537542
rect 98380 536586 98408 538154
rect 99024 538014 99052 540138
rect 99668 539306 99696 540138
rect 99656 539300 99708 539306
rect 99656 539242 99708 539248
rect 99288 538892 99340 538898
rect 99288 538834 99340 538840
rect 99012 538008 99064 538014
rect 99012 537950 99064 537956
rect 98368 536580 98420 536586
rect 98368 536522 98420 536528
rect 99194 532264 99250 532273
rect 99194 532199 99250 532208
rect 98184 492652 98236 492658
rect 98184 492594 98236 492600
rect 98196 491366 98224 492594
rect 99208 492046 99236 532199
rect 99196 492040 99248 492046
rect 99196 491982 99248 491988
rect 99300 491722 99328 538834
rect 100312 538218 100340 540138
rect 100576 539300 100628 539306
rect 100576 539242 100628 539248
rect 100300 538212 100352 538218
rect 100300 538154 100352 538160
rect 99654 538112 99710 538121
rect 99654 538047 99710 538056
rect 99380 537532 99432 537538
rect 99380 537474 99432 537480
rect 99392 536761 99420 537474
rect 99472 536920 99524 536926
rect 99472 536862 99524 536868
rect 99378 536752 99434 536761
rect 99378 536687 99434 536696
rect 99484 536602 99512 536862
rect 99208 491694 99328 491722
rect 99392 536574 99512 536602
rect 99208 491502 99236 491694
rect 99288 491632 99340 491638
rect 99288 491574 99340 491580
rect 99196 491496 99248 491502
rect 99196 491438 99248 491444
rect 98368 491428 98420 491434
rect 98368 491370 98420 491376
rect 98184 491360 98236 491366
rect 98184 491302 98236 491308
rect 97908 491292 97960 491298
rect 97908 491234 97960 491240
rect 94134 489903 94190 489912
rect 73068 489874 73120 489880
rect 98196 489870 98224 491302
rect 98380 489940 98408 491370
rect 99208 489954 99236 491438
rect 99038 489926 99236 489954
rect 98184 489864 98236 489870
rect 98184 489806 98236 489812
rect 99196 489864 99248 489870
rect 99196 489806 99248 489812
rect 99208 489190 99236 489806
rect 99300 489258 99328 491574
rect 99288 489252 99340 489258
rect 99288 489194 99340 489200
rect 99196 489184 99248 489190
rect 99196 489126 99248 489132
rect 69308 460906 69704 460934
rect 69676 440042 69704 460906
rect 99392 442898 99420 536574
rect 99668 533338 99696 538047
rect 100312 536926 100340 538154
rect 100300 536920 100352 536926
rect 100300 536862 100352 536868
rect 99484 533310 99696 533338
rect 99484 446593 99512 533310
rect 99656 492108 99708 492114
rect 99656 492050 99708 492056
rect 99668 489940 99696 492050
rect 100588 466818 100616 539242
rect 100956 535362 100984 540138
rect 102227 540110 102272 540138
rect 102244 538150 102272 540110
rect 102232 538144 102284 538150
rect 102232 538086 102284 538092
rect 100944 535356 100996 535362
rect 100944 535298 100996 535304
rect 102048 535356 102100 535362
rect 102048 535298 102100 535304
rect 100668 491564 100720 491570
rect 100668 491506 100720 491512
rect 100680 491230 100708 491506
rect 100668 491224 100720 491230
rect 100668 491166 100720 491172
rect 100576 466812 100628 466818
rect 100576 466754 100628 466760
rect 100024 465792 100076 465798
rect 100024 465734 100076 465740
rect 99470 446584 99526 446593
rect 99470 446519 99526 446528
rect 99656 444372 99708 444378
rect 99656 444314 99708 444320
rect 99668 443873 99696 444314
rect 99654 443864 99710 443873
rect 99654 443799 99710 443808
rect 99746 443728 99802 443737
rect 99746 443663 99802 443672
rect 99392 442870 99512 442898
rect 99378 442368 99434 442377
rect 99378 442303 99434 442312
rect 99392 441590 99420 442303
rect 99288 441584 99340 441590
rect 99288 441526 99340 441532
rect 99380 441584 99432 441590
rect 99380 441526 99432 441532
rect 97908 440700 97960 440706
rect 97908 440642 97960 440648
rect 69676 440014 70058 440042
rect 69202 439104 69258 439113
rect 69202 439039 69258 439048
rect 69676 431954 69704 440014
rect 70688 432614 70716 440028
rect 71042 439104 71098 439113
rect 71042 439039 71098 439048
rect 70676 432608 70728 432614
rect 70676 432550 70728 432556
rect 69308 431926 69704 431954
rect 69204 397452 69256 397458
rect 69204 397394 69256 397400
rect 68928 394664 68980 394670
rect 68928 394606 68980 394612
rect 68940 393378 68968 394606
rect 68928 393372 68980 393378
rect 68928 393314 68980 393320
rect 68940 353161 68968 393314
rect 69110 380352 69166 380361
rect 69110 380287 69166 380296
rect 68926 353152 68982 353161
rect 68926 353087 68982 353096
rect 68940 352578 68968 353087
rect 68928 352572 68980 352578
rect 68928 352514 68980 352520
rect 68926 347304 68982 347313
rect 68926 347239 68982 347248
rect 68836 346384 68888 346390
rect 68834 346352 68836 346361
rect 68888 346352 68890 346361
rect 68834 346287 68890 346296
rect 68652 345092 68704 345098
rect 68652 345034 68704 345040
rect 68664 345001 68692 345034
rect 68650 344992 68706 345001
rect 68650 344927 68706 344936
rect 67638 343768 67694 343777
rect 67638 343703 67694 343712
rect 67652 343670 67680 343703
rect 67640 343664 67692 343670
rect 67640 343606 67692 343612
rect 67638 342952 67694 342961
rect 67638 342887 67694 342896
rect 67652 342310 67680 342887
rect 67640 342304 67692 342310
rect 67560 342264 67640 342292
rect 66996 338768 67048 338774
rect 66996 338710 67048 338716
rect 66904 327888 66956 327894
rect 66904 327830 66956 327836
rect 66168 318844 66220 318850
rect 66168 318786 66220 318792
rect 65524 299464 65576 299470
rect 65524 299406 65576 299412
rect 65984 295724 66036 295730
rect 65984 295666 66036 295672
rect 65996 262206 66024 295666
rect 66076 269136 66128 269142
rect 66076 269078 66128 269084
rect 65984 262200 66036 262206
rect 65984 262142 66036 262148
rect 65984 256760 66036 256766
rect 65984 256702 66036 256708
rect 65892 247172 65944 247178
rect 65892 247114 65944 247120
rect 64788 245744 64840 245750
rect 64788 245686 64840 245692
rect 64800 238066 64828 245686
rect 64788 238060 64840 238066
rect 64788 238002 64840 238008
rect 65904 204950 65932 247114
rect 65996 239426 66024 256702
rect 65984 239420 66036 239426
rect 65984 239362 66036 239368
rect 66088 225593 66116 269078
rect 66180 251190 66208 318786
rect 67364 302252 67416 302258
rect 67364 302194 67416 302200
rect 67376 261633 67404 302194
rect 67454 298888 67510 298897
rect 67454 298823 67510 298832
rect 67468 298353 67496 298823
rect 67454 298344 67510 298353
rect 67454 298279 67510 298288
rect 67468 283393 67496 298279
rect 67454 283384 67510 283393
rect 67454 283319 67510 283328
rect 67454 271960 67510 271969
rect 67454 271895 67510 271904
rect 67362 261624 67418 261633
rect 67362 261559 67418 261568
rect 66168 251184 66220 251190
rect 66168 251126 66220 251132
rect 67362 248704 67418 248713
rect 67362 248639 67418 248648
rect 67376 232558 67404 248639
rect 67364 232552 67416 232558
rect 67364 232494 67416 232500
rect 66074 225584 66130 225593
rect 66074 225519 66130 225528
rect 65892 204944 65944 204950
rect 65892 204886 65944 204892
rect 67468 198082 67496 271895
rect 67456 198076 67508 198082
rect 67456 198018 67508 198024
rect 67454 129296 67510 129305
rect 67454 129231 67510 129240
rect 65522 128072 65578 128081
rect 65522 128007 65578 128016
rect 65536 127022 65564 128007
rect 65524 127016 65576 127022
rect 65524 126958 65576 126964
rect 66166 125216 66222 125225
rect 66166 125151 66222 125160
rect 66074 123584 66130 123593
rect 66074 123519 66130 123528
rect 66088 122874 66116 123519
rect 66076 122868 66128 122874
rect 66076 122810 66128 122816
rect 65154 120864 65210 120873
rect 65154 120799 65210 120808
rect 65168 120154 65196 120799
rect 65156 120148 65208 120154
rect 65156 120090 65208 120096
rect 65982 102368 66038 102377
rect 65982 102303 66038 102312
rect 65996 84182 66024 102303
rect 66180 100774 66208 125151
rect 67362 122632 67418 122641
rect 67362 122567 67418 122576
rect 66168 100768 66220 100774
rect 66074 100736 66130 100745
rect 66168 100710 66220 100716
rect 66074 100671 66130 100680
rect 66088 88233 66116 100671
rect 67376 93838 67404 122567
rect 67468 94897 67496 129231
rect 67454 94888 67510 94897
rect 67454 94823 67510 94832
rect 67364 93832 67416 93838
rect 67364 93774 67416 93780
rect 66074 88224 66130 88233
rect 66074 88159 66130 88168
rect 65984 84176 66036 84182
rect 65984 84118 66036 84124
rect 66260 71052 66312 71058
rect 66260 70994 66312 71000
rect 64696 49700 64748 49706
rect 64696 49642 64748 49648
rect 64512 27600 64564 27606
rect 64512 27542 64564 27548
rect 63500 24200 63552 24206
rect 63500 24142 63552 24148
rect 63512 16574 63540 24142
rect 66272 16574 66300 70994
rect 67560 21418 67588 342264
rect 67640 342246 67692 342252
rect 67914 341728 67970 341737
rect 67914 341663 67970 341672
rect 68742 341728 68798 341737
rect 68742 341663 68798 341672
rect 67928 341562 67956 341663
rect 67916 341556 67968 341562
rect 67916 341498 67968 341504
rect 67638 341048 67694 341057
rect 67638 340983 67694 340992
rect 67652 340950 67680 340983
rect 67640 340944 67692 340950
rect 67640 340886 67692 340892
rect 67638 340232 67694 340241
rect 67638 340167 67694 340176
rect 67652 339590 67680 340167
rect 67640 339584 67692 339590
rect 67640 339526 67692 339532
rect 68756 305726 68784 341663
rect 68848 338842 68876 346287
rect 68940 339969 68968 347239
rect 68926 339960 68982 339969
rect 68926 339895 68982 339904
rect 68836 338836 68888 338842
rect 68836 338778 68888 338784
rect 69124 330750 69152 380287
rect 69216 363361 69244 397394
rect 69202 363352 69258 363361
rect 69202 363287 69258 363296
rect 69216 362982 69244 363287
rect 69204 362976 69256 362982
rect 69204 362918 69256 362924
rect 69308 340746 69336 431926
rect 70400 400988 70452 400994
rect 70400 400930 70452 400936
rect 70412 400314 70440 400930
rect 70400 400308 70452 400314
rect 70400 400250 70452 400256
rect 71056 389174 71084 439039
rect 71332 435402 71360 440028
rect 71780 439272 71832 439278
rect 71780 439214 71832 439220
rect 71320 435396 71372 435402
rect 71320 435338 71372 435344
rect 71688 406428 71740 406434
rect 71688 406370 71740 406376
rect 71700 405793 71728 406370
rect 71686 405784 71742 405793
rect 71686 405719 71742 405728
rect 71700 389366 71728 405719
rect 71688 389360 71740 389366
rect 71688 389302 71740 389308
rect 70964 389146 71084 389174
rect 69664 388544 69716 388550
rect 69664 388486 69716 388492
rect 69676 369170 69704 388486
rect 69756 388000 69808 388006
rect 69756 387942 69808 387948
rect 69768 385914 69796 387942
rect 69768 385886 70058 385914
rect 70964 385665 70992 389146
rect 71792 387870 71820 439214
rect 71976 438841 72004 440028
rect 72620 438938 72648 440028
rect 72608 438932 72660 438938
rect 72608 438874 72660 438880
rect 71962 438832 72018 438841
rect 71962 438767 72018 438776
rect 73264 438258 73292 440028
rect 73344 438932 73396 438938
rect 73344 438874 73396 438880
rect 73252 438252 73304 438258
rect 73252 438194 73304 438200
rect 73356 389842 73384 438874
rect 73908 438666 73936 440028
rect 73896 438660 73948 438666
rect 73896 438602 73948 438608
rect 74552 433294 74580 440028
rect 75184 439612 75236 439618
rect 75184 439554 75236 439560
rect 74724 434716 74776 434722
rect 74724 434658 74776 434664
rect 74540 433288 74592 433294
rect 74540 433230 74592 433236
rect 74630 407552 74686 407561
rect 74630 407487 74686 407496
rect 74540 400308 74592 400314
rect 74540 400250 74592 400256
rect 73344 389836 73396 389842
rect 73344 389778 73396 389784
rect 73344 389360 73396 389366
rect 73344 389302 73396 389308
rect 71780 387864 71832 387870
rect 71780 387806 71832 387812
rect 72700 387864 72752 387870
rect 72700 387806 72752 387812
rect 72712 385914 72740 387806
rect 73356 385914 73384 389302
rect 74552 389174 74580 400250
rect 74644 393314 74672 407487
rect 74736 394126 74764 434658
rect 75196 407561 75224 439554
rect 75840 434722 75868 440028
rect 76484 436082 76512 440028
rect 76472 436076 76524 436082
rect 76472 436018 76524 436024
rect 77128 435946 77156 440028
rect 77772 437345 77800 440028
rect 77298 437336 77354 437345
rect 77298 437271 77354 437280
rect 77758 437336 77814 437345
rect 77758 437271 77814 437280
rect 76012 435940 76064 435946
rect 76012 435882 76064 435888
rect 77116 435940 77168 435946
rect 77116 435882 77168 435888
rect 75828 434716 75880 434722
rect 75828 434658 75880 434664
rect 75182 407552 75238 407561
rect 75182 407487 75238 407496
rect 75196 407153 75224 407487
rect 75182 407144 75238 407153
rect 75182 407079 75238 407088
rect 75920 403640 75972 403646
rect 75920 403582 75972 403588
rect 75932 403102 75960 403582
rect 75920 403096 75972 403102
rect 75920 403038 75972 403044
rect 74724 394120 74776 394126
rect 74724 394062 74776 394068
rect 74644 393286 74856 393314
rect 74552 389146 74672 389174
rect 74644 385914 74672 389146
rect 72634 385886 72740 385914
rect 73278 385886 73384 385914
rect 74566 385886 74672 385914
rect 74828 385914 74856 393286
rect 75460 391264 75512 391270
rect 75460 391206 75512 391212
rect 75472 390658 75500 391206
rect 75460 390652 75512 390658
rect 75460 390594 75512 390600
rect 75472 385914 75500 390594
rect 75932 386050 75960 403038
rect 76024 386170 76052 435882
rect 77312 392698 77340 437271
rect 78416 437238 78444 440028
rect 78784 440014 79074 440042
rect 78784 438802 78812 440014
rect 78772 438796 78824 438802
rect 78772 438738 78824 438744
rect 77944 437232 77996 437238
rect 77944 437174 77996 437180
rect 78404 437232 78456 437238
rect 78404 437174 78456 437180
rect 77956 431254 77984 437174
rect 77944 431248 77996 431254
rect 77944 431190 77996 431196
rect 77300 392692 77352 392698
rect 77300 392634 77352 392640
rect 77484 388612 77536 388618
rect 77484 388554 77536 388560
rect 77300 388476 77352 388482
rect 77300 388418 77352 388424
rect 77312 388074 77340 388418
rect 77300 388068 77352 388074
rect 77300 388010 77352 388016
rect 76012 386164 76064 386170
rect 76012 386106 76064 386112
rect 75932 386022 76696 386050
rect 76668 385914 76696 386022
rect 77496 385914 77524 388554
rect 77956 387258 77984 431190
rect 78784 396778 78812 438738
rect 79704 437481 79732 440028
rect 78862 437472 78918 437481
rect 78862 437407 78918 437416
rect 79690 437472 79746 437481
rect 79690 437407 79746 437416
rect 78772 396772 78824 396778
rect 78772 396714 78824 396720
rect 78876 389881 78904 437407
rect 80992 437374 81020 440028
rect 81452 440014 81650 440042
rect 80980 437368 81032 437374
rect 80980 437310 81032 437316
rect 80992 436490 81020 437310
rect 80152 436484 80204 436490
rect 80152 436426 80204 436432
rect 80980 436484 81032 436490
rect 80980 436426 81032 436432
rect 80060 400920 80112 400926
rect 80060 400862 80112 400868
rect 80072 400246 80100 400862
rect 80060 400240 80112 400246
rect 80060 400182 80112 400188
rect 79324 390720 79376 390726
rect 79324 390662 79376 390668
rect 78862 389872 78918 389881
rect 78862 389807 78918 389816
rect 78496 388068 78548 388074
rect 78496 388010 78548 388016
rect 77944 387252 77996 387258
rect 77944 387194 77996 387200
rect 78508 385914 78536 388010
rect 74828 385886 75210 385914
rect 75472 385886 75854 385914
rect 76668 385886 77142 385914
rect 77496 385886 77786 385914
rect 78430 385886 78536 385914
rect 79336 385914 79364 390662
rect 80164 387190 80192 436426
rect 81452 436014 81480 440014
rect 82280 438734 82308 440028
rect 82820 439544 82872 439550
rect 82820 439486 82872 439492
rect 82832 438802 82860 439486
rect 82820 438796 82872 438802
rect 82820 438738 82872 438744
rect 82268 438728 82320 438734
rect 82268 438670 82320 438676
rect 82924 437306 82952 440028
rect 83464 438796 83516 438802
rect 83464 438738 83516 438744
rect 82912 437300 82964 437306
rect 82912 437242 82964 437248
rect 81440 436008 81492 436014
rect 81440 435950 81492 435956
rect 80244 400240 80296 400246
rect 80244 400182 80296 400188
rect 80152 387184 80204 387190
rect 80152 387126 80204 387132
rect 80256 386414 80284 400182
rect 81452 399634 81480 435950
rect 82924 431954 82952 437242
rect 82832 431926 82952 431954
rect 81440 399628 81492 399634
rect 81440 399570 81492 399576
rect 82832 394058 82860 431926
rect 83476 396846 83504 438738
rect 83568 438190 83596 440028
rect 84212 438977 84240 440028
rect 84198 438968 84254 438977
rect 84198 438903 84254 438912
rect 83556 438184 83608 438190
rect 83556 438126 83608 438132
rect 84856 435985 84884 440028
rect 86158 440014 86264 440042
rect 85486 438968 85542 438977
rect 85542 438926 85620 438954
rect 85486 438903 85542 438912
rect 84290 435976 84346 435985
rect 84290 435911 84346 435920
rect 84842 435976 84898 435985
rect 84842 435911 84898 435920
rect 83464 396840 83516 396846
rect 83464 396782 83516 396788
rect 82820 394052 82872 394058
rect 82820 393994 82872 394000
rect 81440 393984 81492 393990
rect 81440 393926 81492 393932
rect 83002 393952 83058 393961
rect 81452 388006 81480 393926
rect 83002 393887 83058 393896
rect 83016 393514 83044 393887
rect 83004 393508 83056 393514
rect 83004 393450 83056 393456
rect 82912 392148 82964 392154
rect 82912 392090 82964 392096
rect 82924 391950 82952 392090
rect 82912 391944 82964 391950
rect 82912 391886 82964 391892
rect 81440 388000 81492 388006
rect 81440 387942 81492 387948
rect 82544 388000 82596 388006
rect 82544 387942 82596 387948
rect 80612 386504 80664 386510
rect 80612 386446 80664 386452
rect 80256 386386 80468 386414
rect 80440 385914 80468 386386
rect 79336 385886 79718 385914
rect 80362 385886 80468 385914
rect 80624 385914 80652 386446
rect 82556 385914 82584 387942
rect 83016 385914 83044 393450
rect 83648 392148 83700 392154
rect 83648 392090 83700 392096
rect 83660 385914 83688 392090
rect 84304 386034 84332 435911
rect 85592 431954 85620 438926
rect 86236 437345 86264 440014
rect 86788 437510 86816 440028
rect 87432 438802 87460 440028
rect 88090 440014 88288 440042
rect 87420 438796 87472 438802
rect 87420 438738 87472 438744
rect 86776 437504 86828 437510
rect 87604 437504 87656 437510
rect 86776 437446 86828 437452
rect 87602 437472 87604 437481
rect 87656 437472 87658 437481
rect 87602 437407 87658 437416
rect 86222 437336 86278 437345
rect 86222 437271 86278 437280
rect 85592 431926 85804 431954
rect 85670 401704 85726 401713
rect 85670 401639 85726 401648
rect 84936 399492 84988 399498
rect 84936 399434 84988 399440
rect 84948 390697 84976 399434
rect 84934 390688 84990 390697
rect 84934 390623 84990 390632
rect 84948 389174 84976 390623
rect 84948 389146 85160 389174
rect 84476 386572 84528 386578
rect 84476 386514 84528 386520
rect 84292 386028 84344 386034
rect 84292 385970 84344 385976
rect 80624 385886 81006 385914
rect 82294 385886 82584 385914
rect 82938 385886 83044 385914
rect 83582 385886 83688 385914
rect 84488 385914 84516 386514
rect 85132 385914 85160 389146
rect 85684 385914 85712 401639
rect 85776 398206 85804 431926
rect 85764 398200 85816 398206
rect 85764 398142 85816 398148
rect 86236 392630 86264 437271
rect 87616 398138 87644 437407
rect 88260 437374 88288 440014
rect 88720 439142 88748 440028
rect 88996 440014 89378 440042
rect 88708 439136 88760 439142
rect 88708 439078 88760 439084
rect 88248 437368 88300 437374
rect 88248 437310 88300 437316
rect 88260 402257 88288 437310
rect 88996 437306 89024 440014
rect 90008 438190 90036 440028
rect 91296 438802 91324 440028
rect 91284 438796 91336 438802
rect 91284 438738 91336 438744
rect 91008 438592 91060 438598
rect 91008 438534 91060 438540
rect 91020 438190 91048 438534
rect 89996 438184 90048 438190
rect 89996 438126 90048 438132
rect 91008 438184 91060 438190
rect 91008 438126 91060 438132
rect 88984 437300 89036 437306
rect 88984 437242 89036 437248
rect 88246 402248 88302 402257
rect 88246 402183 88302 402192
rect 88064 399560 88116 399566
rect 88064 399502 88116 399508
rect 88076 399022 88104 399502
rect 87696 399016 87748 399022
rect 87696 398958 87748 398964
rect 88064 399016 88116 399022
rect 88064 398958 88116 398964
rect 87604 398132 87656 398138
rect 87604 398074 87656 398080
rect 86224 392624 86276 392630
rect 86224 392566 86276 392572
rect 86960 388000 87012 388006
rect 86960 387942 87012 387948
rect 86972 387190 87000 387942
rect 87052 387932 87104 387938
rect 87052 387874 87104 387880
rect 86960 387184 87012 387190
rect 86960 387126 87012 387132
rect 87064 385914 87092 387874
rect 87708 385914 87736 398958
rect 88340 398132 88392 398138
rect 88340 398074 88392 398080
rect 88352 385914 88380 398074
rect 88996 393314 89024 437242
rect 89720 410576 89772 410582
rect 89720 410518 89772 410524
rect 89732 409902 89760 410518
rect 89720 409896 89772 409902
rect 89720 409838 89772 409844
rect 88904 393286 89024 393314
rect 88904 388550 88932 393286
rect 88984 392216 89036 392222
rect 88984 392158 89036 392164
rect 88996 391270 89024 392158
rect 88984 391264 89036 391270
rect 88984 391206 89036 391212
rect 88892 388544 88944 388550
rect 88892 388486 88944 388492
rect 89732 385914 89760 409838
rect 89812 406428 89864 406434
rect 89812 406370 89864 406376
rect 89824 402974 89852 406370
rect 89824 402946 90312 402974
rect 90284 385914 90312 402946
rect 91020 392630 91048 438126
rect 91940 436014 91968 440028
rect 92584 439090 92612 440028
rect 92400 439062 92612 439090
rect 91928 436008 91980 436014
rect 91928 435950 91980 435956
rect 92400 404977 92428 439062
rect 92480 439000 92532 439006
rect 92480 438942 92532 438948
rect 92492 405074 92520 438942
rect 92584 438705 92612 439062
rect 93228 439006 93256 440028
rect 93216 439000 93268 439006
rect 93216 438942 93268 438948
rect 92570 438696 92626 438705
rect 92570 438631 92626 438640
rect 93872 438530 93900 440028
rect 94516 439074 94544 440028
rect 94504 439068 94556 439074
rect 94504 439010 94556 439016
rect 95160 438682 95188 440028
rect 96448 439210 96476 440028
rect 97106 440014 97488 440042
rect 96436 439204 96488 439210
rect 96436 439146 96488 439152
rect 96448 438734 96476 439146
rect 95068 438654 95188 438682
rect 96436 438728 96488 438734
rect 96436 438670 96488 438676
rect 93860 438524 93912 438530
rect 93860 438466 93912 438472
rect 95068 436082 95096 438654
rect 95148 438524 95200 438530
rect 95148 438466 95200 438472
rect 95056 436076 95108 436082
rect 95056 436018 95108 436024
rect 92480 405068 92532 405074
rect 92480 405010 92532 405016
rect 92386 404968 92442 404977
rect 92386 404903 92442 404912
rect 95068 398206 95096 436018
rect 95056 398200 95108 398206
rect 95056 398142 95108 398148
rect 93952 396772 94004 396778
rect 93952 396714 94004 396720
rect 91008 392624 91060 392630
rect 91008 392566 91060 392572
rect 92848 388068 92900 388074
rect 92848 388010 92900 388016
rect 91560 387932 91612 387938
rect 91560 387874 91612 387880
rect 91572 385914 91600 387874
rect 92860 385914 92888 388010
rect 93308 388000 93360 388006
rect 93308 387942 93360 387948
rect 84488 385886 84870 385914
rect 85132 385886 85514 385914
rect 85684 385886 86158 385914
rect 87064 385886 87446 385914
rect 87708 385886 88090 385914
rect 88352 385886 88734 385914
rect 89732 385886 90022 385914
rect 90284 385886 90666 385914
rect 91310 385886 91600 385914
rect 92598 385886 92888 385914
rect 70950 385656 71006 385665
rect 70702 385614 70950 385642
rect 70950 385591 71006 385600
rect 93320 385370 93348 387942
rect 93964 385914 93992 396714
rect 95160 393961 95188 438466
rect 97460 437442 97488 440014
rect 97736 439929 97764 440028
rect 97722 439920 97778 439929
rect 97722 439855 97778 439864
rect 97736 438054 97764 439855
rect 97724 438048 97776 438054
rect 97724 437990 97776 437996
rect 97448 437436 97500 437442
rect 97448 437378 97500 437384
rect 97460 431954 97488 437378
rect 97460 431926 97856 431954
rect 95884 399492 95936 399498
rect 95884 399434 95936 399440
rect 95792 393984 95844 393990
rect 95146 393952 95202 393961
rect 95792 393926 95844 393932
rect 95146 393887 95202 393896
rect 95516 389224 95568 389230
rect 95516 389166 95568 389172
rect 94872 388612 94924 388618
rect 94872 388554 94924 388560
rect 94884 385914 94912 388554
rect 95424 388136 95476 388142
rect 95424 388078 95476 388084
rect 93886 385886 93992 385914
rect 94530 385886 94912 385914
rect 95436 385694 95464 388078
rect 95528 385914 95556 389166
rect 95804 386186 95832 393926
rect 95896 388074 95924 399434
rect 97828 396846 97856 431926
rect 97920 397882 97948 440642
rect 98380 437889 98408 440028
rect 99024 438666 99052 440028
rect 99012 438660 99064 438666
rect 99012 438602 99064 438608
rect 98644 438048 98696 438054
rect 98644 437990 98696 437996
rect 98366 437880 98422 437889
rect 98366 437815 98422 437824
rect 98656 400897 98684 437990
rect 99300 437889 99328 441526
rect 99484 441153 99512 442870
rect 99470 441144 99526 441153
rect 99470 441079 99526 441088
rect 99668 438870 99696 440028
rect 99656 438864 99708 438870
rect 99656 438806 99708 438812
rect 99760 438462 99788 443663
rect 100036 438598 100064 465734
rect 100024 438592 100076 438598
rect 100024 438534 100076 438540
rect 99748 438456 99800 438462
rect 99748 438398 99800 438404
rect 99286 437880 99342 437889
rect 99286 437815 99342 437824
rect 99300 407833 99328 437815
rect 99286 407824 99342 407833
rect 99286 407759 99342 407768
rect 98642 400888 98698 400897
rect 98642 400823 98698 400832
rect 97920 397854 98040 397882
rect 98012 397497 98040 397854
rect 97998 397488 98054 397497
rect 97998 397423 98054 397432
rect 97816 396840 97868 396846
rect 97816 396782 97868 396788
rect 96712 395344 96764 395350
rect 96712 395286 96764 395292
rect 95884 388068 95936 388074
rect 95884 388010 95936 388016
rect 95804 386158 96016 386186
rect 95988 385914 96016 386158
rect 96724 385914 96752 395286
rect 98012 385914 98040 397423
rect 100680 394058 100708 491166
rect 101404 490680 101456 490686
rect 101404 490622 101456 490628
rect 101312 458856 101364 458862
rect 101312 458798 101364 458804
rect 101324 458153 101352 458798
rect 101310 458144 101366 458153
rect 101310 458079 101366 458088
rect 101126 400344 101182 400353
rect 101126 400279 101182 400288
rect 100668 394052 100720 394058
rect 100668 393994 100720 394000
rect 101036 392216 101088 392222
rect 101036 392158 101088 392164
rect 99288 389836 99340 389842
rect 99288 389778 99340 389784
rect 99300 385914 99328 389778
rect 100022 388376 100078 388385
rect 100022 388311 100078 388320
rect 100036 385914 100064 388311
rect 101048 385914 101076 392158
rect 95528 385886 95818 385914
rect 95988 385886 96462 385914
rect 96724 385886 97106 385914
rect 98012 385886 98394 385914
rect 99038 385886 99328 385914
rect 99682 385886 100064 385914
rect 100970 385886 101076 385914
rect 101140 385914 101168 400279
rect 101416 392222 101444 490622
rect 101956 471300 102008 471306
rect 101956 471242 102008 471248
rect 101968 470257 101996 471242
rect 101954 470248 102010 470257
rect 101954 470183 102010 470192
rect 101496 466812 101548 466818
rect 101496 466754 101548 466760
rect 101508 440298 101536 466754
rect 101586 451208 101642 451217
rect 101586 451143 101642 451152
rect 101600 448662 101628 451143
rect 101588 448656 101640 448662
rect 101588 448598 101640 448604
rect 101496 440292 101548 440298
rect 101496 440234 101548 440240
rect 101600 429894 101628 448598
rect 102060 441697 102088 535298
rect 102888 534070 102916 540138
rect 103244 538960 103296 538966
rect 103244 538902 103296 538908
rect 102876 534064 102928 534070
rect 102876 534006 102928 534012
rect 102692 491292 102744 491298
rect 102692 491234 102744 491240
rect 102414 485344 102470 485353
rect 102414 485279 102470 485288
rect 102138 485208 102194 485217
rect 102138 485143 102140 485152
rect 102192 485143 102194 485152
rect 102140 485114 102192 485120
rect 102428 485110 102456 485279
rect 102416 485104 102468 485110
rect 102416 485046 102468 485052
rect 102140 482792 102192 482798
rect 102140 482734 102192 482740
rect 102152 482633 102180 482734
rect 102138 482624 102194 482633
rect 102138 482559 102194 482568
rect 102704 481710 102732 491234
rect 102782 487248 102838 487257
rect 102782 487183 102838 487192
rect 102796 487150 102824 487183
rect 102784 487144 102836 487150
rect 102784 487086 102836 487092
rect 102692 481704 102744 481710
rect 102692 481646 102744 481652
rect 102140 481636 102192 481642
rect 102140 481578 102192 481584
rect 102152 481137 102180 481578
rect 102232 481568 102284 481574
rect 102232 481510 102284 481516
rect 102138 481128 102194 481137
rect 102138 481063 102194 481072
rect 102244 480593 102272 481510
rect 102230 480584 102286 480593
rect 102230 480519 102286 480528
rect 102140 480208 102192 480214
rect 102140 480150 102192 480156
rect 102152 479913 102180 480150
rect 102138 479904 102194 479913
rect 102138 479839 102194 479848
rect 102140 477420 102192 477426
rect 102140 477362 102192 477368
rect 102152 477057 102180 477362
rect 102232 477352 102284 477358
rect 102232 477294 102284 477300
rect 102138 477048 102194 477057
rect 102138 476983 102194 476992
rect 102244 476513 102272 477294
rect 102322 477184 102378 477193
rect 102322 477119 102378 477128
rect 102230 476504 102286 476513
rect 102230 476439 102286 476448
rect 102336 476066 102364 477119
rect 102324 476060 102376 476066
rect 102324 476002 102376 476008
rect 102138 475688 102194 475697
rect 102138 475623 102194 475632
rect 102152 475386 102180 475623
rect 102140 475380 102192 475386
rect 102140 475322 102192 475328
rect 102138 475008 102194 475017
rect 102138 474943 102194 474952
rect 102152 474774 102180 474943
rect 102140 474768 102192 474774
rect 102140 474710 102192 474716
rect 102232 474700 102284 474706
rect 102232 474642 102284 474648
rect 102244 474337 102272 474642
rect 102230 474328 102286 474337
rect 102230 474263 102286 474272
rect 102138 472968 102194 472977
rect 102138 472903 102194 472912
rect 102152 472666 102180 472903
rect 102140 472660 102192 472666
rect 102140 472602 102192 472608
rect 102138 472288 102194 472297
rect 102138 472223 102194 472232
rect 102152 472122 102180 472223
rect 102140 472116 102192 472122
rect 102140 472058 102192 472064
rect 102140 471980 102192 471986
rect 102140 471922 102192 471928
rect 102152 471617 102180 471922
rect 102138 471608 102194 471617
rect 102138 471543 102194 471552
rect 102138 470928 102194 470937
rect 102138 470863 102194 470872
rect 102152 470626 102180 470863
rect 102140 470620 102192 470626
rect 102140 470562 102192 470568
rect 102140 469872 102192 469878
rect 102140 469814 102192 469820
rect 102152 469577 102180 469814
rect 102138 469568 102194 469577
rect 102138 469503 102194 469512
rect 102140 469192 102192 469198
rect 102140 469134 102192 469140
rect 102152 468897 102180 469134
rect 102138 468888 102194 468897
rect 102138 468823 102194 468832
rect 102140 467832 102192 467838
rect 102140 467774 102192 467780
rect 102152 467537 102180 467774
rect 102232 467764 102284 467770
rect 102232 467706 102284 467712
rect 102138 467528 102194 467537
rect 102138 467463 102194 467472
rect 102244 466993 102272 467706
rect 102230 466984 102286 466993
rect 102230 466919 102286 466928
rect 102230 466168 102286 466177
rect 102230 466103 102286 466112
rect 102244 465118 102272 466103
rect 102324 465724 102376 465730
rect 102324 465666 102376 465672
rect 102232 465112 102284 465118
rect 102232 465054 102284 465060
rect 102140 465044 102192 465050
rect 102140 464986 102192 464992
rect 102152 464273 102180 464986
rect 102336 464953 102364 465666
rect 102322 464944 102378 464953
rect 102322 464879 102378 464888
rect 102138 464264 102194 464273
rect 102138 464199 102194 464208
rect 102140 463684 102192 463690
rect 102140 463626 102192 463632
rect 102152 463457 102180 463626
rect 102138 463448 102194 463457
rect 102138 463383 102194 463392
rect 102232 462324 102284 462330
rect 102232 462266 102284 462272
rect 102140 462256 102192 462262
rect 102140 462198 102192 462204
rect 102152 462097 102180 462198
rect 102138 462088 102194 462097
rect 102138 462023 102194 462032
rect 102244 461553 102272 462266
rect 102230 461544 102286 461553
rect 102230 461479 102286 461488
rect 102140 460896 102192 460902
rect 102140 460838 102192 460844
rect 102152 460737 102180 460838
rect 102138 460728 102194 460737
rect 102138 460663 102194 460672
rect 102140 460216 102192 460222
rect 102140 460158 102192 460164
rect 102152 460057 102180 460158
rect 102138 460048 102194 460057
rect 102138 459983 102194 459992
rect 103256 459610 103284 538902
rect 103532 537946 103560 540138
rect 103704 539980 103756 539986
rect 103704 539922 103756 539928
rect 103520 537940 103572 537946
rect 103520 537882 103572 537888
rect 103716 537606 103744 539922
rect 104176 539374 104204 540138
rect 104820 539889 104848 540138
rect 105648 540002 105676 540382
rect 105464 539974 105676 540002
rect 104806 539880 104862 539889
rect 104806 539815 104862 539824
rect 104164 539368 104216 539374
rect 104164 539310 104216 539316
rect 104716 539368 104768 539374
rect 104716 539310 104768 539316
rect 103704 537600 103756 537606
rect 103704 537542 103756 537548
rect 104162 536888 104218 536897
rect 104162 536823 104218 536832
rect 103520 490612 103572 490618
rect 103520 490554 103572 490560
rect 103426 488608 103482 488617
rect 103426 488543 103428 488552
rect 103480 488543 103482 488552
rect 103428 488514 103480 488520
rect 103336 488504 103388 488510
rect 103336 488446 103388 488452
rect 103348 487393 103376 488446
rect 103426 487928 103482 487937
rect 103426 487863 103482 487872
rect 103334 487384 103390 487393
rect 103334 487319 103390 487328
rect 103440 487286 103468 487863
rect 103428 487280 103480 487286
rect 103428 487222 103480 487228
rect 103336 487076 103388 487082
rect 103336 487018 103388 487024
rect 103348 486577 103376 487018
rect 103334 486568 103390 486577
rect 103334 486503 103390 486512
rect 103426 477728 103482 477737
rect 103426 477663 103482 477672
rect 103440 477494 103468 477663
rect 103428 477488 103480 477494
rect 103428 477430 103480 477436
rect 103336 476060 103388 476066
rect 103336 476002 103388 476008
rect 102232 459604 102284 459610
rect 102232 459546 102284 459552
rect 103244 459604 103296 459610
rect 103244 459546 103296 459552
rect 102140 459536 102192 459542
rect 102140 459478 102192 459484
rect 102152 459377 102180 459478
rect 102138 459368 102194 459377
rect 102138 459303 102194 459312
rect 102244 458833 102272 459546
rect 102230 458824 102286 458833
rect 102230 458759 102286 458768
rect 102232 457564 102284 457570
rect 102232 457506 102284 457512
rect 102244 455433 102272 457506
rect 102874 456104 102930 456113
rect 102874 456039 102876 456048
rect 102928 456039 102930 456048
rect 102876 456010 102928 456016
rect 102230 455424 102286 455433
rect 102140 455388 102192 455394
rect 102230 455359 102286 455368
rect 102140 455330 102192 455336
rect 102152 454753 102180 455330
rect 102138 454744 102194 454753
rect 102138 454679 102194 454688
rect 102140 454028 102192 454034
rect 102140 453970 102192 453976
rect 102152 453257 102180 453970
rect 102874 453384 102930 453393
rect 102874 453319 102876 453328
rect 102928 453319 102930 453328
rect 102876 453290 102928 453296
rect 102138 453248 102194 453257
rect 102138 453183 102194 453192
rect 102322 452024 102378 452033
rect 102322 451959 102378 451968
rect 102336 451926 102364 451959
rect 102324 451920 102376 451926
rect 102324 451862 102376 451868
rect 102140 451308 102192 451314
rect 102140 451250 102192 451256
rect 102152 450673 102180 451250
rect 102138 450664 102194 450673
rect 102138 450599 102194 450608
rect 102140 449880 102192 449886
rect 102140 449822 102192 449828
rect 102152 449177 102180 449822
rect 102874 449304 102930 449313
rect 102874 449239 102876 449248
rect 102928 449239 102930 449248
rect 102876 449210 102928 449216
rect 102138 449168 102194 449177
rect 102138 449103 102194 449112
rect 102140 448520 102192 448526
rect 102140 448462 102192 448468
rect 102230 448488 102286 448497
rect 102152 447953 102180 448462
rect 102230 448423 102286 448432
rect 102138 447944 102194 447953
rect 102138 447879 102194 447888
rect 102244 447166 102272 448423
rect 102232 447160 102284 447166
rect 102232 447102 102284 447108
rect 102598 446584 102654 446593
rect 102598 446519 102654 446528
rect 102612 445806 102640 446519
rect 102600 445800 102652 445806
rect 102506 445768 102562 445777
rect 102600 445742 102652 445748
rect 102506 445703 102562 445712
rect 103244 445732 103296 445738
rect 102520 445670 102548 445703
rect 103244 445674 103296 445680
rect 102508 445664 102560 445670
rect 102508 445606 102560 445612
rect 103256 445233 103284 445674
rect 103242 445224 103298 445233
rect 103242 445159 103298 445168
rect 102232 445052 102284 445058
rect 102232 444994 102284 445000
rect 102244 443737 102272 444994
rect 102230 443728 102286 443737
rect 102230 443663 102286 443672
rect 102874 443048 102930 443057
rect 102874 442983 102930 442992
rect 102888 442270 102916 442983
rect 102876 442264 102928 442270
rect 102876 442206 102928 442212
rect 102046 441688 102102 441697
rect 102046 441623 102102 441632
rect 102598 441144 102654 441153
rect 102598 441079 102654 441088
rect 102612 440366 102640 441079
rect 102600 440360 102652 440366
rect 102600 440302 102652 440308
rect 102048 440292 102100 440298
rect 102048 440234 102100 440240
rect 102060 439793 102088 440234
rect 102046 439784 102102 439793
rect 102046 439719 102102 439728
rect 101588 429888 101640 429894
rect 101588 429830 101640 429836
rect 102230 395312 102286 395321
rect 102230 395247 102286 395256
rect 101404 392216 101456 392222
rect 101404 392158 101456 392164
rect 102244 388618 102272 395247
rect 103348 390114 103376 476002
rect 103440 391241 103468 477430
rect 103532 438530 103560 490554
rect 104072 471504 104124 471510
rect 104072 471446 104124 471452
rect 104084 465633 104112 471446
rect 104070 465624 104126 465633
rect 104070 465559 104126 465568
rect 103612 457496 103664 457502
rect 103612 457438 103664 457444
rect 103624 455977 103652 457438
rect 103610 455968 103666 455977
rect 103610 455903 103666 455912
rect 104176 445670 104204 536823
rect 104728 528554 104756 539310
rect 104820 536897 104848 539815
rect 105464 538121 105492 539974
rect 105544 539912 105596 539918
rect 105544 539854 105596 539860
rect 105450 538112 105506 538121
rect 105450 538047 105506 538056
rect 104806 536888 104862 536897
rect 104806 536823 104862 536832
rect 104728 528526 104848 528554
rect 104820 445874 104848 528526
rect 104900 487212 104952 487218
rect 104900 487154 104952 487160
rect 104912 487082 104940 487154
rect 104900 487076 104952 487082
rect 104900 487018 104952 487024
rect 105556 482798 105584 539854
rect 105636 539028 105688 539034
rect 105636 538970 105688 538976
rect 105544 482792 105596 482798
rect 105544 482734 105596 482740
rect 104900 481704 104952 481710
rect 104900 481646 104952 481652
rect 104808 445868 104860 445874
rect 104808 445810 104860 445816
rect 104820 445738 104848 445810
rect 104808 445732 104860 445738
rect 104808 445674 104860 445680
rect 104164 445664 104216 445670
rect 104164 445606 104216 445612
rect 103520 438524 103572 438530
rect 103520 438466 103572 438472
rect 103612 391264 103664 391270
rect 103426 391232 103482 391241
rect 103612 391206 103664 391212
rect 103426 391167 103482 391176
rect 103336 390108 103388 390114
rect 103336 390050 103388 390056
rect 103624 389162 103652 391206
rect 103612 389156 103664 389162
rect 103612 389098 103664 389104
rect 102232 388612 102284 388618
rect 102232 388554 102284 388560
rect 102600 388544 102652 388550
rect 102600 388486 102652 388492
rect 102612 385914 102640 388486
rect 103624 385914 103652 389098
rect 104176 387025 104204 445606
rect 104912 437306 104940 481646
rect 105542 479088 105598 479097
rect 105542 479023 105598 479032
rect 105556 478990 105584 479023
rect 105544 478984 105596 478990
rect 105544 478926 105596 478932
rect 105648 448526 105676 538970
rect 105740 487218 105768 567166
rect 105820 555144 105872 555150
rect 105820 555086 105872 555092
rect 105832 539918 105860 555086
rect 105820 539912 105872 539918
rect 105820 539854 105872 539860
rect 105818 539608 105874 539617
rect 105818 539543 105874 539552
rect 105832 539034 105860 539543
rect 105820 539028 105872 539034
rect 105820 538970 105872 538976
rect 106292 538121 106320 625126
rect 106922 587888 106978 587897
rect 106922 587823 106978 587832
rect 106936 586566 106964 587823
rect 106924 586560 106976 586566
rect 106924 586502 106976 586508
rect 106936 584526 106964 586502
rect 107016 585268 107068 585274
rect 107016 585210 107068 585216
rect 106924 584520 106976 584526
rect 106924 584462 106976 584468
rect 106924 583772 106976 583778
rect 106924 583714 106976 583720
rect 106936 575113 106964 583714
rect 107028 577697 107056 585210
rect 107580 582729 107608 632946
rect 108960 586514 108988 634786
rect 108776 586486 108988 586514
rect 107566 582720 107622 582729
rect 107566 582655 107622 582664
rect 107108 582548 107160 582554
rect 107108 582490 107160 582496
rect 107014 577688 107070 577697
rect 107014 577623 107070 577632
rect 106922 575104 106978 575113
rect 106922 575039 106978 575048
rect 107120 574705 107148 582490
rect 108028 580984 108080 580990
rect 108028 580926 108080 580932
rect 108040 580281 108068 580926
rect 108026 580272 108082 580281
rect 108026 580207 108082 580216
rect 108670 578776 108726 578785
rect 108670 578711 108726 578720
rect 108684 578270 108712 578711
rect 108672 578264 108724 578270
rect 108118 578232 108174 578241
rect 108672 578206 108724 578212
rect 108118 578167 108120 578176
rect 108172 578167 108174 578176
rect 108120 578138 108172 578144
rect 108776 576745 108804 586486
rect 108946 580952 109002 580961
rect 108946 580887 108948 580896
rect 109000 580887 109002 580896
rect 108948 580858 109000 580864
rect 108948 579624 109000 579630
rect 108946 579592 108948 579601
rect 109000 579592 109002 579601
rect 108946 579527 109002 579536
rect 108946 577552 109002 577561
rect 108946 577487 108948 577496
rect 109000 577487 109002 577496
rect 108948 577458 109000 577464
rect 108762 576736 108818 576745
rect 108762 576671 108818 576680
rect 108672 576224 108724 576230
rect 108670 576192 108672 576201
rect 108724 576192 108726 576201
rect 108776 576162 108804 576671
rect 108670 576127 108726 576136
rect 108764 576156 108816 576162
rect 108764 576098 108816 576104
rect 107106 574696 107162 574705
rect 107106 574631 107162 574640
rect 108580 574048 108632 574054
rect 108580 573990 108632 573996
rect 108946 574016 109002 574025
rect 108592 572801 108620 573990
rect 108946 573951 108948 573960
rect 109000 573951 109002 573960
rect 108948 573922 109000 573928
rect 108946 573336 109002 573345
rect 108946 573271 109002 573280
rect 108960 573238 108988 573271
rect 108948 573232 109000 573238
rect 108948 573174 109000 573180
rect 107382 572792 107438 572801
rect 107382 572727 107438 572736
rect 108578 572792 108634 572801
rect 108578 572727 108634 572736
rect 106740 551268 106792 551274
rect 106740 551210 106792 551216
rect 106752 551041 106780 551210
rect 106370 551032 106426 551041
rect 106370 550967 106426 550976
rect 106738 551032 106794 551041
rect 106738 550967 106794 550976
rect 106384 538966 106412 550967
rect 106372 538960 106424 538966
rect 106372 538902 106424 538908
rect 106278 538112 106334 538121
rect 106278 538047 106334 538056
rect 107292 489252 107344 489258
rect 107292 489194 107344 489200
rect 105728 487212 105780 487218
rect 105728 487154 105780 487160
rect 106922 486024 106978 486033
rect 106922 485959 106978 485968
rect 106186 478952 106242 478961
rect 106186 478887 106242 478896
rect 106200 467906 106228 478887
rect 106188 467900 106240 467906
rect 106188 467842 106240 467848
rect 106200 467770 106228 467842
rect 106188 467764 106240 467770
rect 106188 467706 106240 467712
rect 106556 463412 106608 463418
rect 106556 463354 106608 463360
rect 106188 463004 106240 463010
rect 106188 462946 106240 462952
rect 106200 462262 106228 462946
rect 106188 462256 106240 462262
rect 106188 462198 106240 462204
rect 106568 460970 106596 463354
rect 106556 460964 106608 460970
rect 106556 460906 106608 460912
rect 106096 460216 106148 460222
rect 106096 460158 106148 460164
rect 106004 448724 106056 448730
rect 106004 448666 106056 448672
rect 106016 448526 106044 448666
rect 105636 448520 105688 448526
rect 105636 448462 105688 448468
rect 106004 448520 106056 448526
rect 106004 448462 106056 448468
rect 105544 440292 105596 440298
rect 105544 440234 105596 440240
rect 104900 437300 104952 437306
rect 104900 437242 104952 437248
rect 105556 395457 105584 440234
rect 106108 405006 106136 460158
rect 106188 449268 106240 449274
rect 106188 449210 106240 449216
rect 106096 405000 106148 405006
rect 106096 404942 106148 404948
rect 105542 395448 105598 395457
rect 105542 395383 105598 395392
rect 106200 393314 106228 449210
rect 106936 398886 106964 485959
rect 106280 398880 106332 398886
rect 106280 398822 106332 398828
rect 106924 398880 106976 398886
rect 106924 398822 106976 398828
rect 106108 393286 106228 393314
rect 104624 388612 104676 388618
rect 104624 388554 104676 388560
rect 104162 387016 104218 387025
rect 104162 386951 104218 386960
rect 101140 385886 101614 385914
rect 102258 385886 102640 385914
rect 103546 385886 103652 385914
rect 104636 385778 104664 388554
rect 106108 386102 106136 393286
rect 106188 392692 106240 392698
rect 106188 392634 106240 392640
rect 106096 386096 106148 386102
rect 106096 386038 106148 386044
rect 106200 385914 106228 392634
rect 106122 385886 106228 385914
rect 106292 385914 106320 398822
rect 107304 393314 107332 489194
rect 107396 481574 107424 572727
rect 108028 572008 108080 572014
rect 108028 571950 108080 571956
rect 108302 571976 108358 571985
rect 108040 571441 108068 571950
rect 108302 571911 108358 571920
rect 108026 571432 108082 571441
rect 108026 571367 108082 571376
rect 108316 571334 108344 571911
rect 108304 571328 108356 571334
rect 108304 571270 108356 571276
rect 107474 560552 107530 560561
rect 107474 560487 107530 560496
rect 107384 481568 107436 481574
rect 107384 481510 107436 481516
rect 107384 478916 107436 478922
rect 107384 478858 107436 478864
rect 107396 449954 107424 478858
rect 107488 469266 107516 560487
rect 108026 559056 108082 559065
rect 108026 558991 108082 559000
rect 108040 558890 108068 558991
rect 108028 558884 108080 558890
rect 108028 558826 108080 558832
rect 107752 558816 107804 558822
rect 107752 558758 107804 558764
rect 107764 557841 107792 558758
rect 108040 558521 108068 558826
rect 108026 558512 108082 558521
rect 108026 558447 108082 558456
rect 107750 557832 107806 557841
rect 107750 557767 107806 557776
rect 107658 542872 107714 542881
rect 107658 542807 107714 542816
rect 107568 481704 107620 481710
rect 107568 481646 107620 481652
rect 107580 481574 107608 481646
rect 107568 481568 107620 481574
rect 107568 481510 107620 481516
rect 107476 469260 107528 469266
rect 107476 469202 107528 469208
rect 107566 467936 107622 467945
rect 107566 467871 107622 467880
rect 107580 465050 107608 467871
rect 107568 465044 107620 465050
rect 107568 464986 107620 464992
rect 107580 464370 107608 464986
rect 107568 464364 107620 464370
rect 107568 464306 107620 464312
rect 107384 449948 107436 449954
rect 107384 449890 107436 449896
rect 107672 449274 107700 542807
rect 107764 471510 107792 557767
rect 108316 556753 108344 571270
rect 108946 569256 109002 569265
rect 108946 569191 109002 569200
rect 108960 568614 108988 569191
rect 108948 568608 109000 568614
rect 108948 568550 109000 568556
rect 108856 568540 108908 568546
rect 108856 568482 108908 568488
rect 108868 567361 108896 568482
rect 108946 567896 109002 567905
rect 108946 567831 109002 567840
rect 108854 567352 108910 567361
rect 108854 567287 108910 567296
rect 108960 567254 108988 567831
rect 108948 567248 109000 567254
rect 108948 567190 109000 567196
rect 108946 566536 109002 566545
rect 108946 566471 108948 566480
rect 109000 566471 109002 566480
rect 108948 566442 109000 566448
rect 108948 565888 109000 565894
rect 108946 565856 108948 565865
rect 109000 565856 109002 565865
rect 108856 565820 108908 565826
rect 108946 565791 109002 565800
rect 108856 565762 108908 565768
rect 108868 565321 108896 565762
rect 108854 565312 108910 565321
rect 108854 565247 108910 565256
rect 108946 563816 109002 563825
rect 108946 563751 109002 563760
rect 108960 563514 108988 563751
rect 108948 563508 109000 563514
rect 108948 563450 109000 563456
rect 108946 563136 109002 563145
rect 108946 563071 109002 563080
rect 108854 562456 108910 562465
rect 108854 562391 108910 562400
rect 108868 560998 108896 562391
rect 108960 562358 108988 563071
rect 108948 562352 109000 562358
rect 108948 562294 109000 562300
rect 108946 561096 109002 561105
rect 108946 561031 108948 561040
rect 109000 561031 109002 561040
rect 108948 561002 109000 561008
rect 108856 560992 108908 560998
rect 108856 560934 108908 560940
rect 108946 560552 109002 560561
rect 109052 560538 109080 658378
rect 109408 647284 109460 647290
rect 109460 647232 109540 647234
rect 109408 647226 109540 647232
rect 109420 647206 109540 647226
rect 109314 645960 109370 645969
rect 109002 560510 109080 560538
rect 109144 645918 109314 645946
rect 108946 560487 109002 560496
rect 108946 559736 109002 559745
rect 108946 559671 109002 559680
rect 108960 559570 108988 559671
rect 108948 559564 109000 559570
rect 108948 559506 109000 559512
rect 108946 558376 109002 558385
rect 108946 558311 109002 558320
rect 108960 558210 108988 558311
rect 108948 558204 109000 558210
rect 108948 558146 109000 558152
rect 108948 557184 109000 557190
rect 108946 557152 108948 557161
rect 109000 557152 109002 557161
rect 108946 557087 109002 557096
rect 108302 556744 108358 556753
rect 108302 556679 108358 556688
rect 108854 555656 108910 555665
rect 108854 555591 108910 555600
rect 108868 554810 108896 555591
rect 108856 554804 108908 554810
rect 108856 554746 108908 554752
rect 108948 554736 109000 554742
rect 108948 554678 109000 554684
rect 108960 554441 108988 554678
rect 108946 554432 109002 554441
rect 108946 554367 109002 554376
rect 108948 554056 109000 554062
rect 108948 553998 109000 554004
rect 108960 553761 108988 553998
rect 108946 553752 109002 553761
rect 108946 553687 109002 553696
rect 108302 552936 108358 552945
rect 108302 552871 108358 552880
rect 108316 552022 108344 552871
rect 108946 552256 109002 552265
rect 108946 552191 109002 552200
rect 108960 552090 108988 552191
rect 108948 552084 109000 552090
rect 108948 552026 109000 552032
rect 108304 552016 108356 552022
rect 108304 551958 108356 551964
rect 108026 540016 108082 540025
rect 108026 539951 108082 539960
rect 108040 539646 108068 539951
rect 108028 539640 108080 539646
rect 108028 539582 108080 539588
rect 107752 471504 107804 471510
rect 107752 471446 107804 471452
rect 108316 463418 108344 551958
rect 108946 551576 109002 551585
rect 108946 551511 109002 551520
rect 108960 550662 108988 551511
rect 108948 550656 109000 550662
rect 108948 550598 109000 550604
rect 108854 550216 108910 550225
rect 108854 550151 108910 550160
rect 108868 548554 108896 550151
rect 109144 549953 109172 645918
rect 109314 645895 109370 645904
rect 109342 640070 109448 640098
rect 109420 637673 109448 640070
rect 109512 639849 109540 647206
rect 109590 640520 109646 640529
rect 109590 640455 109646 640464
rect 109498 639840 109554 639849
rect 109498 639775 109554 639784
rect 109406 637664 109462 637673
rect 109406 637599 109462 637608
rect 109604 625154 109632 640455
rect 109682 638888 109738 638897
rect 109682 638823 109738 638832
rect 109420 625126 109632 625154
rect 109130 549944 109186 549953
rect 109130 549879 109186 549888
rect 108948 549228 109000 549234
rect 108948 549170 109000 549176
rect 108960 549001 108988 549170
rect 108946 548992 109002 549001
rect 108946 548927 109002 548936
rect 108856 548548 108908 548554
rect 108856 548490 108908 548496
rect 108946 547496 109002 547505
rect 108946 547431 109002 547440
rect 108960 547194 108988 547431
rect 108948 547188 109000 547194
rect 108948 547130 109000 547136
rect 108762 546952 108818 546961
rect 108762 546887 108818 546896
rect 108776 538214 108804 546887
rect 108946 546136 109002 546145
rect 108946 546071 109002 546080
rect 108960 545698 108988 546071
rect 108948 545692 109000 545698
rect 108948 545634 109000 545640
rect 108854 545456 108910 545465
rect 108854 545391 108910 545400
rect 108868 544406 108896 545391
rect 108946 544776 109002 544785
rect 108946 544711 109002 544720
rect 108960 544474 108988 544711
rect 108948 544468 109000 544474
rect 108948 544410 109000 544416
rect 108856 544400 108908 544406
rect 108856 544342 108908 544348
rect 108854 544096 108910 544105
rect 108854 544031 108910 544040
rect 108868 543794 108896 544031
rect 109420 543794 109448 625126
rect 109696 573986 109724 638823
rect 110432 574530 110460 672551
rect 110510 665816 110566 665825
rect 110510 665751 110566 665760
rect 110420 574524 110472 574530
rect 110420 574466 110472 574472
rect 109684 573980 109736 573986
rect 109684 573922 109736 573928
rect 109696 573374 109724 573922
rect 109684 573368 109736 573374
rect 109684 573310 109736 573316
rect 110524 567254 110552 665751
rect 110616 658481 110644 697546
rect 111798 678736 111854 678745
rect 111798 678671 111854 678680
rect 111812 677686 111840 678671
rect 112350 678056 112406 678065
rect 112350 677991 112406 678000
rect 111800 677680 111852 677686
rect 111800 677622 111852 677628
rect 112364 677618 112392 677991
rect 112352 677612 112404 677618
rect 112352 677554 112404 677560
rect 111798 677376 111854 677385
rect 111798 677311 111854 677320
rect 111812 676326 111840 677311
rect 112718 676696 112774 676705
rect 112718 676631 112774 676640
rect 111800 676320 111852 676326
rect 111800 676262 111852 676268
rect 112732 676258 112760 676631
rect 113100 676297 113128 702510
rect 113180 681012 113232 681018
rect 113180 680954 113232 680960
rect 113086 676288 113142 676297
rect 112720 676252 112772 676258
rect 113086 676223 113142 676232
rect 112720 676194 112772 676200
rect 111982 676016 112038 676025
rect 111982 675951 112038 675960
rect 111996 674898 112024 675951
rect 113100 675481 113128 676223
rect 113086 675472 113142 675481
rect 113086 675407 113142 675416
rect 111984 674892 112036 674898
rect 111984 674834 112036 674840
rect 112074 674656 112130 674665
rect 112074 674591 112130 674600
rect 111800 672036 111852 672042
rect 111800 671978 111852 671984
rect 111812 671809 111840 671978
rect 111798 671800 111854 671809
rect 111798 671735 111854 671744
rect 111798 671256 111854 671265
rect 111798 671191 111854 671200
rect 111812 670750 111840 671191
rect 111800 670744 111852 670750
rect 111800 670686 111852 670692
rect 111798 670576 111854 670585
rect 111798 670511 111854 670520
rect 111812 669526 111840 670511
rect 111800 669520 111852 669526
rect 111800 669462 111852 669468
rect 111800 669384 111852 669390
rect 111798 669352 111800 669361
rect 111852 669352 111854 669361
rect 111798 669287 111854 669296
rect 111982 667176 112038 667185
rect 111982 667111 112038 667120
rect 111798 666632 111854 666641
rect 111798 666567 111800 666576
rect 111852 666567 111854 666576
rect 111800 666538 111852 666544
rect 111798 665272 111854 665281
rect 111798 665207 111800 665216
rect 111852 665207 111854 665216
rect 111800 665178 111852 665184
rect 111798 663912 111854 663921
rect 111798 663847 111854 663856
rect 111812 663814 111840 663847
rect 111800 663808 111852 663814
rect 111800 663750 111852 663756
rect 111798 662552 111854 662561
rect 111798 662487 111854 662496
rect 111812 662454 111840 662487
rect 111800 662448 111852 662454
rect 111800 662390 111852 662396
rect 111156 661564 111208 661570
rect 111156 661506 111208 661512
rect 111168 661201 111196 661506
rect 111154 661192 111210 661201
rect 111154 661127 111210 661136
rect 110602 658472 110658 658481
rect 110602 658407 110604 658416
rect 110656 658407 110658 658416
rect 110604 658378 110656 658384
rect 110616 658347 110644 658378
rect 110602 654256 110658 654265
rect 110602 654191 110658 654200
rect 110512 567248 110564 567254
rect 110512 567190 110564 567196
rect 110616 557190 110644 654191
rect 111168 640334 111196 661127
rect 111798 659016 111854 659025
rect 111798 658951 111854 658960
rect 111076 640306 111196 640334
rect 111076 563514 111104 640306
rect 111708 564188 111760 564194
rect 111708 564130 111760 564136
rect 111156 563848 111208 563854
rect 111156 563790 111208 563796
rect 111064 563508 111116 563514
rect 111064 563450 111116 563456
rect 110604 557184 110656 557190
rect 110604 557126 110656 557132
rect 110616 556850 110644 557126
rect 110604 556844 110656 556850
rect 110604 556786 110656 556792
rect 109776 555416 109828 555422
rect 109776 555358 109828 555364
rect 109684 551336 109736 551342
rect 109684 551278 109736 551284
rect 108856 543788 108908 543794
rect 108856 543730 108908 543736
rect 109408 543788 109460 543794
rect 109408 543730 109460 543736
rect 108948 543720 109000 543726
rect 108948 543662 109000 543668
rect 108960 543561 108988 543662
rect 108946 543552 109002 543561
rect 108946 543487 109002 543496
rect 108854 542056 108910 542065
rect 108854 541991 108910 542000
rect 108868 541006 108896 541991
rect 108856 541000 108908 541006
rect 108856 540942 108908 540948
rect 108948 540932 109000 540938
rect 108948 540874 109000 540880
rect 108960 540841 108988 540874
rect 108946 540832 109002 540841
rect 108946 540767 109002 540776
rect 108776 538186 108988 538214
rect 108394 469296 108450 469305
rect 108394 469231 108450 469240
rect 108304 463412 108356 463418
rect 108304 463354 108356 463360
rect 108304 458924 108356 458930
rect 108304 458866 108356 458872
rect 108316 457570 108344 458866
rect 108304 457564 108356 457570
rect 108304 457506 108356 457512
rect 107660 449268 107712 449274
rect 107660 449210 107712 449216
rect 107476 448656 107528 448662
rect 107476 448598 107528 448604
rect 107488 396914 107516 448598
rect 108408 437374 108436 469231
rect 108960 456822 108988 538186
rect 109040 530732 109092 530738
rect 109040 530674 109092 530680
rect 109052 481545 109080 530674
rect 109130 491328 109186 491337
rect 109130 491263 109186 491272
rect 109144 491230 109172 491263
rect 109696 491230 109724 551278
rect 109788 537878 109816 555358
rect 111064 550588 111116 550594
rect 111064 550530 111116 550536
rect 109868 549160 109920 549166
rect 109868 549102 109920 549108
rect 109776 537872 109828 537878
rect 109776 537814 109828 537820
rect 109776 491496 109828 491502
rect 109776 491438 109828 491444
rect 109132 491224 109184 491230
rect 109132 491166 109184 491172
rect 109684 491224 109736 491230
rect 109684 491166 109736 491172
rect 109682 489968 109738 489977
rect 109682 489903 109738 489912
rect 109038 481536 109094 481545
rect 109038 481471 109094 481480
rect 108488 456816 108540 456822
rect 108488 456758 108540 456764
rect 108948 456816 109000 456822
rect 108948 456758 109000 456764
rect 108500 455394 108528 456758
rect 108488 455388 108540 455394
rect 108488 455330 108540 455336
rect 108948 454980 109000 454986
rect 108948 454922 109000 454928
rect 108854 452568 108910 452577
rect 108854 452503 108910 452512
rect 108764 442264 108816 442270
rect 108764 442206 108816 442212
rect 108396 437368 108448 437374
rect 108396 437310 108448 437316
rect 107476 396908 107528 396914
rect 107476 396850 107528 396856
rect 108304 396704 108356 396710
rect 108304 396646 108356 396652
rect 107660 394052 107712 394058
rect 107660 393994 107712 394000
rect 107212 393286 107332 393314
rect 107212 386510 107240 393286
rect 107672 387802 107700 393994
rect 108316 387938 108344 396646
rect 108776 394058 108804 442206
rect 108868 399498 108896 452503
rect 108856 399492 108908 399498
rect 108856 399434 108908 399440
rect 108960 395321 108988 454922
rect 108946 395312 109002 395321
rect 108946 395247 109002 395256
rect 108764 394052 108816 394058
rect 108764 393994 108816 394000
rect 109696 387977 109724 489903
rect 109788 390182 109816 491438
rect 109880 491434 109908 549102
rect 110420 541000 110472 541006
rect 110420 540942 110472 540948
rect 110432 540870 110460 540942
rect 110420 540864 110472 540870
rect 110420 540806 110472 540812
rect 111076 528630 111104 550530
rect 111168 549166 111196 563790
rect 111248 563712 111300 563718
rect 111248 563654 111300 563660
rect 111156 549160 111208 549166
rect 111156 549102 111208 549108
rect 111156 540864 111208 540870
rect 111156 540806 111208 540812
rect 111064 528624 111116 528630
rect 111064 528566 111116 528572
rect 110420 493944 110472 493950
rect 110420 493886 110472 493892
rect 110432 493406 110460 493886
rect 110420 493400 110472 493406
rect 110420 493342 110472 493348
rect 110420 492788 110472 492794
rect 110420 492730 110472 492736
rect 109868 491428 109920 491434
rect 109868 491370 109920 491376
rect 109880 398818 109908 491370
rect 109868 398812 109920 398818
rect 109868 398754 109920 398760
rect 110328 391264 110380 391270
rect 110328 391206 110380 391212
rect 109776 390176 109828 390182
rect 109776 390118 109828 390124
rect 109682 387968 109738 387977
rect 108304 387932 108356 387938
rect 109682 387903 109738 387912
rect 108304 387874 108356 387880
rect 107660 387796 107712 387802
rect 107660 387738 107712 387744
rect 107200 386504 107252 386510
rect 107200 386446 107252 386452
rect 106292 385886 106766 385914
rect 107212 385778 107240 386446
rect 108316 386034 108344 387874
rect 108488 387796 108540 387802
rect 108488 387738 108540 387744
rect 108500 386646 108528 387738
rect 108488 386640 108540 386646
rect 108488 386582 108540 386588
rect 108304 386028 108356 386034
rect 108304 385970 108356 385976
rect 108500 385778 108528 386582
rect 109696 385914 109724 387903
rect 110340 385914 110368 391206
rect 110432 389162 110460 492730
rect 110512 491360 110564 491366
rect 110512 491302 110564 491308
rect 110524 491201 110552 491302
rect 110510 491192 110566 491201
rect 110510 491127 110566 491136
rect 110604 482792 110656 482798
rect 110604 482734 110656 482740
rect 110512 394120 110564 394126
rect 110512 394062 110564 394068
rect 110420 389156 110472 389162
rect 110420 389098 110472 389104
rect 110432 388482 110460 389098
rect 110420 388476 110472 388482
rect 110420 388418 110472 388424
rect 110524 386050 110552 394062
rect 110616 387122 110644 482734
rect 111076 459678 111104 528566
rect 111168 478922 111196 540806
rect 111260 538898 111288 563654
rect 111248 538892 111300 538898
rect 111248 538834 111300 538840
rect 111720 493950 111748 564130
rect 111812 561066 111840 658951
rect 111890 654936 111946 654945
rect 111890 654871 111946 654880
rect 111800 561060 111852 561066
rect 111800 561002 111852 561008
rect 111904 558822 111932 654871
rect 111996 650978 112024 667111
rect 112088 654134 112116 674591
rect 112718 669896 112774 669905
rect 112718 669831 112774 669840
rect 112732 669458 112760 669831
rect 112720 669452 112772 669458
rect 112720 669394 112772 669400
rect 112350 664456 112406 664465
rect 112350 664391 112406 664400
rect 112364 663882 112392 664391
rect 112352 663876 112404 663882
rect 112352 663818 112404 663824
rect 112350 660376 112406 660385
rect 112350 660311 112406 660320
rect 112364 659734 112392 660311
rect 112534 659832 112590 659841
rect 112534 659767 112536 659776
rect 112588 659767 112590 659776
rect 112536 659738 112588 659744
rect 112352 659728 112404 659734
rect 112352 659670 112404 659676
rect 112534 656976 112590 656985
rect 112534 656911 112536 656920
rect 112588 656911 112590 656920
rect 112536 656882 112588 656888
rect 112350 656296 112406 656305
rect 112350 656231 112406 656240
rect 112364 655586 112392 656231
rect 112536 655648 112588 655654
rect 112534 655616 112536 655625
rect 112588 655616 112590 655625
rect 112352 655580 112404 655586
rect 112534 655551 112590 655560
rect 112352 655522 112404 655528
rect 112088 654106 112300 654134
rect 111996 650950 112208 650978
rect 112074 650856 112130 650865
rect 112074 650791 112130 650800
rect 111982 650176 112038 650185
rect 112088 650146 112116 650791
rect 111982 650111 112038 650120
rect 112076 650140 112128 650146
rect 111996 650078 112024 650111
rect 112076 650082 112128 650088
rect 111984 650072 112036 650078
rect 111984 650014 112036 650020
rect 111982 648136 112038 648145
rect 111982 648071 112038 648080
rect 111892 558816 111944 558822
rect 111892 558758 111944 558764
rect 111996 551274 112024 648071
rect 112180 647290 112208 650950
rect 112168 647284 112220 647290
rect 112168 647226 112220 647232
rect 112272 639674 112300 654106
rect 113086 652896 113142 652905
rect 113192 652882 113220 680954
rect 113836 661570 113864 702714
rect 114560 670744 114612 670750
rect 114560 670686 114612 670692
rect 113824 661564 113876 661570
rect 113824 661506 113876 661512
rect 113142 652854 113312 652882
rect 113086 652831 113142 652840
rect 112534 651536 112590 651545
rect 112534 651471 112590 651480
rect 112548 651438 112576 651471
rect 112536 651432 112588 651438
rect 112536 651374 112588 651380
rect 113086 649496 113142 649505
rect 113086 649431 113142 649440
rect 112994 648816 113050 648825
rect 112994 648751 113050 648760
rect 113008 648718 113036 648751
rect 112996 648712 113048 648718
rect 112996 648654 113048 648660
rect 113100 648650 113128 649431
rect 113088 648644 113140 648650
rect 113088 648586 113140 648592
rect 113086 647456 113142 647465
rect 113086 647391 113142 647400
rect 113100 647290 113128 647391
rect 113088 647284 113140 647290
rect 113088 647226 113140 647232
rect 112994 645416 113050 645425
rect 112994 645351 113050 645360
rect 113008 644570 113036 645351
rect 113086 644736 113142 644745
rect 113086 644671 113142 644680
rect 112996 644564 113048 644570
rect 112996 644506 113048 644512
rect 113100 644502 113128 644671
rect 113088 644496 113140 644502
rect 113088 644438 113140 644444
rect 112812 644360 112864 644366
rect 112812 644302 112864 644308
rect 112824 643521 112852 644302
rect 112810 643512 112866 643521
rect 112810 643447 112866 643456
rect 113086 642696 113142 642705
rect 113086 642631 113142 642640
rect 112626 642152 112682 642161
rect 112626 642087 112628 642096
rect 112680 642087 112682 642096
rect 112628 642058 112680 642064
rect 113100 641782 113128 642631
rect 113088 641776 113140 641782
rect 113088 641718 113140 641724
rect 112902 639976 112958 639985
rect 112902 639911 112958 639920
rect 112260 639668 112312 639674
rect 112260 639610 112312 639616
rect 112916 638994 112944 639911
rect 112904 638988 112956 638994
rect 112904 638930 112956 638936
rect 113178 638616 113234 638625
rect 113178 638551 113234 638560
rect 112904 559632 112956 559638
rect 112904 559574 112956 559580
rect 112628 551404 112680 551410
rect 112628 551346 112680 551352
rect 111984 551268 112036 551274
rect 111984 551210 112036 551216
rect 112260 536784 112312 536790
rect 112260 536726 112312 536732
rect 112272 536382 112300 536726
rect 112260 536376 112312 536382
rect 112260 536318 112312 536324
rect 111800 494080 111852 494086
rect 111800 494022 111852 494028
rect 111708 493944 111760 493950
rect 111708 493886 111760 493892
rect 111156 478916 111208 478922
rect 111156 478858 111208 478864
rect 111064 459672 111116 459678
rect 111064 459614 111116 459620
rect 111076 459542 111104 459614
rect 111064 459536 111116 459542
rect 111064 459478 111116 459484
rect 111812 454986 111840 494022
rect 112536 491224 112588 491230
rect 112536 491166 112588 491172
rect 112444 489184 112496 489190
rect 112444 489126 112496 489132
rect 111892 477556 111944 477562
rect 111892 477498 111944 477504
rect 111904 477358 111932 477498
rect 111892 477352 111944 477358
rect 111892 477294 111944 477300
rect 111800 454980 111852 454986
rect 111800 454922 111852 454928
rect 110604 387116 110656 387122
rect 110604 387058 110656 387064
rect 112456 386578 112484 489126
rect 112548 388686 112576 491166
rect 112640 489258 112668 551346
rect 112916 536382 112944 559574
rect 112996 555552 113048 555558
rect 112996 555494 113048 555500
rect 112904 536376 112956 536382
rect 112904 536318 112956 536324
rect 113008 492114 113036 555494
rect 113088 555484 113140 555490
rect 113088 555426 113140 555432
rect 112996 492108 113048 492114
rect 112996 492050 113048 492056
rect 112628 489252 112680 489258
rect 112628 489194 112680 489200
rect 113100 477562 113128 555426
rect 113192 539646 113220 638551
rect 113284 554810 113312 652854
rect 113456 585200 113508 585206
rect 113456 585142 113508 585148
rect 113364 582480 113416 582486
rect 113364 582422 113416 582428
rect 113376 564194 113404 582422
rect 113468 568585 113496 585142
rect 114572 573238 114600 670686
rect 115216 638625 115244 703054
rect 116584 702908 116636 702914
rect 116584 702850 116636 702856
rect 115296 702704 115348 702710
rect 115296 702646 115348 702652
rect 115308 644473 115336 702646
rect 115940 648712 115992 648718
rect 115940 648654 115992 648660
rect 115294 644464 115350 644473
rect 115294 644399 115350 644408
rect 115308 644366 115336 644399
rect 115296 644360 115348 644366
rect 115296 644302 115348 644308
rect 115202 638616 115258 638625
rect 115202 638551 115258 638560
rect 115848 618248 115900 618254
rect 115848 618190 115900 618196
rect 114652 583908 114704 583914
rect 114652 583850 114704 583856
rect 114560 573232 114612 573238
rect 114560 573174 114612 573180
rect 113454 568576 113510 568585
rect 113454 568511 113510 568520
rect 113548 567248 113600 567254
rect 113548 567190 113600 567196
rect 113364 564188 113416 564194
rect 113364 564130 113416 564136
rect 113560 555490 113588 567190
rect 113824 563508 113876 563514
rect 113824 563450 113876 563456
rect 113548 555484 113600 555490
rect 113548 555426 113600 555432
rect 113272 554804 113324 554810
rect 113272 554746 113324 554752
rect 113272 543788 113324 543794
rect 113272 543730 113324 543736
rect 113180 539640 113232 539646
rect 113180 539582 113232 539588
rect 113180 536376 113232 536382
rect 113180 536318 113232 536324
rect 113088 477556 113140 477562
rect 113088 477498 113140 477504
rect 112628 445868 112680 445874
rect 112628 445810 112680 445816
rect 112640 392601 112668 445810
rect 113192 442513 113220 536318
rect 113284 448662 113312 543730
rect 113836 472054 113864 563450
rect 114100 554804 114152 554810
rect 114100 554746 114152 554752
rect 114112 553450 114140 554746
rect 114100 553444 114152 553450
rect 114100 553386 114152 553392
rect 114572 539578 114600 573174
rect 114560 539572 114612 539578
rect 114560 539514 114612 539520
rect 114560 495576 114612 495582
rect 114560 495518 114612 495524
rect 113916 493944 113968 493950
rect 113916 493886 113968 493892
rect 113824 472048 113876 472054
rect 113824 471990 113876 471996
rect 113928 467158 113956 493886
rect 114466 493368 114522 493377
rect 114466 493303 114522 493312
rect 114480 492726 114508 493303
rect 114468 492720 114520 492726
rect 114468 492662 114520 492668
rect 114468 485172 114520 485178
rect 114468 485114 114520 485120
rect 114480 485081 114508 485114
rect 114466 485072 114522 485081
rect 114466 485007 114522 485016
rect 113916 467152 113968 467158
rect 113916 467094 113968 467100
rect 113272 448656 113324 448662
rect 113272 448598 113324 448604
rect 113178 442504 113234 442513
rect 113178 442439 113234 442448
rect 114100 398812 114152 398818
rect 114100 398754 114152 398760
rect 112626 392592 112682 392601
rect 112626 392527 112682 392536
rect 113914 390824 113970 390833
rect 113914 390759 113970 390768
rect 112536 388680 112588 388686
rect 112536 388622 112588 388628
rect 112548 387682 112576 388622
rect 112548 387654 112668 387682
rect 112168 386572 112220 386578
rect 112168 386514 112220 386520
rect 112444 386572 112496 386578
rect 112444 386514 112496 386520
rect 110524 386022 110920 386050
rect 109342 385886 109724 385914
rect 109986 385886 110368 385914
rect 110892 385914 110920 386022
rect 112180 385914 112208 386514
rect 112640 385914 112668 387654
rect 113928 385914 113956 390759
rect 114112 390726 114140 398754
rect 114572 396710 114600 495518
rect 114664 494834 114692 583850
rect 114744 581052 114796 581058
rect 114744 580994 114796 581000
rect 114756 563854 114784 580994
rect 114744 563848 114796 563854
rect 114744 563790 114796 563796
rect 115204 545692 115256 545698
rect 115204 545634 115256 545640
rect 115216 545193 115244 545634
rect 115202 545184 115258 545193
rect 115202 545119 115258 545128
rect 115204 539572 115256 539578
rect 115204 539514 115256 539520
rect 114744 534812 114796 534818
rect 114744 534754 114796 534760
rect 114652 494828 114704 494834
rect 114652 494770 114704 494776
rect 114652 492856 114704 492862
rect 114652 492798 114704 492804
rect 114664 406434 114692 492798
rect 114756 465798 114784 534754
rect 115216 481642 115244 539514
rect 115860 536858 115888 618190
rect 115952 550594 115980 648654
rect 116596 643074 116624 702850
rect 129004 700392 129056 700398
rect 129004 700334 129056 700340
rect 129016 687954 129044 700334
rect 136652 692102 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 700398 154160 703520
rect 170324 702434 170352 703520
rect 202800 703322 202828 703520
rect 201500 703316 201552 703322
rect 201500 703258 201552 703264
rect 202788 703316 202840 703322
rect 202788 703258 202840 703264
rect 169772 702406 170352 702434
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 136640 692096 136692 692102
rect 136640 692038 136692 692044
rect 169772 690674 169800 702406
rect 188344 700392 188396 700398
rect 188344 700334 188396 700340
rect 169760 690668 169812 690674
rect 169760 690610 169812 690616
rect 129004 687948 129056 687954
rect 129004 687890 129056 687896
rect 188356 683806 188384 700334
rect 188344 683800 188396 683806
rect 188344 683742 188396 683748
rect 196624 683188 196676 683194
rect 196624 683130 196676 683136
rect 125692 681760 125744 681766
rect 125692 681702 125744 681708
rect 118700 677680 118752 677686
rect 118700 677622 118752 677628
rect 117412 662448 117464 662454
rect 117412 662390 117464 662396
rect 116032 643068 116084 643074
rect 116032 643010 116084 643016
rect 116584 643068 116636 643074
rect 116584 643010 116636 643016
rect 116044 642122 116072 643010
rect 116032 642116 116084 642122
rect 116032 642058 116084 642064
rect 115940 550588 115992 550594
rect 115940 550530 115992 550536
rect 116044 544474 116072 642058
rect 117320 638444 117372 638450
rect 117320 638386 117372 638392
rect 116122 587344 116178 587353
rect 116122 587279 116178 587288
rect 116136 551410 116164 587279
rect 116214 583944 116270 583953
rect 116214 583879 116270 583888
rect 116228 563718 116256 583879
rect 116398 578232 116454 578241
rect 116398 578167 116454 578176
rect 116412 577522 116440 578167
rect 116400 577516 116452 577522
rect 116400 577458 116452 577464
rect 116308 576224 116360 576230
rect 116306 576192 116308 576201
rect 116360 576192 116362 576201
rect 116306 576127 116362 576136
rect 117134 576192 117190 576201
rect 117134 576127 117190 576136
rect 117148 575550 117176 576127
rect 117136 575544 117188 575550
rect 117136 575486 117188 575492
rect 116216 563712 116268 563718
rect 116216 563654 116268 563660
rect 116584 553444 116636 553450
rect 116584 553386 116636 553392
rect 116124 551404 116176 551410
rect 116124 551346 116176 551352
rect 116032 544468 116084 544474
rect 116032 544410 116084 544416
rect 115848 536852 115900 536858
rect 115848 536794 115900 536800
rect 115940 492040 115992 492046
rect 115940 491982 115992 491988
rect 115848 481772 115900 481778
rect 115848 481714 115900 481720
rect 115860 481642 115888 481714
rect 115204 481636 115256 481642
rect 115204 481578 115256 481584
rect 115848 481636 115900 481642
rect 115848 481578 115900 481584
rect 115296 478984 115348 478990
rect 115296 478926 115348 478932
rect 114744 465792 114796 465798
rect 114744 465734 114796 465740
rect 114652 406428 114704 406434
rect 114652 406370 114704 406376
rect 114560 396704 114612 396710
rect 114560 396646 114612 396652
rect 114100 390720 114152 390726
rect 114100 390662 114152 390668
rect 110892 385886 111274 385914
rect 111918 385886 112208 385914
rect 112562 385886 112668 385914
rect 113850 385886 113956 385914
rect 114112 385914 114140 390662
rect 114928 390176 114980 390182
rect 114928 390118 114980 390124
rect 114468 389972 114520 389978
rect 114468 389914 114520 389920
rect 114480 388618 114508 389914
rect 114468 388612 114520 388618
rect 114468 388554 114520 388560
rect 114940 387938 114968 390118
rect 115204 390108 115256 390114
rect 115204 390050 115256 390056
rect 114928 387932 114980 387938
rect 114928 387874 114980 387880
rect 114112 385886 114494 385914
rect 114940 385778 114968 387874
rect 104636 385750 104834 385778
rect 107212 385750 107410 385778
rect 108500 385750 108698 385778
rect 114940 385750 115138 385778
rect 95424 385688 95476 385694
rect 95424 385630 95476 385636
rect 71792 385354 71990 385370
rect 92952 385354 93348 385370
rect 71780 385348 71990 385354
rect 71832 385342 71990 385348
rect 92940 385348 93348 385354
rect 71780 385290 71832 385296
rect 92992 385342 93348 385348
rect 104190 385354 104480 385370
rect 104190 385348 104492 385354
rect 104190 385342 104440 385348
rect 92940 385290 92992 385296
rect 104440 385290 104492 385296
rect 115216 373994 115244 390050
rect 115308 374649 115336 478926
rect 115848 406428 115900 406434
rect 115848 406370 115900 406376
rect 115860 406337 115888 406370
rect 115846 406328 115902 406337
rect 115846 406263 115902 406272
rect 115848 394800 115900 394806
rect 115848 394742 115900 394748
rect 115860 394670 115888 394742
rect 115848 394664 115900 394670
rect 115848 394606 115900 394612
rect 115848 389904 115900 389910
rect 115848 389846 115900 389852
rect 115860 385914 115888 389846
rect 115952 388550 115980 491982
rect 116044 451926 116072 544410
rect 116596 463690 116624 553386
rect 117332 536586 117360 638386
rect 117424 565826 117452 662390
rect 117594 587480 117650 587489
rect 117594 587415 117650 587424
rect 117412 565820 117464 565826
rect 117412 565762 117464 565768
rect 117424 564466 117452 565762
rect 117412 564460 117464 564466
rect 117412 564402 117464 564408
rect 117504 561060 117556 561066
rect 117504 561002 117556 561008
rect 117320 536580 117372 536586
rect 117320 536522 117372 536528
rect 117332 535498 117360 536522
rect 117320 535492 117372 535498
rect 117320 535434 117372 535440
rect 117228 488572 117280 488578
rect 117228 488514 117280 488520
rect 117240 488481 117268 488514
rect 117226 488472 117282 488481
rect 117148 488430 117226 488458
rect 117148 480254 117176 488430
rect 117226 488407 117282 488416
rect 117226 485752 117282 485761
rect 117226 485687 117282 485696
rect 117240 485110 117268 485687
rect 117228 485104 117280 485110
rect 117228 485046 117280 485052
rect 117410 485072 117466 485081
rect 117240 484430 117268 485046
rect 117410 485007 117466 485016
rect 117228 484424 117280 484430
rect 117228 484366 117280 484372
rect 117148 480226 117268 480254
rect 117240 463690 117268 480226
rect 116584 463684 116636 463690
rect 116584 463626 116636 463632
rect 117228 463684 117280 463690
rect 117228 463626 117280 463632
rect 116032 451920 116084 451926
rect 116032 451862 116084 451868
rect 116044 451586 116072 451862
rect 116032 451580 116084 451586
rect 116032 451522 116084 451528
rect 116584 451580 116636 451586
rect 116584 451522 116636 451528
rect 115940 388544 115992 388550
rect 115940 388486 115992 388492
rect 115940 387116 115992 387122
rect 115940 387058 115992 387064
rect 115782 385886 115888 385914
rect 115952 378593 115980 387058
rect 116400 381540 116452 381546
rect 116400 381482 116452 381488
rect 116412 380905 116440 381482
rect 116398 380896 116454 380905
rect 116398 380831 116454 380840
rect 115938 378584 115994 378593
rect 115938 378519 115994 378528
rect 115478 377496 115534 377505
rect 115478 377431 115534 377440
rect 115294 374640 115350 374649
rect 115294 374575 115350 374584
rect 115216 373966 115336 373994
rect 115308 371929 115336 373966
rect 115492 373153 115520 377431
rect 115478 373144 115534 373153
rect 115478 373079 115534 373088
rect 115848 371952 115900 371958
rect 115294 371920 115350 371929
rect 115848 371894 115900 371900
rect 115294 371855 115350 371864
rect 69664 369164 69716 369170
rect 69664 369106 69716 369112
rect 115294 367024 115350 367033
rect 115294 366959 115350 366968
rect 69662 349888 69718 349897
rect 69662 349823 69718 349832
rect 69676 349110 69704 349823
rect 69664 349104 69716 349110
rect 69664 349046 69716 349052
rect 69296 340740 69348 340746
rect 69296 340682 69348 340688
rect 69676 334694 69704 349046
rect 69756 340740 69808 340746
rect 69756 340682 69808 340688
rect 69768 340082 69796 340682
rect 70400 340264 70452 340270
rect 70400 340206 70452 340212
rect 69768 340068 70058 340082
rect 69768 340054 70072 340068
rect 70044 337142 70072 340054
rect 70032 337136 70084 337142
rect 70032 337078 70084 337084
rect 70412 336530 70440 340206
rect 70504 340054 70702 340082
rect 70504 337890 70532 340054
rect 70492 337884 70544 337890
rect 70492 337826 70544 337832
rect 70400 336524 70452 336530
rect 70400 336466 70452 336472
rect 69664 334688 69716 334694
rect 69664 334630 69716 334636
rect 69112 330744 69164 330750
rect 69112 330686 69164 330692
rect 70400 326392 70452 326398
rect 70400 326334 70452 326340
rect 68836 307828 68888 307834
rect 68836 307770 68888 307776
rect 68744 305720 68796 305726
rect 68744 305662 68796 305668
rect 68652 299464 68704 299470
rect 68652 299406 68704 299412
rect 68664 298314 68692 299406
rect 68652 298308 68704 298314
rect 68652 298250 68704 298256
rect 67640 291168 67692 291174
rect 67640 291110 67692 291116
rect 67652 290873 67680 291110
rect 67638 290864 67694 290873
rect 67638 290799 67694 290808
rect 67638 290184 67694 290193
rect 67638 290119 67694 290128
rect 67652 289882 67680 290119
rect 67640 289876 67692 289882
rect 67640 289818 67692 289824
rect 67638 288824 67694 288833
rect 67638 288759 67694 288768
rect 67652 288454 67680 288759
rect 67640 288448 67692 288454
rect 67640 288390 67692 288396
rect 68664 288153 68692 298250
rect 68744 292664 68796 292670
rect 68744 292606 68796 292612
rect 68650 288144 68706 288153
rect 68650 288079 68706 288088
rect 67638 287464 67694 287473
rect 67638 287399 67694 287408
rect 67652 287094 67680 287399
rect 67640 287088 67692 287094
rect 67640 287030 67692 287036
rect 67822 287056 67878 287065
rect 67732 287020 67784 287026
rect 67822 286991 67878 287000
rect 67732 286962 67784 286968
rect 67640 286952 67692 286958
rect 67640 286894 67692 286900
rect 67652 286113 67680 286894
rect 67744 286793 67772 286962
rect 67730 286784 67786 286793
rect 67730 286719 67786 286728
rect 67638 286104 67694 286113
rect 67638 286039 67694 286048
rect 67836 285734 67864 286991
rect 67824 285728 67876 285734
rect 67824 285670 67876 285676
rect 67640 285660 67692 285666
rect 67640 285602 67692 285608
rect 67652 285433 67680 285602
rect 67638 285424 67694 285433
rect 67638 285359 67694 285368
rect 67638 284472 67694 284481
rect 67638 284407 67694 284416
rect 67652 284374 67680 284407
rect 67640 284368 67692 284374
rect 67640 284310 67692 284316
rect 67640 282872 67692 282878
rect 67640 282814 67692 282820
rect 67652 282169 67680 282814
rect 67638 282160 67694 282169
rect 67638 282095 67694 282104
rect 67638 280392 67694 280401
rect 67638 280327 67694 280336
rect 67652 280226 67680 280327
rect 67640 280220 67692 280226
rect 67640 280162 67692 280168
rect 67732 280152 67784 280158
rect 67732 280094 67784 280100
rect 67744 279857 67772 280094
rect 67730 279848 67786 279857
rect 67730 279783 67786 279792
rect 67640 279472 67692 279478
rect 67640 279414 67692 279420
rect 67652 279313 67680 279414
rect 67638 279304 67694 279313
rect 67638 279239 67694 279248
rect 67638 277672 67694 277681
rect 67638 277607 67694 277616
rect 67652 277438 67680 277607
rect 67640 277432 67692 277438
rect 67640 277374 67692 277380
rect 67822 276992 67878 277001
rect 67822 276927 67878 276936
rect 67640 276684 67692 276690
rect 67640 276626 67692 276632
rect 67652 275913 67680 276626
rect 67638 275904 67694 275913
rect 67638 275839 67694 275848
rect 67638 274952 67694 274961
rect 67638 274887 67694 274896
rect 67652 274718 67680 274887
rect 67640 274712 67692 274718
rect 67640 274654 67692 274660
rect 67732 274644 67784 274650
rect 67732 274586 67784 274592
rect 67744 274553 67772 274586
rect 67730 274544 67786 274553
rect 67730 274479 67786 274488
rect 67638 273592 67694 273601
rect 67638 273527 67694 273536
rect 67652 273290 67680 273527
rect 67640 273284 67692 273290
rect 67640 273226 67692 273232
rect 67732 271856 67784 271862
rect 67732 271798 67784 271804
rect 67638 271008 67694 271017
rect 67638 270943 67694 270952
rect 67652 270570 67680 270943
rect 67744 270881 67772 271798
rect 67730 270872 67786 270881
rect 67730 270807 67786 270816
rect 67640 270564 67692 270570
rect 67640 270506 67692 270512
rect 67732 270496 67784 270502
rect 67732 270438 67784 270444
rect 67744 269793 67772 270438
rect 67836 269822 67864 276927
rect 68756 276593 68784 292606
rect 68848 278633 68876 307770
rect 69020 299532 69072 299538
rect 69020 299474 69072 299480
rect 69032 298353 69060 299474
rect 69018 298344 69074 298353
rect 69018 298279 69074 298288
rect 69112 298172 69164 298178
rect 69112 298114 69164 298120
rect 68928 295588 68980 295594
rect 68928 295530 68980 295536
rect 68834 278624 68890 278633
rect 68834 278559 68890 278568
rect 68742 276584 68798 276593
rect 68742 276519 68798 276528
rect 68742 272232 68798 272241
rect 68742 272167 68798 272176
rect 68190 270192 68246 270201
rect 68190 270127 68246 270136
rect 67824 269816 67876 269822
rect 67730 269784 67786 269793
rect 67824 269758 67876 269764
rect 67730 269719 67786 269728
rect 68204 269142 68232 270127
rect 68192 269136 68244 269142
rect 68192 269078 68244 269084
rect 67640 269068 67692 269074
rect 67640 269010 67692 269016
rect 67652 268433 67680 269010
rect 68558 268832 68614 268841
rect 68558 268767 68614 268776
rect 67638 268424 67694 268433
rect 67638 268359 67694 268368
rect 67732 267708 67784 267714
rect 67732 267650 67784 267656
rect 67638 267064 67694 267073
rect 67638 266999 67640 267008
rect 67692 266999 67694 267008
rect 67640 266970 67692 266976
rect 67744 266937 67772 267650
rect 67730 266928 67786 266937
rect 67730 266863 67786 266872
rect 67732 266348 67784 266354
rect 67732 266290 67784 266296
rect 67638 265432 67694 265441
rect 67638 265367 67694 265376
rect 67652 264994 67680 265367
rect 67744 265033 67772 266290
rect 67730 265024 67786 265033
rect 67640 264988 67692 264994
rect 68572 264994 68600 268767
rect 67730 264959 67786 264968
rect 68560 264988 68612 264994
rect 67640 264930 67692 264936
rect 68560 264930 68612 264936
rect 67730 264208 67786 264217
rect 67730 264143 67786 264152
rect 67640 263696 67692 263702
rect 67638 263664 67640 263673
rect 67692 263664 67694 263673
rect 67744 263634 67772 264143
rect 67638 263599 67694 263608
rect 67732 263628 67784 263634
rect 67732 263570 67784 263576
rect 67640 263560 67692 263566
rect 67638 263528 67640 263537
rect 67692 263528 67694 263537
rect 67638 263463 67694 263472
rect 68560 262948 68612 262954
rect 68560 262890 68612 262896
rect 67638 262304 67694 262313
rect 67638 262239 67640 262248
rect 67692 262239 67694 262248
rect 67640 262210 67692 262216
rect 67732 262200 67784 262206
rect 67730 262168 67732 262177
rect 67784 262168 67786 262177
rect 67730 262103 67786 262112
rect 67640 260840 67692 260846
rect 67638 260808 67640 260817
rect 67692 260808 67694 260817
rect 67638 260743 67694 260752
rect 67730 258632 67786 258641
rect 67730 258567 67786 258576
rect 67744 258126 67772 258567
rect 67732 258120 67784 258126
rect 67732 258062 67784 258068
rect 67640 258052 67692 258058
rect 67640 257994 67692 258000
rect 67652 257961 67680 257994
rect 67638 257952 67694 257961
rect 67638 257887 67694 257896
rect 68006 256864 68062 256873
rect 68006 256799 68062 256808
rect 68020 256766 68048 256799
rect 68008 256760 68060 256766
rect 68008 256702 68060 256708
rect 67638 255368 67694 255377
rect 67638 255303 67640 255312
rect 67692 255303 67694 255312
rect 67640 255274 67692 255280
rect 67732 255264 67784 255270
rect 67730 255232 67732 255241
rect 67784 255232 67786 255241
rect 67640 255196 67692 255202
rect 67730 255167 67786 255176
rect 67640 255138 67692 255144
rect 67652 254833 67680 255138
rect 67638 254824 67694 254833
rect 67638 254759 67694 254768
rect 67640 253904 67692 253910
rect 67638 253872 67640 253881
rect 67692 253872 67694 253881
rect 67638 253807 67694 253816
rect 67638 251832 67694 251841
rect 67638 251767 67694 251776
rect 67652 251258 67680 251767
rect 68572 251433 68600 262890
rect 68558 251424 68614 251433
rect 68558 251359 68614 251368
rect 67640 251252 67692 251258
rect 67640 251194 67692 251200
rect 67732 251184 67784 251190
rect 67730 251152 67732 251161
rect 67784 251152 67786 251161
rect 67730 251087 67786 251096
rect 68466 249928 68522 249937
rect 68466 249863 68522 249872
rect 67638 249112 67694 249121
rect 67638 249047 67694 249056
rect 67652 248538 67680 249047
rect 67640 248532 67692 248538
rect 67640 248474 67692 248480
rect 67730 247752 67786 247761
rect 67730 247687 67786 247696
rect 67638 247208 67694 247217
rect 67744 247178 67772 247687
rect 67638 247143 67694 247152
rect 67732 247172 67784 247178
rect 67652 247110 67680 247143
rect 67732 247114 67784 247120
rect 67640 247104 67692 247110
rect 67640 247046 67692 247052
rect 67730 246392 67786 246401
rect 67730 246327 67786 246336
rect 67638 245848 67694 245857
rect 67638 245783 67694 245792
rect 67652 245750 67680 245783
rect 67640 245744 67692 245750
rect 67640 245686 67692 245692
rect 67744 245682 67772 246327
rect 67732 245676 67784 245682
rect 67732 245618 67784 245624
rect 67640 245608 67692 245614
rect 67640 245550 67692 245556
rect 67652 245313 67680 245550
rect 67638 245304 67694 245313
rect 67638 245239 67694 245248
rect 67732 244248 67784 244254
rect 67732 244190 67784 244196
rect 67640 244180 67692 244186
rect 67640 244122 67692 244128
rect 67652 243817 67680 244122
rect 67638 243808 67694 243817
rect 67638 243743 67694 243752
rect 67744 243681 67772 244190
rect 67730 243672 67786 243681
rect 67730 243607 67786 243616
rect 68480 243574 68508 249863
rect 68468 243568 68520 243574
rect 68468 243510 68520 243516
rect 68650 240952 68706 240961
rect 68650 240887 68706 240896
rect 68664 240106 68692 240887
rect 68652 240100 68704 240106
rect 68652 240042 68704 240048
rect 68756 236609 68784 272167
rect 68836 264988 68888 264994
rect 68836 264930 68888 264936
rect 68742 236600 68798 236609
rect 68742 236535 68798 236544
rect 68848 226953 68876 264930
rect 68940 262954 68968 295530
rect 69020 289196 69072 289202
rect 69020 289138 69072 289144
rect 68928 262948 68980 262954
rect 68928 262890 68980 262896
rect 68928 243568 68980 243574
rect 68928 243510 68980 243516
rect 68834 226944 68890 226953
rect 68834 226879 68890 226888
rect 68940 220114 68968 243510
rect 68928 220108 68980 220114
rect 68928 220050 68980 220056
rect 69032 186969 69060 289138
rect 69124 260273 69152 298114
rect 69204 295452 69256 295458
rect 69204 295394 69256 295400
rect 69216 281353 69244 295394
rect 70412 291977 70440 326334
rect 70504 302938 70532 337826
rect 71332 336394 71360 340068
rect 71976 336462 72004 340068
rect 73218 339810 73246 340068
rect 73172 339782 73246 339810
rect 73172 337770 73200 339782
rect 73908 339318 73936 340068
rect 73896 339312 73948 339318
rect 73896 339254 73948 339260
rect 73080 337742 73200 337770
rect 71964 336456 72016 336462
rect 71964 336398 72016 336404
rect 72424 336456 72476 336462
rect 72424 336398 72476 336404
rect 71320 336388 71372 336394
rect 71320 336330 71372 336336
rect 71332 319530 71360 336330
rect 71780 335164 71832 335170
rect 71780 335106 71832 335112
rect 71320 319524 71372 319530
rect 71320 319466 71372 319472
rect 71044 306468 71096 306474
rect 71044 306410 71096 306416
rect 70492 302932 70544 302938
rect 70492 302874 70544 302880
rect 70412 291949 70702 291977
rect 71056 291922 71084 306410
rect 71792 296002 71820 335106
rect 72436 312594 72464 336398
rect 73080 335170 73108 337742
rect 73068 335164 73120 335170
rect 73068 335106 73120 335112
rect 73804 332648 73856 332654
rect 73804 332590 73856 332596
rect 72424 312588 72476 312594
rect 72424 312530 72476 312536
rect 71780 295996 71832 296002
rect 71780 295938 71832 295944
rect 71320 294704 71372 294710
rect 71320 294646 71372 294652
rect 71332 291963 71360 294646
rect 71964 294636 72016 294642
rect 71964 294578 72016 294584
rect 71688 292392 71740 292398
rect 71686 292360 71688 292369
rect 71740 292360 71742 292369
rect 71686 292295 71742 292304
rect 71976 291963 72004 294578
rect 72608 294568 72660 294574
rect 72608 294510 72660 294516
rect 73250 294536 73306 294545
rect 72620 291963 72648 294510
rect 73250 294471 73306 294480
rect 73264 291963 73292 294471
rect 73816 292670 73844 332590
rect 73908 311234 73936 339254
rect 74552 337958 74580 340068
rect 75182 339960 75238 339969
rect 75840 339930 75868 340068
rect 75182 339895 75238 339904
rect 75828 339924 75880 339930
rect 74540 337952 74592 337958
rect 74540 337894 74592 337900
rect 74630 333296 74686 333305
rect 74630 333231 74686 333240
rect 73896 311228 73948 311234
rect 73896 311170 73948 311176
rect 74644 294250 74672 333231
rect 75196 316810 75224 339895
rect 75828 339866 75880 339872
rect 75276 337952 75328 337958
rect 75276 337894 75328 337900
rect 75288 323678 75316 337894
rect 75840 337550 75868 339866
rect 76484 339250 76512 340068
rect 76472 339244 76524 339250
rect 76472 339186 76524 339192
rect 76484 338230 76512 339186
rect 76472 338224 76524 338230
rect 76472 338166 76524 338172
rect 75828 337544 75880 337550
rect 75828 337486 75880 337492
rect 76564 337136 76616 337142
rect 76564 337078 76616 337084
rect 75276 323672 75328 323678
rect 75276 323614 75328 323620
rect 75276 322448 75328 322454
rect 75276 322390 75328 322396
rect 75184 316804 75236 316810
rect 75184 316746 75236 316752
rect 75288 306374 75316 322390
rect 75920 315308 75972 315314
rect 75920 315250 75972 315256
rect 75932 306374 75960 315250
rect 76576 314022 76604 337078
rect 76656 333872 76708 333878
rect 76656 333814 76708 333820
rect 76668 333470 76696 333814
rect 77128 333470 77156 340068
rect 78416 339522 78444 340068
rect 79076 339810 79104 340068
rect 79076 339782 79456 339810
rect 78404 339516 78456 339522
rect 78404 339458 78456 339464
rect 77484 338768 77536 338774
rect 77484 338710 77536 338716
rect 77404 336054 77432 336085
rect 77392 336048 77444 336054
rect 77390 336016 77392 336025
rect 77444 336016 77446 336025
rect 77390 335951 77446 335960
rect 76656 333464 76708 333470
rect 76656 333406 76708 333412
rect 77116 333464 77168 333470
rect 77116 333406 77168 333412
rect 76668 315353 76696 333406
rect 76654 315344 76710 315353
rect 76654 315279 76710 315288
rect 76564 314016 76616 314022
rect 76564 313958 76616 313964
rect 75288 306346 75408 306374
rect 75932 306346 76604 306374
rect 75000 297424 75052 297430
rect 75000 297366 75052 297372
rect 75012 294574 75040 297366
rect 75000 294568 75052 294574
rect 75000 294510 75052 294516
rect 74644 294222 75316 294250
rect 75184 294160 75236 294166
rect 75184 294102 75236 294108
rect 74540 294092 74592 294098
rect 74540 294034 74592 294040
rect 73804 292664 73856 292670
rect 73804 292606 73856 292612
rect 73896 292664 73948 292670
rect 73896 292606 73948 292612
rect 73908 291963 73936 292606
rect 74552 291963 74580 294034
rect 75196 291963 75224 294102
rect 75288 291938 75316 294222
rect 75380 292398 75408 306346
rect 76472 296744 76524 296750
rect 76472 296686 76524 296692
rect 75368 292392 75420 292398
rect 75368 292334 75420 292340
rect 76484 291963 76512 296686
rect 76576 291938 76604 306346
rect 77404 291977 77432 335951
rect 77496 306374 77524 338710
rect 78416 337482 78444 339458
rect 78404 337476 78456 337482
rect 78404 337418 78456 337424
rect 79428 332586 79456 339782
rect 79704 339425 79732 340068
rect 80946 339810 80974 340068
rect 80808 339782 80974 339810
rect 79690 339416 79746 339425
rect 79690 339351 79746 339360
rect 79704 338298 79732 339351
rect 79692 338292 79744 338298
rect 79692 338234 79744 338240
rect 80808 336734 80836 339782
rect 80796 336728 80848 336734
rect 80796 336670 80848 336676
rect 79416 332580 79468 332586
rect 79416 332522 79468 332528
rect 79324 323740 79376 323746
rect 79324 323682 79376 323688
rect 77496 306346 78076 306374
rect 77404 291949 77786 291977
rect 78048 291938 78076 306346
rect 79140 302320 79192 302326
rect 79140 302262 79192 302268
rect 79048 294228 79100 294234
rect 79048 294170 79100 294176
rect 79060 294030 79088 294170
rect 79048 294024 79100 294030
rect 79048 293966 79100 293972
rect 79060 291963 79088 293966
rect 79152 291938 79180 302262
rect 79336 296714 79364 323682
rect 79428 307086 79456 332522
rect 80704 323604 80756 323610
rect 80704 323546 80756 323552
rect 79416 307080 79468 307086
rect 79416 307022 79468 307028
rect 79244 296686 79364 296714
rect 79244 294234 79272 296686
rect 80336 295316 80388 295322
rect 80336 295258 80388 295264
rect 79232 294228 79284 294234
rect 79232 294170 79284 294176
rect 80348 291963 80376 295258
rect 80716 294545 80744 323546
rect 80808 320890 80836 336670
rect 81636 333810 81664 340068
rect 82280 339454 82308 340068
rect 82268 339448 82320 339454
rect 82268 339390 82320 339396
rect 83464 338224 83516 338230
rect 83464 338166 83516 338172
rect 82820 337340 82872 337346
rect 82820 337282 82872 337288
rect 82832 336598 82860 337282
rect 82820 336592 82872 336598
rect 82820 336534 82872 336540
rect 81624 333804 81676 333810
rect 81624 333746 81676 333752
rect 81636 332722 81664 333746
rect 81624 332716 81676 332722
rect 81624 332658 81676 332664
rect 82084 332716 82136 332722
rect 82084 332658 82136 332664
rect 80796 320884 80848 320890
rect 80796 320826 80848 320832
rect 82096 301578 82124 332658
rect 82084 301572 82136 301578
rect 82084 301514 82136 301520
rect 83476 298790 83504 338166
rect 83568 338026 83596 340068
rect 83648 338292 83700 338298
rect 83648 338234 83700 338240
rect 83556 338020 83608 338026
rect 83556 337962 83608 337968
rect 83556 313336 83608 313342
rect 83556 313278 83608 313284
rect 83464 298784 83516 298790
rect 83464 298726 83516 298732
rect 82268 298376 82320 298382
rect 82268 298318 82320 298324
rect 81622 294672 81678 294681
rect 81622 294607 81678 294616
rect 80702 294536 80758 294545
rect 80702 294471 80758 294480
rect 80978 292632 81034 292641
rect 80978 292567 81034 292576
rect 80992 291963 81020 292567
rect 81636 291963 81664 294607
rect 82280 291963 82308 298318
rect 83568 296714 83596 313278
rect 83660 305658 83688 338234
rect 84212 337822 84240 340068
rect 84856 339425 84884 340068
rect 84842 339416 84898 339425
rect 84842 339351 84898 339360
rect 84200 337816 84252 337822
rect 84200 337758 84252 337764
rect 84856 337346 84884 339351
rect 86144 337754 86172 340068
rect 86132 337748 86184 337754
rect 86132 337690 86184 337696
rect 84844 337340 84896 337346
rect 84844 337282 84896 337288
rect 86224 336048 86276 336054
rect 86224 335990 86276 335996
rect 85580 329112 85632 329118
rect 85580 329054 85632 329060
rect 84292 318164 84344 318170
rect 84292 318106 84344 318112
rect 84304 306374 84332 318106
rect 84304 306346 84976 306374
rect 83648 305652 83700 305658
rect 83648 305594 83700 305600
rect 84200 300892 84252 300898
rect 84200 300834 84252 300840
rect 83476 296686 83596 296714
rect 82912 294772 82964 294778
rect 82912 294714 82964 294720
rect 82924 291963 82952 294714
rect 83476 294710 83504 296686
rect 83556 295656 83608 295662
rect 83556 295598 83608 295604
rect 83464 294704 83516 294710
rect 83464 294646 83516 294652
rect 83568 291963 83596 295598
rect 84212 291963 84240 300834
rect 84844 294908 84896 294914
rect 84844 294850 84896 294856
rect 84856 291963 84884 294850
rect 84948 291977 84976 306346
rect 85592 294250 85620 329054
rect 86236 295322 86264 335990
rect 86316 335232 86368 335238
rect 86316 335174 86368 335180
rect 86328 334830 86356 335174
rect 86788 334830 86816 340068
rect 87432 339454 87460 340068
rect 88736 339810 88764 340068
rect 89318 339810 89346 340068
rect 88736 339782 89024 339810
rect 87420 339448 87472 339454
rect 87420 339390 87472 339396
rect 87696 339448 87748 339454
rect 87696 339390 87748 339396
rect 87604 338156 87656 338162
rect 87604 338098 87656 338104
rect 86868 337748 86920 337754
rect 86868 337690 86920 337696
rect 86880 337346 86908 337690
rect 86868 337340 86920 337346
rect 86868 337282 86920 337288
rect 86316 334824 86368 334830
rect 86316 334766 86368 334772
rect 86776 334824 86828 334830
rect 86776 334766 86828 334772
rect 86328 312662 86356 334766
rect 86316 312656 86368 312662
rect 86316 312598 86368 312604
rect 87616 304298 87644 338098
rect 87708 335306 87736 339390
rect 88996 336666 89024 339782
rect 89088 339782 89346 339810
rect 90024 339810 90052 340068
rect 90024 339782 90404 339810
rect 88984 336660 89036 336666
rect 88984 336602 89036 336608
rect 87696 335300 87748 335306
rect 87696 335242 87748 335248
rect 88340 326460 88392 326466
rect 88340 326402 88392 326408
rect 87604 304292 87656 304298
rect 87604 304234 87656 304240
rect 87604 302388 87656 302394
rect 87604 302330 87656 302336
rect 87512 299736 87564 299742
rect 87512 299678 87564 299684
rect 86224 295316 86276 295322
rect 86224 295258 86276 295264
rect 87420 294704 87472 294710
rect 87420 294646 87472 294652
rect 85592 294222 86264 294250
rect 86132 294160 86184 294166
rect 86132 294102 86184 294108
rect 84948 291949 85514 291977
rect 86144 291963 86172 294102
rect 86236 291977 86264 294222
rect 86236 291949 86802 291977
rect 87432 291963 87460 294646
rect 87524 291977 87552 299678
rect 87616 294166 87644 302330
rect 88352 296714 88380 326402
rect 88996 305697 89024 336602
rect 89088 333946 89116 339782
rect 90376 336530 90404 339782
rect 91296 337754 91324 340068
rect 91744 338768 91796 338774
rect 91744 338710 91796 338716
rect 91284 337748 91336 337754
rect 91284 337690 91336 337696
rect 91008 337408 91060 337414
rect 91008 337350 91060 337356
rect 90364 336524 90416 336530
rect 90364 336466 90416 336472
rect 89076 333940 89128 333946
rect 89076 333882 89128 333888
rect 89088 309806 89116 333882
rect 89720 310548 89772 310554
rect 89720 310490 89772 310496
rect 89076 309800 89128 309806
rect 89076 309742 89128 309748
rect 88982 305688 89038 305697
rect 88982 305623 89038 305632
rect 88352 296686 89024 296714
rect 88706 294808 88762 294817
rect 88706 294743 88762 294752
rect 87604 294160 87656 294166
rect 87604 294102 87656 294108
rect 87524 291949 88090 291977
rect 88720 291963 88748 294743
rect 88996 291977 89024 296686
rect 89732 291977 89760 310490
rect 90376 304366 90404 336466
rect 91020 314634 91048 337350
rect 91008 314628 91060 314634
rect 91008 314570 91060 314576
rect 90364 304360 90416 304366
rect 90364 304302 90416 304308
rect 90272 303680 90324 303686
rect 90272 303622 90324 303628
rect 90284 291977 90312 303622
rect 91282 298752 91338 298761
rect 91282 298687 91338 298696
rect 91296 298217 91324 298687
rect 91282 298208 91338 298217
rect 91282 298143 91338 298152
rect 88996 291949 89378 291977
rect 89732 291949 90022 291977
rect 90284 291949 90666 291977
rect 91296 291963 91324 298143
rect 91756 294914 91784 338710
rect 91940 337414 91968 340068
rect 92584 339386 92612 340068
rect 92572 339380 92624 339386
rect 92572 339322 92624 339328
rect 93124 339380 93176 339386
rect 93124 339322 93176 339328
rect 91928 337408 91980 337414
rect 91928 337350 91980 337356
rect 93136 308446 93164 339322
rect 93228 331226 93256 340068
rect 94516 332586 94544 340068
rect 95160 339386 95188 340068
rect 94596 339380 94648 339386
rect 94596 339322 94648 339328
rect 95148 339380 95200 339386
rect 95148 339322 95200 339328
rect 94504 332580 94556 332586
rect 94504 332522 94556 332528
rect 93216 331220 93268 331226
rect 93216 331162 93268 331168
rect 94608 329186 94636 339322
rect 95804 333985 95832 340068
rect 95790 333976 95846 333985
rect 95790 333911 95846 333920
rect 95804 332625 95832 333911
rect 95790 332616 95846 332625
rect 95790 332551 95846 332560
rect 96526 332616 96582 332625
rect 96526 332551 96582 332560
rect 94596 329180 94648 329186
rect 94596 329122 94648 329128
rect 95332 322244 95384 322250
rect 95332 322186 95384 322192
rect 93216 318232 93268 318238
rect 93216 318174 93268 318180
rect 93124 308440 93176 308446
rect 93124 308382 93176 308388
rect 93228 296714 93256 318174
rect 93952 316872 94004 316878
rect 93952 316814 94004 316820
rect 93964 306374 93992 316814
rect 93964 306346 94636 306374
rect 93860 298240 93912 298246
rect 93860 298182 93912 298188
rect 92952 296686 93256 296714
rect 91744 294908 91796 294914
rect 91744 294850 91796 294856
rect 91928 292868 91980 292874
rect 91928 292810 91980 292816
rect 91940 291963 91968 292810
rect 92952 292738 92980 296686
rect 93216 295520 93268 295526
rect 93216 295462 93268 295468
rect 92572 292732 92624 292738
rect 92572 292674 92624 292680
rect 92940 292732 92992 292738
rect 92940 292674 92992 292680
rect 92584 291963 92612 292674
rect 93228 291963 93256 295462
rect 93872 291963 93900 298182
rect 94504 294908 94556 294914
rect 94504 294850 94556 294856
rect 94516 291963 94544 294850
rect 94608 291938 94636 306346
rect 95344 291977 95372 322186
rect 96540 296041 96568 332551
rect 97092 331974 97120 340068
rect 97752 339810 97780 340068
rect 97752 339782 97948 339810
rect 97920 336530 97948 339782
rect 97908 336524 97960 336530
rect 97908 336466 97960 336472
rect 97816 332512 97868 332518
rect 97816 332454 97868 332460
rect 97828 331974 97856 332454
rect 97080 331968 97132 331974
rect 97080 331910 97132 331916
rect 97816 331968 97868 331974
rect 97816 331910 97868 331916
rect 97356 302932 97408 302938
rect 97356 302874 97408 302880
rect 97080 297492 97132 297498
rect 97080 297434 97132 297440
rect 97092 296818 97120 297434
rect 97080 296812 97132 296818
rect 97080 296754 97132 296760
rect 96526 296032 96582 296041
rect 96526 295967 96582 295976
rect 96436 292596 96488 292602
rect 96436 292538 96488 292544
rect 95344 291949 95818 291977
rect 96448 291963 96476 292538
rect 97092 291963 97120 296754
rect 97368 291938 97396 302874
rect 97828 302841 97856 331910
rect 97814 302832 97870 302841
rect 97814 302767 97870 302776
rect 97920 293185 97948 336466
rect 98380 334762 98408 340068
rect 98644 338836 98696 338842
rect 98644 338778 98696 338784
rect 98368 334756 98420 334762
rect 98368 334698 98420 334704
rect 98656 306374 98684 338778
rect 99668 337822 99696 340068
rect 99656 337816 99708 337822
rect 99656 337758 99708 337764
rect 98736 337476 98788 337482
rect 98736 337418 98788 337424
rect 98748 311137 98776 337418
rect 100312 336598 100340 340068
rect 100668 337816 100720 337822
rect 100668 337758 100720 337764
rect 100300 336592 100352 336598
rect 100300 336534 100352 336540
rect 99288 315376 99340 315382
rect 99288 315318 99340 315324
rect 98734 311128 98790 311137
rect 98734 311063 98790 311072
rect 98656 306346 98776 306374
rect 98552 301640 98604 301646
rect 98552 301582 98604 301588
rect 97906 293176 97962 293185
rect 97906 293111 97962 293120
rect 98368 292596 98420 292602
rect 98368 292538 98420 292544
rect 98380 291963 98408 292538
rect 98564 291938 98592 301582
rect 98748 292602 98776 306346
rect 99300 294098 99328 315318
rect 100680 310486 100708 337758
rect 100956 336734 100984 340068
rect 102198 339810 102226 340068
rect 102152 339782 102226 339810
rect 102152 337736 102180 339782
rect 102060 337708 102180 337736
rect 100944 336728 100996 336734
rect 100944 336670 100996 336676
rect 101956 336728 102008 336734
rect 101956 336670 102008 336676
rect 101404 319456 101456 319462
rect 101404 319398 101456 319404
rect 100668 310480 100720 310486
rect 100668 310422 100720 310428
rect 99380 305040 99432 305046
rect 99380 304982 99432 304988
rect 99288 294092 99340 294098
rect 99288 294034 99340 294040
rect 99300 293282 99328 294034
rect 99288 293276 99340 293282
rect 99288 293218 99340 293224
rect 98736 292596 98788 292602
rect 98736 292538 98788 292544
rect 99392 291977 99420 304982
rect 101416 294642 101444 319398
rect 101968 308582 101996 336670
rect 102060 335345 102088 337708
rect 102046 335336 102102 335345
rect 102046 335271 102102 335280
rect 101956 308576 102008 308582
rect 101956 308518 102008 308524
rect 102060 297401 102088 335271
rect 102888 317422 102916 340068
rect 103532 337482 103560 340068
rect 104820 337890 104848 340068
rect 105464 339250 105492 340068
rect 105452 339244 105504 339250
rect 105452 339186 105504 339192
rect 104808 337884 104860 337890
rect 104808 337826 104860 337832
rect 103612 337748 103664 337754
rect 103612 337690 103664 337696
rect 103520 337476 103572 337482
rect 103520 337418 103572 337424
rect 103060 337272 103112 337278
rect 103060 337214 103112 337220
rect 103072 334626 103100 337214
rect 103624 335209 103652 337690
rect 104164 337544 104216 337550
rect 104164 337486 104216 337492
rect 103610 335200 103666 335209
rect 103610 335135 103666 335144
rect 103060 334620 103112 334626
rect 103060 334562 103112 334568
rect 103612 327752 103664 327758
rect 103612 327694 103664 327700
rect 102876 317416 102928 317422
rect 102876 317358 102928 317364
rect 103624 316034 103652 327694
rect 103532 316006 103652 316034
rect 102140 299668 102192 299674
rect 102140 299610 102192 299616
rect 102046 297392 102102 297401
rect 102046 297327 102102 297336
rect 101404 294636 101456 294642
rect 101404 294578 101456 294584
rect 101588 294092 101640 294098
rect 101588 294034 101640 294040
rect 100944 294024 100996 294030
rect 100944 293966 100996 293972
rect 99392 291949 99682 291977
rect 100956 291963 100984 293966
rect 101600 291963 101628 294034
rect 102152 291977 102180 299610
rect 102876 296948 102928 296954
rect 102876 296890 102928 296896
rect 102152 291949 102258 291977
rect 102888 291963 102916 296890
rect 103532 291963 103560 316006
rect 103612 310480 103664 310486
rect 103612 310422 103664 310428
rect 103624 296714 103652 310422
rect 104176 304434 104204 337486
rect 104820 337278 104848 337826
rect 104808 337272 104860 337278
rect 104808 337214 104860 337220
rect 106108 336394 106136 340068
rect 106188 339244 106240 339250
rect 106188 339186 106240 339192
rect 106096 336388 106148 336394
rect 106096 336330 106148 336336
rect 104806 335200 104862 335209
rect 104806 335135 104862 335144
rect 104716 325032 104768 325038
rect 104716 324974 104768 324980
rect 104728 323746 104756 324974
rect 104716 323740 104768 323746
rect 104716 323682 104768 323688
rect 104820 307154 104848 335135
rect 104900 330812 104952 330818
rect 104900 330754 104952 330760
rect 104808 307148 104860 307154
rect 104808 307090 104860 307096
rect 104164 304428 104216 304434
rect 104164 304370 104216 304376
rect 103624 296686 104296 296714
rect 104162 294536 104218 294545
rect 104162 294471 104218 294480
rect 104176 291963 104204 294471
rect 104268 291977 104296 296686
rect 104912 294370 104940 330754
rect 106108 309874 106136 336330
rect 106096 309868 106148 309874
rect 106096 309810 106148 309816
rect 106200 308514 106228 339186
rect 107396 337550 107424 340068
rect 107476 339516 107528 339522
rect 107476 339458 107528 339464
rect 107384 337544 107436 337550
rect 107384 337486 107436 337492
rect 107488 322386 107516 339458
rect 108040 333946 108068 340068
rect 108028 333940 108080 333946
rect 108028 333882 108080 333888
rect 107568 333328 107620 333334
rect 107568 333270 107620 333276
rect 107476 322380 107528 322386
rect 107476 322322 107528 322328
rect 106188 308508 106240 308514
rect 106188 308450 106240 308456
rect 104992 300144 105044 300150
rect 104992 300086 105044 300092
rect 104900 294364 104952 294370
rect 104900 294306 104952 294312
rect 104268 291949 104834 291977
rect 105004 291938 105032 300086
rect 107292 297016 107344 297022
rect 107292 296958 107344 296964
rect 106740 294840 106792 294846
rect 106740 294782 106792 294788
rect 105820 294364 105872 294370
rect 105820 294306 105872 294312
rect 105832 291977 105860 294306
rect 105832 291949 106122 291977
rect 106752 291963 106780 294782
rect 107304 294778 107332 296958
rect 107292 294772 107344 294778
rect 107292 294714 107344 294720
rect 107580 292738 107608 333270
rect 108040 331906 108068 333882
rect 108028 331900 108080 331906
rect 108028 331842 108080 331848
rect 107752 327956 107804 327962
rect 107752 327898 107804 327904
rect 107658 327720 107714 327729
rect 107658 327655 107714 327664
rect 107672 294370 107700 327655
rect 107660 294364 107712 294370
rect 107660 294306 107712 294312
rect 107384 292732 107436 292738
rect 107384 292674 107436 292680
rect 107568 292732 107620 292738
rect 107568 292674 107620 292680
rect 107396 291963 107424 292674
rect 107764 291977 107792 327898
rect 108684 313342 108712 340068
rect 109972 337754 110000 340068
rect 109960 337748 110012 337754
rect 109960 337690 110012 337696
rect 110236 337544 110288 337550
rect 110236 337486 110288 337492
rect 110248 336841 110276 337486
rect 110234 336832 110290 336841
rect 110234 336767 110290 336776
rect 110616 336734 110644 340068
rect 111260 339697 111288 340068
rect 111246 339688 111302 339697
rect 111246 339623 111302 339632
rect 111064 339584 111116 339590
rect 111064 339526 111116 339532
rect 110604 336728 110656 336734
rect 110604 336670 110656 336676
rect 109040 334688 109092 334694
rect 109040 334630 109092 334636
rect 109052 333266 109080 334630
rect 109040 333260 109092 333266
rect 109040 333202 109092 333208
rect 111076 327826 111104 339526
rect 111064 327820 111116 327826
rect 111064 327762 111116 327768
rect 110328 325712 110380 325718
rect 110328 325654 110380 325660
rect 108672 313336 108724 313342
rect 108672 313278 108724 313284
rect 110340 300966 110368 325654
rect 111260 318102 111288 339623
rect 112548 338026 112576 340068
rect 113192 339318 113220 340068
rect 113180 339312 113232 339318
rect 113180 339254 113232 339260
rect 113732 339312 113784 339318
rect 113732 339254 113784 339260
rect 112536 338020 112588 338026
rect 112536 337962 112588 337968
rect 111800 337748 111852 337754
rect 111800 337690 111852 337696
rect 111812 337385 111840 337690
rect 111798 337376 111854 337385
rect 111798 337311 111854 337320
rect 111616 336796 111668 336802
rect 111616 336738 111668 336744
rect 111248 318096 111300 318102
rect 111248 318038 111300 318044
rect 111064 314696 111116 314702
rect 111064 314638 111116 314644
rect 111076 301646 111104 314638
rect 111628 302462 111656 336738
rect 111708 336728 111760 336734
rect 111708 336670 111760 336676
rect 111800 336728 111852 336734
rect 111800 336670 111852 336676
rect 111720 336462 111748 336670
rect 111708 336456 111760 336462
rect 111708 336398 111760 336404
rect 111156 302456 111208 302462
rect 111156 302398 111208 302404
rect 111616 302456 111668 302462
rect 111616 302398 111668 302404
rect 111064 301640 111116 301646
rect 111064 301582 111116 301588
rect 109684 300960 109736 300966
rect 109684 300902 109736 300908
rect 110328 300960 110380 300966
rect 110328 300902 110380 300908
rect 108396 294364 108448 294370
rect 108396 294306 108448 294312
rect 109316 294364 109368 294370
rect 109316 294306 109368 294312
rect 108408 291977 108436 294306
rect 107764 291949 108054 291977
rect 108408 291949 108698 291977
rect 109328 291963 109356 294306
rect 109696 291977 109724 300902
rect 111168 294914 111196 302398
rect 111248 294976 111300 294982
rect 111248 294918 111300 294924
rect 111156 294908 111208 294914
rect 111156 294850 111208 294856
rect 109696 291949 109986 291977
rect 111260 291963 111288 294918
rect 111720 293282 111748 336398
rect 111812 336394 111840 336670
rect 111800 336388 111852 336394
rect 111800 336330 111852 336336
rect 113744 335354 113772 339254
rect 113836 338094 113864 340068
rect 113824 338088 113876 338094
rect 113824 338030 113876 338036
rect 113836 336802 113864 338030
rect 113824 336796 113876 336802
rect 113824 336738 113876 336744
rect 113744 335326 113864 335354
rect 111800 330676 111852 330682
rect 111800 330618 111852 330624
rect 111708 293276 111760 293282
rect 111708 293218 111760 293224
rect 111812 291977 111840 330618
rect 112444 327820 112496 327826
rect 112444 327762 112496 327768
rect 112456 294370 112484 327762
rect 113836 318170 113864 335326
rect 115124 335306 115152 340068
rect 115112 335300 115164 335306
rect 115112 335242 115164 335248
rect 115124 334014 115152 335242
rect 115112 334008 115164 334014
rect 115112 333950 115164 333956
rect 115204 330744 115256 330750
rect 115204 330686 115256 330692
rect 114560 323672 114612 323678
rect 114560 323614 114612 323620
rect 113824 318164 113876 318170
rect 113824 318106 113876 318112
rect 113824 309868 113876 309874
rect 113824 309810 113876 309816
rect 113836 298450 113864 309810
rect 113824 298444 113876 298450
rect 113824 298386 113876 298392
rect 113836 296714 113864 298386
rect 113744 296686 113864 296714
rect 112444 294364 112496 294370
rect 112444 294306 112496 294312
rect 113744 291977 113772 296686
rect 114468 295996 114520 296002
rect 114468 295938 114520 295944
rect 113824 294636 113876 294642
rect 113824 294578 113876 294584
rect 111812 291949 111918 291977
rect 113206 291949 113772 291977
rect 113836 291963 113864 294578
rect 114480 291963 114508 295938
rect 114572 291977 114600 323614
rect 115216 292806 115244 330686
rect 115308 325718 115336 366959
rect 115860 353297 115888 371894
rect 115938 364304 115994 364313
rect 115938 364239 115994 364248
rect 115846 353288 115902 353297
rect 115846 353223 115902 353232
rect 115662 339824 115718 339833
rect 115662 339759 115718 339768
rect 115676 339590 115704 339759
rect 115664 339584 115716 339590
rect 115664 339526 115716 339532
rect 115768 338065 115796 340068
rect 115754 338056 115810 338065
rect 115754 337991 115810 338000
rect 115388 334008 115440 334014
rect 115388 333950 115440 333956
rect 115296 325712 115348 325718
rect 115296 325654 115348 325660
rect 115400 318238 115428 333950
rect 115952 333334 115980 364239
rect 116596 346390 116624 451522
rect 116676 392488 116728 392494
rect 116676 392430 116728 392436
rect 116688 392018 116716 392430
rect 116676 392012 116728 392018
rect 116676 391954 116728 391960
rect 116688 370025 116716 391954
rect 117424 379545 117452 485007
rect 117516 469878 117544 561002
rect 117608 551342 117636 587415
rect 118712 584066 118740 677622
rect 122932 677612 122984 677618
rect 122932 677554 122984 677560
rect 120356 676320 120408 676326
rect 120356 676262 120408 676268
rect 118792 666596 118844 666602
rect 118792 666538 118844 666544
rect 118620 584038 118740 584066
rect 118620 583522 118648 584038
rect 118700 583976 118752 583982
rect 118700 583918 118752 583924
rect 118712 583710 118740 583918
rect 118700 583704 118752 583710
rect 118700 583646 118752 583652
rect 118620 583494 118740 583522
rect 118712 580922 118740 583494
rect 118700 580916 118752 580922
rect 118700 580858 118752 580864
rect 118712 579737 118740 580858
rect 118698 579728 118754 579737
rect 118698 579663 118754 579672
rect 118804 576854 118832 666538
rect 119344 650140 119396 650146
rect 119344 650082 119396 650088
rect 119356 643754 119384 650082
rect 119344 643748 119396 643754
rect 119344 643690 119396 643696
rect 118884 636948 118936 636954
rect 118884 636890 118936 636896
rect 118896 618254 118924 636890
rect 120080 635724 120132 635730
rect 120080 635666 120132 635672
rect 118884 618248 118936 618254
rect 118884 618190 118936 618196
rect 118882 587208 118938 587217
rect 118882 587143 118938 587152
rect 118712 576826 118832 576854
rect 118712 569922 118740 576826
rect 118620 569894 118740 569922
rect 118620 568614 118648 569894
rect 118608 568608 118660 568614
rect 118608 568550 118660 568556
rect 117596 551336 117648 551342
rect 117596 551278 117648 551284
rect 117594 497448 117650 497457
rect 117594 497383 117650 497392
rect 117504 469872 117556 469878
rect 117504 469814 117556 469820
rect 117516 469334 117544 469814
rect 117504 469328 117556 469334
rect 117504 469270 117556 469276
rect 117504 463684 117556 463690
rect 117504 463626 117556 463632
rect 117516 384985 117544 463626
rect 117608 440910 117636 497383
rect 118620 477630 118648 568550
rect 118790 545184 118846 545193
rect 118790 545119 118846 545128
rect 118608 477624 118660 477630
rect 118608 477566 118660 477572
rect 118620 477426 118648 477566
rect 118700 477556 118752 477562
rect 118700 477498 118752 477504
rect 118608 477420 118660 477426
rect 118608 477362 118660 477368
rect 117688 469328 117740 469334
rect 117688 469270 117740 469276
rect 117596 440904 117648 440910
rect 117596 440846 117648 440852
rect 117594 396672 117650 396681
rect 117594 396607 117650 396616
rect 117502 384976 117558 384985
rect 117502 384911 117558 384920
rect 117410 379536 117466 379545
rect 117410 379471 117466 379480
rect 116674 370016 116730 370025
rect 116674 369951 116730 369960
rect 117318 365256 117374 365265
rect 117318 365191 117374 365200
rect 117332 364410 117360 365191
rect 117320 364404 117372 364410
rect 117320 364346 117372 364352
rect 117608 357105 117636 396607
rect 117700 362234 117728 469270
rect 118712 392494 118740 477498
rect 118804 459649 118832 545119
rect 118896 533526 118924 587143
rect 119528 583704 119580 583710
rect 119528 583646 119580 583652
rect 119344 580304 119396 580310
rect 119344 580246 119396 580252
rect 119356 538286 119384 580246
rect 119436 564460 119488 564466
rect 119436 564402 119488 564408
rect 119344 538280 119396 538286
rect 119344 538222 119396 538228
rect 119356 538082 119384 538222
rect 119344 538076 119396 538082
rect 119344 538018 119396 538024
rect 119448 537538 119476 564402
rect 119540 555558 119568 583646
rect 119528 555552 119580 555558
rect 119528 555494 119580 555500
rect 119436 537532 119488 537538
rect 119436 537474 119488 537480
rect 120092 536654 120120 635666
rect 120262 585304 120318 585313
rect 120262 585239 120318 585248
rect 120172 581732 120224 581738
rect 120172 581674 120224 581680
rect 120184 539374 120212 581674
rect 120172 539368 120224 539374
rect 120172 539310 120224 539316
rect 120080 536648 120132 536654
rect 120080 536590 120132 536596
rect 120092 536110 120120 536590
rect 120080 536104 120132 536110
rect 120080 536046 120132 536052
rect 119344 535492 119396 535498
rect 119344 535434 119396 535440
rect 118884 533520 118936 533526
rect 118884 533462 118936 533468
rect 118790 459640 118846 459649
rect 118790 459575 118846 459584
rect 118792 453348 118844 453354
rect 118792 453290 118844 453296
rect 118804 453257 118832 453290
rect 118790 453248 118846 453257
rect 118790 453183 118846 453192
rect 119356 438938 119384 535434
rect 120276 499574 120304 585239
rect 120368 579630 120396 676262
rect 121552 676252 121604 676258
rect 121552 676194 121604 676200
rect 121460 638376 121512 638382
rect 121460 638318 121512 638324
rect 120356 579624 120408 579630
rect 120356 579566 120408 579572
rect 121092 579624 121144 579630
rect 121092 579566 121144 579572
rect 121104 578338 121132 579566
rect 121092 578332 121144 578338
rect 121092 578274 121144 578280
rect 121472 538014 121500 638318
rect 121564 633010 121592 676194
rect 121644 655648 121696 655654
rect 121644 655590 121696 655596
rect 121552 633004 121604 633010
rect 121552 632946 121604 632952
rect 121552 632868 121604 632874
rect 121552 632810 121604 632816
rect 121460 538008 121512 538014
rect 121460 537950 121512 537956
rect 121472 536926 121500 537950
rect 121460 536920 121512 536926
rect 121460 536862 121512 536868
rect 121564 534818 121592 632810
rect 121656 558210 121684 655590
rect 122840 638920 122892 638926
rect 122840 638862 122892 638868
rect 121736 588600 121788 588606
rect 121736 588542 121788 588548
rect 121748 581641 121776 588542
rect 121734 581632 121790 581641
rect 121734 581567 121790 581576
rect 121736 581528 121788 581534
rect 121736 581470 121788 581476
rect 121644 558204 121696 558210
rect 121644 558146 121696 558152
rect 121552 534812 121604 534818
rect 121552 534754 121604 534760
rect 120724 530664 120776 530670
rect 120724 530606 120776 530612
rect 120092 499546 120304 499574
rect 120092 494018 120120 499546
rect 120080 494012 120132 494018
rect 120080 493954 120132 493960
rect 120092 493406 120120 493954
rect 120080 493400 120132 493406
rect 120080 493342 120132 493348
rect 120172 492108 120224 492114
rect 120172 492050 120224 492056
rect 120080 477624 120132 477630
rect 120080 477566 120132 477572
rect 119988 465044 120040 465050
rect 119988 464986 120040 464992
rect 119436 459672 119488 459678
rect 119436 459614 119488 459620
rect 119344 438932 119396 438938
rect 119344 438874 119396 438880
rect 119356 438666 119384 438874
rect 119344 438660 119396 438666
rect 119344 438602 119396 438608
rect 118792 394800 118844 394806
rect 118792 394742 118844 394748
rect 118804 394670 118832 394742
rect 118792 394664 118844 394670
rect 118792 394606 118844 394612
rect 118700 392488 118752 392494
rect 118700 392430 118752 392436
rect 119448 389638 119476 459614
rect 119620 398200 119672 398206
rect 119620 398142 119672 398148
rect 119436 389632 119488 389638
rect 119436 389574 119488 389580
rect 119344 388000 119396 388006
rect 119344 387942 119396 387948
rect 118514 384976 118570 384985
rect 118514 384911 118570 384920
rect 118528 384810 118556 384911
rect 118516 384804 118568 384810
rect 118516 384746 118568 384752
rect 118608 384396 118660 384402
rect 118608 384338 118660 384344
rect 118620 384305 118648 384338
rect 118606 384296 118662 384305
rect 118606 384231 118662 384240
rect 118606 383616 118662 383625
rect 118606 383551 118662 383560
rect 118620 383110 118648 383551
rect 118608 383104 118660 383110
rect 118608 383046 118660 383052
rect 118606 382256 118662 382265
rect 118606 382191 118608 382200
rect 118660 382191 118662 382200
rect 118608 382162 118660 382168
rect 118608 381608 118660 381614
rect 118606 381576 118608 381585
rect 118660 381576 118662 381585
rect 118606 381511 118662 381520
rect 118332 380180 118384 380186
rect 118332 380122 118384 380128
rect 118344 379545 118372 380122
rect 118330 379536 118386 379545
rect 118330 379471 118386 379480
rect 118606 378856 118662 378865
rect 118606 378791 118662 378800
rect 118620 378758 118648 378791
rect 118608 378752 118660 378758
rect 118608 378694 118660 378700
rect 118056 378208 118108 378214
rect 118054 378176 118056 378185
rect 118108 378176 118110 378185
rect 118054 378111 118110 378120
rect 118240 378140 118292 378146
rect 118240 378082 118292 378088
rect 118252 376825 118280 378082
rect 118238 376816 118294 376825
rect 118238 376751 118294 376760
rect 118148 376712 118200 376718
rect 118148 376654 118200 376660
rect 118160 375465 118188 376654
rect 118606 376136 118662 376145
rect 119356 376106 119384 387942
rect 119436 387864 119488 387870
rect 119436 387806 119488 387812
rect 119448 383042 119476 387806
rect 119436 383036 119488 383042
rect 119436 382978 119488 382984
rect 118606 376071 118662 376080
rect 119344 376100 119396 376106
rect 118146 375456 118202 375465
rect 118620 375426 118648 376071
rect 119344 376042 119396 376048
rect 118146 375391 118202 375400
rect 118608 375420 118660 375426
rect 118608 375362 118660 375368
rect 118608 373992 118660 373998
rect 119632 373994 119660 398142
rect 120000 394806 120028 464986
rect 119988 394800 120040 394806
rect 119988 394742 120040 394748
rect 120092 383654 120120 477566
rect 120184 422278 120212 492050
rect 120736 436150 120764 530606
rect 121458 498264 121514 498273
rect 121458 498199 121460 498208
rect 121512 498199 121514 498208
rect 121460 498170 121512 498176
rect 121460 474768 121512 474774
rect 121460 474710 121512 474716
rect 121472 474638 121500 474710
rect 121460 474632 121512 474638
rect 121460 474574 121512 474580
rect 121460 472116 121512 472122
rect 121460 472058 121512 472064
rect 121472 471986 121500 472058
rect 121460 471980 121512 471986
rect 121460 471922 121512 471928
rect 121656 465050 121684 558146
rect 121748 555422 121776 581470
rect 121736 555416 121788 555422
rect 121736 555358 121788 555364
rect 122852 537946 122880 638862
rect 122944 580990 122972 677554
rect 123024 669520 123076 669526
rect 123024 669462 123076 669468
rect 122932 580984 122984 580990
rect 122932 580926 122984 580932
rect 123036 574054 123064 669462
rect 124404 665236 124456 665242
rect 124404 665178 124456 665184
rect 124128 639600 124180 639606
rect 124128 639542 124180 639548
rect 124140 638926 124168 639542
rect 124128 638920 124180 638926
rect 124128 638862 124180 638868
rect 124312 638512 124364 638518
rect 124312 638454 124364 638460
rect 124220 638240 124272 638246
rect 124220 638182 124272 638188
rect 123116 584044 123168 584050
rect 123116 583986 123168 583992
rect 123024 574048 123076 574054
rect 123024 573990 123076 573996
rect 122930 572792 122986 572801
rect 122930 572727 122986 572736
rect 122944 540258 122972 572727
rect 122932 540252 122984 540258
rect 122932 540194 122984 540200
rect 122840 537940 122892 537946
rect 122840 537882 122892 537888
rect 122852 536858 122880 537882
rect 121736 536852 121788 536858
rect 121736 536794 121788 536800
rect 122840 536852 122892 536858
rect 122840 536794 122892 536800
rect 121644 465044 121696 465050
rect 121644 464986 121696 464992
rect 121460 463752 121512 463758
rect 121460 463694 121512 463700
rect 120264 436144 120316 436150
rect 120264 436086 120316 436092
rect 120724 436144 120776 436150
rect 120724 436086 120776 436092
rect 120276 436014 120304 436086
rect 120264 436008 120316 436014
rect 120264 435950 120316 435956
rect 120172 422272 120224 422278
rect 120172 422214 120224 422220
rect 120184 389910 120212 422214
rect 120264 392624 120316 392630
rect 120264 392566 120316 392572
rect 120276 392018 120304 392566
rect 120264 392012 120316 392018
rect 120264 391954 120316 391960
rect 120816 392012 120868 392018
rect 120816 391954 120868 391960
rect 120172 389904 120224 389910
rect 120172 389846 120224 389852
rect 120092 383626 120212 383654
rect 118608 373934 118660 373940
rect 119448 373966 119660 373994
rect 118620 373425 118648 373934
rect 118606 373416 118662 373425
rect 118606 373351 118662 373360
rect 117872 372768 117924 372774
rect 117870 372736 117872 372745
rect 117924 372736 117926 372745
rect 117870 372671 117926 372680
rect 117778 371376 117834 371385
rect 117778 371311 117834 371320
rect 117792 371278 117820 371311
rect 117780 371272 117832 371278
rect 117780 371214 117832 371220
rect 118606 370696 118662 370705
rect 118606 370631 118662 370640
rect 118620 370530 118648 370631
rect 118608 370524 118660 370530
rect 118608 370466 118660 370472
rect 118606 370016 118662 370025
rect 118662 369974 118740 370002
rect 118606 369951 118662 369960
rect 118424 369844 118476 369850
rect 118424 369786 118476 369792
rect 118436 368665 118464 369786
rect 118712 369170 118740 369974
rect 118700 369164 118752 369170
rect 118700 369106 118752 369112
rect 119344 368688 119396 368694
rect 118422 368656 118478 368665
rect 119344 368630 119396 368636
rect 118422 368591 118478 368600
rect 118606 367976 118662 367985
rect 118606 367911 118662 367920
rect 117780 367872 117832 367878
rect 117780 367814 117832 367820
rect 117792 367305 117820 367814
rect 118620 367810 118648 367911
rect 118608 367804 118660 367810
rect 118608 367746 118660 367752
rect 117778 367296 117834 367305
rect 117778 367231 117834 367240
rect 118148 367056 118200 367062
rect 118148 366998 118200 367004
rect 118160 365945 118188 366998
rect 118146 365936 118202 365945
rect 118146 365871 118202 365880
rect 118056 365696 118108 365702
rect 118056 365638 118108 365644
rect 118068 364585 118096 365638
rect 118054 364576 118110 364585
rect 118054 364511 118110 364520
rect 118148 364268 118200 364274
rect 118148 364210 118200 364216
rect 118160 363225 118188 364210
rect 118146 363216 118202 363225
rect 118146 363151 118202 363160
rect 117964 362908 118016 362914
rect 117964 362850 118016 362856
rect 117976 362545 118004 362850
rect 117962 362536 118018 362545
rect 117962 362471 118018 362480
rect 117688 362228 117740 362234
rect 117688 362170 117740 362176
rect 117700 361865 117728 362170
rect 117686 361856 117742 361865
rect 117686 361791 117742 361800
rect 118606 361176 118662 361185
rect 118606 361111 118662 361120
rect 118620 360874 118648 361111
rect 118608 360868 118660 360874
rect 118608 360810 118660 360816
rect 117962 360224 118018 360233
rect 117962 360159 118018 360168
rect 118148 360188 118200 360194
rect 117594 357096 117650 357105
rect 117594 357031 117650 357040
rect 117780 354068 117832 354074
rect 117780 354010 117832 354016
rect 117792 353705 117820 354010
rect 117778 353696 117834 353705
rect 117778 353631 117834 353640
rect 117412 351892 117464 351898
rect 117412 351834 117464 351840
rect 117424 351665 117452 351834
rect 117410 351656 117466 351665
rect 117410 351591 117466 351600
rect 117502 347712 117558 347721
rect 117502 347647 117558 347656
rect 116584 346384 116636 346390
rect 116584 346326 116636 346332
rect 117320 346384 117372 346390
rect 117320 346326 117372 346332
rect 117332 342145 117360 346326
rect 117318 342136 117374 342145
rect 117318 342071 117374 342080
rect 117320 340876 117372 340882
rect 117320 340818 117372 340824
rect 117332 340105 117360 340818
rect 117412 340808 117464 340814
rect 117410 340776 117412 340785
rect 117464 340776 117466 340785
rect 117410 340711 117466 340720
rect 117318 340096 117374 340105
rect 117318 340031 117374 340040
rect 117424 339522 117452 340711
rect 117412 339516 117464 339522
rect 117412 339458 117464 339464
rect 117516 339250 117544 347647
rect 117780 343596 117832 343602
rect 117780 343538 117832 343544
rect 117792 342825 117820 343538
rect 117778 342816 117834 342825
rect 117778 342751 117834 342760
rect 117504 339244 117556 339250
rect 117504 339186 117556 339192
rect 117226 337920 117282 337929
rect 117226 337855 117282 337864
rect 117240 336841 117268 337855
rect 117226 336832 117282 336841
rect 117226 336767 117282 336776
rect 115940 333328 115992 333334
rect 115940 333270 115992 333276
rect 115388 318232 115440 318238
rect 115388 318174 115440 318180
rect 116674 318064 116730 318073
rect 116674 317999 116730 318008
rect 115296 317484 115348 317490
rect 115296 317426 115348 317432
rect 115308 296002 115336 317426
rect 116688 316878 116716 317999
rect 116676 316872 116728 316878
rect 116676 316814 116728 316820
rect 116676 313948 116728 313954
rect 116676 313890 116728 313896
rect 116584 312656 116636 312662
rect 116584 312598 116636 312604
rect 115296 295996 115348 296002
rect 115296 295938 115348 295944
rect 115204 292800 115256 292806
rect 115204 292742 115256 292748
rect 115756 292800 115808 292806
rect 115756 292742 115808 292748
rect 114572 291949 115138 291977
rect 115768 291963 115796 292742
rect 116596 292097 116624 312598
rect 116688 296886 116716 313890
rect 116676 296880 116728 296886
rect 116676 296822 116728 296828
rect 116582 292088 116638 292097
rect 116582 292023 116638 292032
rect 116688 291977 116716 296822
rect 117240 296714 117268 336767
rect 117976 336530 118004 360159
rect 118148 360130 118200 360136
rect 118160 359145 118188 360130
rect 118606 359816 118662 359825
rect 118606 359751 118662 359760
rect 118620 359514 118648 359751
rect 118608 359508 118660 359514
rect 118608 359450 118660 359456
rect 118146 359136 118202 359145
rect 118146 359071 118202 359080
rect 118056 358760 118108 358766
rect 118056 358702 118108 358708
rect 118068 338094 118096 358702
rect 118606 358456 118662 358465
rect 118606 358391 118662 358400
rect 118620 358086 118648 358391
rect 118608 358080 118660 358086
rect 118608 358022 118660 358028
rect 118606 357096 118662 357105
rect 118606 357031 118662 357040
rect 118620 356794 118648 357031
rect 118608 356788 118660 356794
rect 118608 356730 118660 356736
rect 118606 356416 118662 356425
rect 118606 356351 118662 356360
rect 118620 356114 118648 356351
rect 118608 356108 118660 356114
rect 118608 356050 118660 356056
rect 118516 356040 118568 356046
rect 118516 355982 118568 355988
rect 118528 355745 118556 355982
rect 118514 355736 118570 355745
rect 118514 355671 118570 355680
rect 118608 354408 118660 354414
rect 118606 354376 118608 354385
rect 118660 354376 118662 354385
rect 118606 354311 118662 354320
rect 118608 351824 118660 351830
rect 118608 351766 118660 351772
rect 118620 350985 118648 351766
rect 118606 350976 118662 350985
rect 118606 350911 118662 350920
rect 118608 350532 118660 350538
rect 118608 350474 118660 350480
rect 118620 350305 118648 350474
rect 118606 350296 118662 350305
rect 118606 350231 118662 350240
rect 118608 349104 118660 349110
rect 118608 349046 118660 349052
rect 118516 349036 118568 349042
rect 118516 348978 118568 348984
rect 118528 348265 118556 348978
rect 118620 348945 118648 349046
rect 118606 348936 118662 348945
rect 118606 348871 118662 348880
rect 118514 348256 118570 348265
rect 118514 348191 118570 348200
rect 118606 347576 118662 347585
rect 118606 347511 118662 347520
rect 118620 347070 118648 347511
rect 118608 347064 118660 347070
rect 118608 347006 118660 347012
rect 118608 346384 118660 346390
rect 118608 346326 118660 346332
rect 118514 346216 118570 346225
rect 118514 346151 118570 346160
rect 118528 345098 118556 346151
rect 118620 345545 118648 346326
rect 118606 345536 118662 345545
rect 118606 345471 118662 345480
rect 118516 345092 118568 345098
rect 118516 345034 118568 345040
rect 118608 345024 118660 345030
rect 118608 344966 118660 344972
rect 118620 344865 118648 344966
rect 118606 344856 118662 344865
rect 118606 344791 118662 344800
rect 118606 343496 118662 343505
rect 118606 343431 118662 343440
rect 118620 342922 118648 343431
rect 118608 342916 118660 342922
rect 118608 342858 118660 342864
rect 118514 342136 118570 342145
rect 118514 342071 118570 342080
rect 118148 341624 118200 341630
rect 118148 341566 118200 341572
rect 118056 338088 118108 338094
rect 118056 338030 118108 338036
rect 117964 336524 118016 336530
rect 117964 336466 118016 336472
rect 118160 332518 118188 341566
rect 118528 341562 118556 342071
rect 118516 341556 118568 341562
rect 118516 341498 118568 341504
rect 118148 332512 118200 332518
rect 118148 332454 118200 332460
rect 117872 303748 117924 303754
rect 117872 303690 117924 303696
rect 117884 300830 117912 303690
rect 117872 300824 117924 300830
rect 117872 300766 117924 300772
rect 117964 300212 118016 300218
rect 117964 300154 118016 300160
rect 117976 299606 118004 300154
rect 117964 299600 118016 299606
rect 117964 299542 118016 299548
rect 117148 296686 117268 296714
rect 117044 295316 117096 295322
rect 117044 295258 117096 295264
rect 116426 291949 116716 291977
rect 117056 291963 117084 295258
rect 117148 293321 117176 296686
rect 117228 295384 117280 295390
rect 117228 295326 117280 295332
rect 117240 294710 117268 295326
rect 117228 294704 117280 294710
rect 117228 294646 117280 294652
rect 117688 294704 117740 294710
rect 117688 294646 117740 294652
rect 117134 293312 117190 293321
rect 117134 293247 117190 293256
rect 117504 292868 117556 292874
rect 117504 292810 117556 292816
rect 71044 291916 71096 291922
rect 75288 291910 75842 291938
rect 76576 291910 77130 291938
rect 78048 291910 78418 291938
rect 79152 291910 79706 291938
rect 94608 291910 95162 291938
rect 97368 291910 97738 291938
rect 98564 291910 99026 291938
rect 105004 291910 105466 291938
rect 117516 291922 117544 292810
rect 117700 291963 117728 294646
rect 117976 291938 118004 299542
rect 118974 295216 119030 295225
rect 118974 295151 119030 295160
rect 118700 294024 118752 294030
rect 118700 293966 118752 293972
rect 110880 291916 110932 291922
rect 71044 291858 71096 291864
rect 110630 291864 110880 291870
rect 112812 291916 112864 291922
rect 110630 291858 110932 291864
rect 112562 291864 112812 291870
rect 112562 291858 112864 291864
rect 117504 291916 117556 291922
rect 117976 291910 118346 291938
rect 118712 291922 118740 293966
rect 118988 291963 119016 295151
rect 119356 294817 119384 368630
rect 119448 360602 119476 373966
rect 120080 371884 120132 371890
rect 120080 371826 120132 371832
rect 120092 367878 120120 371826
rect 120184 370530 120212 383626
rect 120172 370524 120224 370530
rect 120172 370466 120224 370472
rect 120080 367872 120132 367878
rect 120080 367814 120132 367820
rect 119528 364472 119580 364478
rect 119528 364414 119580 364420
rect 119436 360596 119488 360602
rect 119436 360538 119488 360544
rect 119448 337958 119476 360538
rect 119436 337952 119488 337958
rect 119436 337894 119488 337900
rect 119342 294808 119398 294817
rect 119342 294743 119398 294752
rect 119540 294681 119568 364414
rect 119710 361584 119766 361593
rect 119710 361519 119766 361528
rect 119724 337929 119752 361519
rect 120724 359508 120776 359514
rect 120724 359450 120776 359456
rect 119710 337920 119766 337929
rect 119710 337855 119766 337864
rect 120080 311228 120132 311234
rect 120080 311170 120132 311176
rect 120092 310486 120120 311170
rect 120080 310480 120132 310486
rect 120080 310422 120132 310428
rect 120080 305720 120132 305726
rect 120080 305662 120132 305668
rect 119620 294772 119672 294778
rect 119620 294714 119672 294720
rect 119526 294672 119582 294681
rect 119526 294607 119582 294616
rect 119632 291924 119660 294714
rect 118700 291916 118752 291922
rect 117504 291858 117556 291864
rect 118700 291858 118752 291864
rect 110630 291842 110920 291858
rect 112562 291842 112852 291858
rect 69768 291230 70058 291258
rect 69768 289202 69796 291230
rect 69756 289196 69808 289202
rect 69756 289138 69808 289144
rect 69202 281344 69258 281353
rect 69202 281279 69258 281288
rect 69110 260264 69166 260273
rect 69110 260199 69166 260208
rect 69202 255912 69258 255921
rect 69202 255847 69258 255856
rect 69110 244352 69166 244361
rect 69110 244287 69166 244296
rect 69124 202230 69152 244287
rect 69216 231198 69244 255847
rect 120092 249665 120120 305662
rect 120736 287065 120764 359450
rect 120828 331226 120856 391954
rect 120908 389632 120960 389638
rect 120908 389574 120960 389580
rect 120920 350606 120948 389574
rect 121000 369232 121052 369238
rect 121000 369174 121052 369180
rect 121012 358766 121040 369174
rect 121000 358760 121052 358766
rect 121000 358702 121052 358708
rect 121472 354414 121500 463694
rect 121550 456104 121606 456113
rect 121550 456039 121552 456048
rect 121604 456039 121606 456048
rect 121552 456010 121604 456016
rect 121748 439385 121776 536794
rect 122838 494728 122894 494737
rect 122838 494663 122894 494672
rect 122748 474632 122800 474638
rect 122748 474574 122800 474580
rect 121550 439376 121606 439385
rect 121550 439311 121606 439320
rect 121734 439376 121790 439385
rect 121734 439311 121790 439320
rect 121564 439142 121592 439311
rect 121552 439136 121604 439142
rect 121552 439078 121604 439084
rect 121552 388680 121604 388686
rect 121552 388622 121604 388628
rect 121564 387870 121592 388622
rect 121552 387864 121604 387870
rect 121550 387832 121552 387841
rect 121604 387832 121606 387841
rect 121550 387767 121606 387776
rect 121552 386028 121604 386034
rect 121552 385970 121604 385976
rect 121564 385150 121592 385970
rect 121552 385144 121604 385150
rect 121552 385086 121604 385092
rect 121460 354408 121512 354414
rect 121460 354350 121512 354356
rect 121472 354006 121500 354350
rect 121460 354000 121512 354006
rect 121460 353942 121512 353948
rect 120908 350600 120960 350606
rect 120908 350542 120960 350548
rect 121564 336054 121592 385086
rect 122656 385076 122708 385082
rect 122656 385018 122708 385024
rect 121644 360868 121696 360874
rect 121644 360810 121696 360816
rect 121656 338774 121684 360810
rect 121644 338768 121696 338774
rect 121644 338710 121696 338716
rect 121552 336048 121604 336054
rect 121552 335990 121604 335996
rect 122668 331294 122696 385018
rect 122760 367810 122788 474574
rect 122852 398138 122880 494663
rect 123128 493338 123156 583986
rect 123576 578332 123628 578338
rect 123576 578274 123628 578280
rect 123484 536852 123536 536858
rect 123484 536794 123536 536800
rect 123116 493332 123168 493338
rect 123116 493274 123168 493280
rect 123496 444446 123524 536794
rect 123588 488578 123616 578274
rect 124232 536518 124260 638182
rect 124324 540870 124352 638454
rect 124416 568546 124444 665178
rect 125600 635588 125652 635594
rect 125600 635530 125652 635536
rect 124496 582412 124548 582418
rect 124496 582354 124548 582360
rect 124404 568540 124456 568546
rect 124404 568482 124456 568488
rect 124312 540864 124364 540870
rect 124312 540806 124364 540812
rect 124220 536512 124272 536518
rect 124220 536454 124272 536460
rect 124232 535498 124260 536454
rect 124220 535492 124272 535498
rect 124220 535434 124272 535440
rect 124220 533384 124272 533390
rect 124220 533326 124272 533332
rect 123576 488572 123628 488578
rect 123576 488514 123628 488520
rect 124128 487280 124180 487286
rect 124128 487222 124180 487228
rect 124140 487082 124168 487222
rect 124128 487076 124180 487082
rect 124128 487018 124180 487024
rect 123576 448724 123628 448730
rect 123576 448666 123628 448672
rect 123484 444440 123536 444446
rect 123484 444382 123536 444388
rect 122840 398132 122892 398138
rect 122840 398074 122892 398080
rect 122840 394800 122892 394806
rect 122840 394742 122892 394748
rect 122748 367804 122800 367810
rect 122748 367746 122800 367752
rect 122852 358086 122880 394742
rect 123588 372026 123616 448666
rect 123668 386640 123720 386646
rect 123668 386582 123720 386588
rect 123576 372020 123628 372026
rect 123576 371962 123628 371968
rect 123484 367124 123536 367130
rect 123484 367066 123536 367072
rect 122840 358080 122892 358086
rect 122840 358022 122892 358028
rect 122196 331288 122248 331294
rect 122196 331230 122248 331236
rect 122656 331288 122708 331294
rect 122656 331230 122708 331236
rect 120816 331220 120868 331226
rect 120816 331162 120868 331168
rect 122104 327888 122156 327894
rect 122104 327830 122156 327836
rect 120816 310480 120868 310486
rect 120816 310422 120868 310428
rect 120828 289785 120856 310422
rect 121460 291984 121512 291990
rect 121460 291926 121512 291932
rect 121472 291825 121500 291926
rect 121458 291816 121514 291825
rect 121458 291751 121514 291760
rect 121550 291136 121606 291145
rect 121550 291071 121606 291080
rect 121458 290456 121514 290465
rect 121458 290391 121514 290400
rect 121472 289882 121500 290391
rect 121564 289950 121592 291071
rect 121552 289944 121604 289950
rect 121552 289886 121604 289892
rect 121460 289876 121512 289882
rect 121460 289818 121512 289824
rect 121552 289808 121604 289814
rect 120814 289776 120870 289785
rect 121552 289750 121604 289756
rect 120814 289711 120870 289720
rect 121564 289105 121592 289750
rect 121550 289096 121606 289105
rect 121550 289031 121606 289040
rect 121458 288416 121514 288425
rect 121458 288351 121460 288360
rect 121512 288351 121514 288360
rect 121460 288322 121512 288328
rect 121552 288312 121604 288318
rect 121552 288254 121604 288260
rect 121564 287745 121592 288254
rect 121550 287736 121606 287745
rect 121550 287671 121606 287680
rect 120722 287056 120778 287065
rect 120722 286991 120778 287000
rect 121552 287020 121604 287026
rect 120736 285734 120764 286991
rect 121552 286962 121604 286968
rect 120724 285728 120776 285734
rect 121564 285705 121592 286962
rect 120724 285670 120776 285676
rect 121550 285696 121606 285705
rect 121460 285660 121512 285666
rect 121550 285631 121606 285640
rect 121460 285602 121512 285608
rect 121472 285025 121500 285602
rect 121552 285592 121604 285598
rect 121552 285534 121604 285540
rect 121458 285016 121514 285025
rect 121458 284951 121514 284960
rect 121564 284345 121592 285534
rect 121550 284336 121606 284345
rect 121460 284300 121512 284306
rect 121550 284271 121606 284280
rect 121460 284242 121512 284248
rect 121472 283665 121500 284242
rect 121458 283656 121514 283665
rect 121458 283591 121514 283600
rect 121458 282976 121514 282985
rect 121458 282911 121460 282920
rect 121512 282911 121514 282920
rect 121460 282882 121512 282888
rect 121458 281616 121514 281625
rect 121458 281551 121460 281560
rect 121512 281551 121514 281560
rect 121460 281522 121512 281528
rect 121552 281512 121604 281518
rect 121552 281454 121604 281460
rect 121564 280945 121592 281454
rect 121550 280936 121606 280945
rect 121550 280871 121606 280880
rect 121458 280256 121514 280265
rect 121458 280191 121460 280200
rect 121512 280191 121514 280200
rect 121460 280162 121512 280168
rect 121552 280152 121604 280158
rect 121552 280094 121604 280100
rect 121564 279585 121592 280094
rect 121550 279576 121606 279585
rect 121550 279511 121606 279520
rect 121458 278896 121514 278905
rect 121458 278831 121514 278840
rect 121472 278798 121500 278831
rect 121460 278792 121512 278798
rect 121460 278734 121512 278740
rect 121552 278724 121604 278730
rect 121552 278666 121604 278672
rect 121564 278225 121592 278666
rect 121550 278216 121606 278225
rect 121550 278151 121606 278160
rect 120814 277536 120870 277545
rect 120814 277471 120870 277480
rect 120722 269376 120778 269385
rect 120722 269311 120778 269320
rect 120632 251184 120684 251190
rect 120632 251126 120684 251132
rect 120644 251025 120672 251126
rect 120170 251016 120226 251025
rect 120170 250951 120226 250960
rect 120630 251016 120686 251025
rect 120630 250951 120686 250960
rect 120078 249656 120134 249665
rect 120078 249591 120134 249600
rect 120092 248470 120120 249591
rect 120080 248464 120132 248470
rect 120080 248406 120132 248412
rect 120080 246356 120132 246362
rect 120080 246298 120132 246304
rect 69846 241632 69902 241641
rect 69846 241567 69902 241576
rect 69860 239494 69888 241567
rect 119988 240168 120040 240174
rect 69952 240094 70058 240122
rect 119646 240094 119752 240122
rect 119988 240110 120040 240116
rect 69848 239488 69900 239494
rect 69848 239430 69900 239436
rect 69952 238474 69980 240094
rect 70400 239828 70452 239834
rect 70400 239770 70452 239776
rect 69940 238468 69992 238474
rect 69940 238410 69992 238416
rect 69204 231192 69256 231198
rect 69204 231134 69256 231140
rect 69112 202224 69164 202230
rect 69112 202166 69164 202172
rect 70412 195430 70440 239770
rect 70688 238754 70716 240037
rect 71320 239834 71348 240037
rect 71780 239964 71832 239970
rect 71780 239906 71832 239912
rect 71308 239828 71360 239834
rect 71308 239770 71360 239776
rect 70504 238726 70716 238754
rect 70504 223514 70532 238726
rect 71792 233209 71820 239906
rect 71976 238202 72004 240037
rect 72620 238678 72648 240037
rect 72608 238672 72660 238678
rect 72608 238614 72660 238620
rect 71964 238196 72016 238202
rect 71964 238138 72016 238144
rect 73264 238134 73292 240037
rect 73896 239850 73924 240037
rect 73816 239822 73924 239850
rect 72424 238128 72476 238134
rect 72424 238070 72476 238076
rect 73252 238128 73304 238134
rect 73252 238070 73304 238076
rect 71778 233200 71834 233209
rect 71778 233135 71834 233144
rect 70492 223508 70544 223514
rect 70492 223450 70544 223456
rect 70400 195424 70452 195430
rect 70400 195366 70452 195372
rect 72436 191146 72464 238070
rect 73816 222018 73844 239822
rect 74552 238754 74580 240037
rect 74552 238726 74672 238754
rect 74540 233912 74592 233918
rect 74540 233854 74592 233860
rect 73804 222012 73856 222018
rect 73804 221954 73856 221960
rect 74552 213382 74580 233854
rect 74644 226166 74672 238726
rect 75196 233918 75224 240037
rect 75840 234433 75868 240037
rect 75920 239828 75972 239834
rect 75920 239770 75972 239776
rect 75826 234424 75882 234433
rect 75826 234359 75882 234368
rect 75184 233912 75236 233918
rect 75184 233854 75236 233860
rect 74632 226160 74684 226166
rect 74632 226102 74684 226108
rect 75932 224738 75960 239770
rect 76484 238754 76512 240037
rect 77116 239834 77144 240037
rect 77104 239828 77156 239834
rect 77104 239770 77156 239776
rect 77300 239828 77352 239834
rect 77300 239770 77352 239776
rect 76564 239488 76616 239494
rect 76564 239430 76616 239436
rect 76024 238726 76512 238754
rect 76024 230450 76052 238726
rect 76012 230444 76064 230450
rect 76012 230386 76064 230392
rect 75920 224732 75972 224738
rect 75920 224674 75972 224680
rect 74540 213376 74592 213382
rect 74540 213318 74592 213324
rect 72424 191140 72476 191146
rect 72424 191082 72476 191088
rect 76576 189922 76604 239430
rect 77312 217462 77340 239770
rect 77772 238754 77800 240037
rect 78404 239834 78432 240037
rect 78392 239828 78444 239834
rect 78392 239770 78444 239776
rect 79060 238754 79088 240037
rect 79704 238754 79732 240037
rect 80348 238754 80376 240037
rect 77404 238726 77800 238754
rect 78692 238726 79088 238754
rect 79244 238726 79732 238754
rect 80072 238726 80376 238754
rect 77404 228954 77432 238726
rect 77392 228948 77444 228954
rect 77392 228890 77444 228896
rect 77300 217456 77352 217462
rect 77300 217398 77352 217404
rect 78692 195294 78720 238726
rect 78864 238196 78916 238202
rect 78864 238138 78916 238144
rect 78876 230382 78904 238138
rect 78864 230376 78916 230382
rect 78864 230318 78916 230324
rect 79244 222086 79272 238726
rect 80072 226302 80100 238726
rect 80992 237454 81020 240037
rect 80980 237448 81032 237454
rect 80980 237390 81032 237396
rect 81636 234462 81664 240037
rect 82084 239420 82136 239426
rect 82084 239362 82136 239368
rect 81624 234456 81676 234462
rect 81624 234398 81676 234404
rect 80060 226296 80112 226302
rect 80060 226238 80112 226244
rect 82096 223582 82124 239362
rect 82280 238746 82308 240037
rect 82924 238882 82952 240037
rect 82912 238876 82964 238882
rect 82912 238818 82964 238824
rect 83568 238746 83596 240037
rect 82268 238740 82320 238746
rect 82268 238682 82320 238688
rect 83556 238740 83608 238746
rect 83556 238682 83608 238688
rect 83464 238128 83516 238134
rect 83464 238070 83516 238076
rect 82084 223576 82136 223582
rect 82084 223518 82136 223524
rect 79232 222080 79284 222086
rect 79232 222022 79284 222028
rect 83476 215218 83504 238070
rect 83568 229770 83596 238682
rect 84212 233986 84240 240037
rect 84292 239828 84344 239834
rect 84292 239770 84344 239776
rect 84200 233980 84252 233986
rect 84200 233922 84252 233928
rect 84304 233866 84332 239770
rect 84856 238754 84884 240037
rect 85488 239834 85516 240037
rect 85476 239828 85528 239834
rect 85476 239770 85528 239776
rect 85672 238944 85724 238950
rect 85672 238886 85724 238892
rect 84212 233838 84332 233866
rect 84396 238726 84884 238754
rect 83556 229764 83608 229770
rect 83556 229706 83608 229712
rect 83464 215212 83516 215218
rect 83464 215154 83516 215160
rect 78680 195288 78732 195294
rect 78680 195230 78732 195236
rect 76564 189916 76616 189922
rect 76564 189858 76616 189864
rect 84212 188426 84240 233838
rect 84292 233776 84344 233782
rect 84292 233718 84344 233724
rect 84304 219366 84332 233718
rect 84396 220658 84424 238726
rect 85684 235890 85712 238886
rect 86144 237386 86172 240037
rect 86788 238950 86816 240037
rect 86960 239828 87012 239834
rect 86960 239770 87012 239776
rect 86776 238944 86828 238950
rect 86776 238886 86828 238892
rect 86224 237448 86276 237454
rect 86224 237390 86276 237396
rect 86132 237380 86184 237386
rect 86132 237322 86184 237328
rect 86144 237153 86172 237322
rect 86130 237144 86186 237153
rect 86130 237079 86186 237088
rect 85672 235884 85724 235890
rect 85672 235826 85724 235832
rect 84384 220652 84436 220658
rect 84384 220594 84436 220600
rect 84292 219360 84344 219366
rect 84292 219302 84344 219308
rect 86236 210526 86264 237390
rect 86224 210520 86276 210526
rect 86224 210462 86276 210468
rect 86972 200870 87000 239770
rect 87432 238754 87460 240037
rect 88064 239834 88092 240037
rect 88052 239828 88104 239834
rect 88052 239770 88104 239776
rect 87064 238726 87460 238754
rect 87064 227594 87092 238726
rect 88720 238678 88748 240037
rect 88708 238672 88760 238678
rect 88708 238614 88760 238620
rect 88984 238060 89036 238066
rect 88984 238002 89036 238008
rect 87052 227588 87104 227594
rect 87052 227530 87104 227536
rect 88996 219434 89024 238002
rect 89364 235890 89392 240037
rect 90008 238754 90036 240037
rect 90640 239850 90668 240037
rect 89732 238726 90036 238754
rect 90560 239822 90668 239850
rect 89352 235884 89404 235890
rect 89352 235826 89404 235832
rect 88984 219428 89036 219434
rect 88984 219370 89036 219376
rect 89732 207806 89760 238726
rect 90560 229770 90588 239822
rect 91296 235686 91324 240037
rect 91940 238754 91968 240037
rect 92480 239828 92532 239834
rect 92480 239770 92532 239776
rect 91756 238726 91968 238754
rect 91284 235680 91336 235686
rect 91284 235622 91336 235628
rect 91756 234530 91784 238726
rect 91744 234524 91796 234530
rect 91744 234466 91796 234472
rect 91756 231849 91784 234466
rect 91742 231840 91798 231849
rect 91742 231775 91798 231784
rect 90548 229764 90600 229770
rect 90548 229706 90600 229712
rect 89720 207800 89772 207806
rect 89720 207742 89772 207748
rect 92492 206990 92520 239770
rect 92584 221610 92612 240037
rect 93216 239834 93244 240037
rect 93204 239828 93256 239834
rect 93204 239770 93256 239776
rect 92572 221604 92624 221610
rect 92572 221546 92624 221552
rect 93872 217530 93900 240037
rect 94516 238754 94544 240037
rect 93964 238726 94544 238754
rect 93964 220726 93992 238726
rect 95160 234530 95188 240037
rect 95240 239828 95292 239834
rect 95240 239770 95292 239776
rect 95148 234524 95200 234530
rect 95148 234466 95200 234472
rect 93952 220720 94004 220726
rect 93952 220662 94004 220668
rect 93860 217524 93912 217530
rect 93860 217466 93912 217472
rect 95252 208350 95280 239770
rect 95804 237250 95832 240037
rect 96436 239834 96464 240037
rect 96424 239828 96476 239834
rect 96424 239770 96476 239776
rect 97092 238754 97120 240037
rect 96632 238726 97120 238754
rect 95792 237244 95844 237250
rect 95792 237186 95844 237192
rect 96632 227050 96660 238726
rect 97736 235822 97764 240037
rect 98380 235958 98408 240037
rect 99012 239850 99040 240037
rect 98932 239822 99040 239850
rect 99380 239828 99432 239834
rect 98368 235952 98420 235958
rect 98368 235894 98420 235900
rect 97724 235816 97776 235822
rect 97724 235758 97776 235764
rect 96620 227044 96672 227050
rect 96620 226986 96672 226992
rect 98932 219434 98960 239822
rect 99380 239770 99432 239776
rect 98012 219406 98960 219434
rect 95240 208344 95292 208350
rect 95240 208286 95292 208292
rect 92480 206984 92532 206990
rect 92480 206926 92532 206932
rect 98012 204270 98040 219406
rect 98000 204264 98052 204270
rect 98000 204206 98052 204212
rect 99392 203658 99420 239770
rect 99668 238754 99696 240037
rect 100300 239834 100328 240037
rect 100944 239850 100972 240037
rect 100288 239828 100340 239834
rect 100288 239770 100340 239776
rect 100760 239828 100812 239834
rect 100760 239770 100812 239776
rect 100864 239822 100972 239850
rect 101588 239834 101616 240037
rect 101576 239828 101628 239834
rect 99484 238726 99696 238754
rect 99484 231810 99512 238726
rect 99472 231804 99524 231810
rect 99472 231746 99524 231752
rect 100772 206446 100800 239770
rect 100864 224262 100892 239822
rect 101576 239770 101628 239776
rect 102140 239828 102192 239834
rect 102140 239770 102192 239776
rect 100852 224256 100904 224262
rect 100852 224198 100904 224204
rect 100760 206440 100812 206446
rect 100760 206382 100812 206388
rect 99380 203652 99432 203658
rect 99380 203594 99432 203600
rect 86960 200864 87012 200870
rect 86960 200806 87012 200812
rect 102152 198150 102180 239770
rect 102244 213926 102272 240037
rect 102876 239834 102904 240037
rect 102864 239828 102916 239834
rect 102864 239770 102916 239776
rect 103532 235754 103560 240037
rect 104176 239442 104204 240037
rect 104808 239850 104836 240037
rect 103624 239414 104204 239442
rect 104728 239822 104836 239850
rect 103520 235748 103572 235754
rect 103520 235690 103572 235696
rect 103624 231130 103652 239414
rect 104728 238754 104756 239822
rect 105464 238754 105492 240037
rect 103716 238726 104756 238754
rect 104912 238726 105492 238754
rect 103612 231124 103664 231130
rect 103612 231066 103664 231072
rect 103716 215286 103744 238726
rect 104164 231192 104216 231198
rect 104164 231134 104216 231140
rect 103704 215280 103756 215286
rect 103704 215222 103756 215228
rect 102232 213920 102284 213926
rect 102232 213862 102284 213868
rect 104176 199578 104204 231134
rect 104912 209778 104940 238726
rect 106108 235958 106136 240037
rect 106096 235952 106148 235958
rect 106096 235894 106148 235900
rect 106752 234394 106780 240037
rect 107396 237318 107424 240037
rect 108040 238754 108068 240037
rect 108672 239850 108700 240037
rect 109960 239850 109988 240037
rect 110604 239850 110632 240037
rect 107672 238726 108068 238754
rect 108592 239822 108700 239850
rect 109880 239822 109988 239850
rect 110420 239828 110472 239834
rect 107384 237312 107436 237318
rect 107384 237254 107436 237260
rect 106740 234388 106792 234394
rect 106740 234330 106792 234336
rect 106924 232552 106976 232558
rect 106924 232494 106976 232500
rect 106936 211886 106964 232494
rect 106924 211880 106976 211886
rect 106924 211822 106976 211828
rect 104900 209772 104952 209778
rect 104900 209714 104952 209720
rect 107672 205630 107700 238726
rect 108592 219434 108620 239822
rect 109880 231674 109908 239822
rect 110420 239770 110472 239776
rect 110524 239822 110632 239850
rect 111248 239834 111276 240037
rect 111892 239850 111920 240037
rect 111236 239828 111288 239834
rect 109868 231668 109920 231674
rect 109868 231610 109920 231616
rect 109880 219434 109908 231610
rect 107764 219406 108620 219434
rect 109696 219406 109908 219434
rect 107764 218006 107792 219406
rect 107752 218000 107804 218006
rect 107752 217942 107804 217948
rect 107660 205624 107712 205630
rect 107660 205566 107712 205572
rect 104164 199572 104216 199578
rect 104164 199514 104216 199520
rect 102140 198144 102192 198150
rect 102140 198086 102192 198092
rect 84200 188420 84252 188426
rect 84200 188362 84252 188368
rect 69018 186960 69074 186969
rect 69018 186895 69074 186904
rect 102048 185020 102100 185026
rect 102048 184962 102100 184968
rect 100668 184952 100720 184958
rect 100668 184894 100720 184900
rect 97816 178084 97868 178090
rect 97816 178026 97868 178032
rect 97828 176769 97856 178026
rect 100680 176769 100708 184894
rect 102060 177721 102088 184962
rect 107568 183592 107620 183598
rect 107568 183534 107620 183540
rect 105728 182436 105780 182442
rect 105728 182378 105780 182384
rect 105740 177721 105768 182378
rect 107580 177721 107608 183534
rect 102046 177712 102102 177721
rect 102046 177647 102102 177656
rect 105726 177712 105782 177721
rect 105726 177647 105782 177656
rect 107566 177712 107622 177721
rect 107566 177647 107622 177656
rect 109696 177342 109724 219406
rect 110432 187134 110460 239770
rect 110524 227730 110552 239822
rect 111236 239770 111288 239776
rect 111812 239822 111920 239850
rect 110512 227724 110564 227730
rect 110512 227666 110564 227672
rect 110524 226370 110552 227666
rect 110512 226364 110564 226370
rect 110512 226306 110564 226312
rect 111064 226364 111116 226370
rect 111064 226306 111116 226312
rect 111076 209098 111104 226306
rect 111064 209092 111116 209098
rect 111064 209034 111116 209040
rect 111812 193934 111840 239822
rect 112548 238814 112576 240037
rect 111892 238808 111944 238814
rect 111892 238750 111944 238756
rect 112536 238808 112588 238814
rect 112536 238750 112588 238756
rect 111904 229838 111932 238750
rect 111892 229832 111944 229838
rect 111892 229774 111944 229780
rect 113192 209710 113220 240037
rect 113836 235754 113864 240037
rect 114480 238814 114508 240037
rect 114560 239828 114612 239834
rect 114560 239770 114612 239776
rect 114468 238808 114520 238814
rect 114468 238750 114520 238756
rect 113824 235748 113876 235754
rect 113824 235690 113876 235696
rect 114572 216646 114600 239770
rect 115124 238542 115152 240037
rect 115756 239834 115784 240037
rect 115744 239828 115796 239834
rect 115744 239770 115796 239776
rect 116412 238754 116440 240037
rect 117056 239018 117084 240037
rect 117044 239012 117096 239018
rect 117044 238954 117096 238960
rect 115952 238726 116440 238754
rect 115112 238536 115164 238542
rect 115112 238478 115164 238484
rect 114560 216640 114612 216646
rect 114560 216582 114612 216588
rect 115952 210594 115980 238726
rect 117700 234734 117728 240037
rect 118344 238610 118372 240037
rect 118988 238754 119016 240037
rect 118804 238726 119016 238754
rect 118332 238604 118384 238610
rect 118332 238546 118384 238552
rect 118608 235612 118660 235618
rect 118608 235554 118660 235560
rect 118620 234734 118648 235554
rect 117688 234728 117740 234734
rect 117688 234670 117740 234676
rect 118608 234728 118660 234734
rect 118608 234670 118660 234676
rect 115940 210588 115992 210594
rect 115940 210530 115992 210536
rect 113180 209704 113232 209710
rect 113180 209646 113232 209652
rect 111800 193928 111852 193934
rect 111800 193870 111852 193876
rect 118620 191049 118648 234670
rect 118700 233912 118752 233918
rect 118700 233854 118752 233860
rect 118712 211818 118740 233854
rect 118804 229022 118832 238726
rect 119724 233918 119752 240094
rect 120000 238474 120028 240110
rect 120092 238882 120120 246298
rect 120080 238876 120132 238882
rect 120080 238818 120132 238824
rect 119988 238468 120040 238474
rect 119988 238410 120040 238416
rect 119712 233912 119764 233918
rect 119712 233854 119764 233860
rect 119344 229900 119396 229906
rect 119344 229842 119396 229848
rect 118792 229016 118844 229022
rect 118792 228958 118844 228964
rect 118700 211812 118752 211818
rect 118700 211754 118752 211760
rect 118606 191040 118662 191049
rect 118606 190975 118662 190984
rect 110420 187128 110472 187134
rect 110420 187070 110472 187076
rect 119356 185638 119384 229842
rect 120184 225622 120212 250951
rect 120172 225616 120224 225622
rect 120172 225558 120224 225564
rect 120736 199345 120764 269311
rect 120828 240106 120856 277471
rect 121460 277364 121512 277370
rect 121460 277306 121512 277312
rect 121472 276865 121500 277306
rect 121458 276856 121514 276865
rect 121458 276791 121514 276800
rect 121458 276176 121514 276185
rect 121458 276111 121514 276120
rect 121472 276078 121500 276111
rect 121460 276072 121512 276078
rect 121460 276014 121512 276020
rect 121550 275496 121606 275505
rect 121550 275431 121606 275440
rect 121564 274854 121592 275431
rect 121552 274848 121604 274854
rect 121458 274816 121514 274825
rect 121552 274790 121604 274796
rect 121458 274751 121460 274760
rect 121512 274751 121514 274760
rect 121460 274722 121512 274728
rect 122116 274718 122144 327830
rect 122208 324970 122236 331230
rect 122196 324964 122248 324970
rect 122196 324906 122248 324912
rect 122840 316736 122892 316742
rect 122840 316678 122892 316684
rect 122746 286376 122802 286385
rect 122852 286362 122880 316678
rect 123496 295322 123524 367066
rect 123576 362976 123628 362982
rect 123576 362918 123628 362924
rect 123484 295316 123536 295322
rect 123484 295258 123536 295264
rect 123588 295225 123616 362918
rect 123680 329798 123708 386582
rect 124140 384402 124168 487018
rect 124232 446486 124260 533326
rect 124508 530602 124536 582354
rect 125508 568540 125560 568546
rect 125508 568482 125560 568488
rect 125520 567866 125548 568482
rect 125508 567860 125560 567866
rect 125508 567802 125560 567808
rect 124864 536920 124916 536926
rect 124864 536862 124916 536868
rect 124496 530596 124548 530602
rect 124496 530538 124548 530544
rect 124310 495544 124366 495553
rect 124310 495479 124312 495488
rect 124364 495479 124366 495488
rect 124312 495450 124364 495456
rect 124312 494828 124364 494834
rect 124312 494770 124364 494776
rect 124220 446480 124272 446486
rect 124220 446422 124272 446428
rect 124220 438796 124272 438802
rect 124220 438738 124272 438744
rect 124128 384396 124180 384402
rect 124128 384338 124180 384344
rect 124128 378752 124180 378758
rect 124126 378720 124128 378729
rect 124180 378720 124182 378729
rect 124126 378655 124182 378664
rect 124232 332586 124260 438738
rect 124324 389978 124352 494770
rect 124404 446480 124456 446486
rect 124404 446422 124456 446428
rect 124416 438802 124444 446422
rect 124876 438870 124904 536862
rect 125612 533390 125640 635530
rect 125704 583710 125732 681702
rect 125784 674892 125836 674898
rect 125784 674834 125836 674840
rect 125692 583704 125744 583710
rect 125692 583646 125744 583652
rect 125796 578202 125824 674834
rect 196636 672042 196664 683130
rect 196624 672036 196676 672042
rect 196624 671978 196676 671984
rect 128452 669452 128504 669458
rect 128452 669394 128504 669400
rect 128360 637016 128412 637022
rect 128360 636958 128412 636964
rect 126980 635656 127032 635662
rect 126980 635598 127032 635604
rect 125968 586628 126020 586634
rect 125968 586570 126020 586576
rect 125876 580984 125928 580990
rect 125876 580926 125928 580932
rect 125784 578196 125836 578202
rect 125784 578138 125836 578144
rect 125692 538280 125744 538286
rect 125692 538222 125744 538228
rect 125600 533384 125652 533390
rect 125600 533326 125652 533332
rect 125600 484424 125652 484430
rect 125600 484366 125652 484372
rect 125508 439136 125560 439142
rect 125508 439078 125560 439084
rect 125520 438870 125548 439078
rect 124864 438864 124916 438870
rect 124864 438806 124916 438812
rect 125508 438864 125560 438870
rect 125508 438806 125560 438812
rect 124404 438796 124456 438802
rect 124404 438738 124456 438744
rect 124402 392592 124458 392601
rect 124402 392527 124458 392536
rect 124312 389972 124364 389978
rect 124312 389914 124364 389920
rect 124312 384804 124364 384810
rect 124312 384746 124364 384752
rect 124324 382974 124352 384746
rect 124312 382968 124364 382974
rect 124312 382910 124364 382916
rect 124416 336462 124444 392527
rect 125508 383104 125560 383110
rect 125508 383046 125560 383052
rect 125520 382702 125548 383046
rect 125508 382696 125560 382702
rect 125508 382638 125560 382644
rect 124956 365764 125008 365770
rect 124956 365706 125008 365712
rect 124864 356720 124916 356726
rect 124864 356662 124916 356668
rect 124876 339454 124904 356662
rect 124864 339448 124916 339454
rect 124864 339390 124916 339396
rect 124404 336456 124456 336462
rect 124404 336398 124456 336404
rect 124220 332580 124272 332586
rect 124220 332522 124272 332528
rect 124220 331220 124272 331226
rect 124220 331162 124272 331168
rect 123668 329792 123720 329798
rect 123668 329734 123720 329740
rect 123760 297016 123812 297022
rect 123760 296958 123812 296964
rect 123574 295216 123630 295225
rect 123574 295151 123630 295160
rect 123668 291304 123720 291310
rect 123668 291246 123720 291252
rect 123576 289196 123628 289202
rect 123576 289138 123628 289144
rect 123588 287054 123616 289138
rect 123680 289134 123708 291246
rect 123668 289128 123720 289134
rect 123668 289070 123720 289076
rect 123588 287026 123708 287054
rect 122802 286334 122880 286362
rect 122746 286311 122802 286320
rect 123576 283008 123628 283014
rect 123576 282950 123628 282956
rect 122194 282296 122250 282305
rect 122194 282231 122250 282240
rect 121552 274712 121604 274718
rect 121552 274654 121604 274660
rect 122104 274712 122156 274718
rect 122104 274654 122156 274660
rect 121564 274145 121592 274654
rect 121550 274136 121606 274145
rect 121550 274071 121606 274080
rect 121458 273456 121514 273465
rect 121458 273391 121514 273400
rect 121472 273358 121500 273391
rect 121460 273352 121512 273358
rect 121460 273294 121512 273300
rect 121460 273216 121512 273222
rect 121460 273158 121512 273164
rect 121472 272785 121500 273158
rect 121458 272776 121514 272785
rect 121458 272711 121514 272720
rect 121458 271416 121514 271425
rect 121458 271351 121514 271360
rect 121472 270570 121500 271351
rect 121460 270564 121512 270570
rect 121460 270506 121512 270512
rect 121550 270056 121606 270065
rect 121550 269991 121606 270000
rect 121564 269142 121592 269991
rect 121552 269136 121604 269142
rect 121552 269078 121604 269084
rect 121460 269068 121512 269074
rect 121460 269010 121512 269016
rect 121472 268705 121500 269010
rect 121458 268696 121514 268705
rect 121458 268631 121514 268640
rect 121458 268016 121514 268025
rect 121458 267951 121514 267960
rect 121472 267782 121500 267951
rect 121460 267776 121512 267782
rect 121460 267718 121512 267724
rect 121550 267336 121606 267345
rect 121550 267271 121606 267280
rect 121458 266656 121514 266665
rect 121458 266591 121514 266600
rect 121472 266490 121500 266591
rect 121460 266484 121512 266490
rect 121460 266426 121512 266432
rect 121564 266422 121592 267271
rect 121552 266416 121604 266422
rect 121552 266358 121604 266364
rect 121550 265976 121606 265985
rect 121550 265911 121606 265920
rect 121458 265296 121514 265305
rect 121458 265231 121514 265240
rect 121472 265062 121500 265231
rect 121460 265056 121512 265062
rect 121460 264998 121512 265004
rect 121564 264994 121592 265911
rect 121552 264988 121604 264994
rect 121552 264930 121604 264936
rect 121550 263936 121606 263945
rect 121550 263871 121606 263880
rect 121564 263634 121592 263871
rect 121552 263628 121604 263634
rect 121552 263570 121604 263576
rect 121460 263560 121512 263566
rect 121460 263502 121512 263508
rect 121472 263265 121500 263502
rect 121458 263256 121514 263265
rect 121458 263191 121514 263200
rect 121460 262812 121512 262818
rect 121460 262754 121512 262760
rect 121472 262585 121500 262754
rect 121458 262576 121514 262585
rect 121458 262511 121514 262520
rect 121552 262200 121604 262206
rect 121552 262142 121604 262148
rect 121460 261928 121512 261934
rect 121458 261896 121460 261905
rect 121512 261896 121514 261905
rect 121458 261831 121514 261840
rect 121564 261225 121592 262142
rect 121550 261216 121606 261225
rect 121550 261151 121606 261160
rect 121460 260840 121512 260846
rect 121460 260782 121512 260788
rect 121472 260545 121500 260782
rect 121458 260536 121514 260545
rect 121458 260471 121514 260480
rect 121458 259856 121514 259865
rect 121458 259791 121514 259800
rect 121472 259486 121500 259791
rect 121460 259480 121512 259486
rect 121460 259422 121512 259428
rect 121552 259412 121604 259418
rect 121552 259354 121604 259360
rect 121564 258505 121592 259354
rect 121642 259176 121698 259185
rect 121642 259111 121698 259120
rect 121550 258496 121606 258505
rect 121550 258431 121606 258440
rect 121656 258126 121684 259111
rect 121644 258120 121696 258126
rect 121644 258062 121696 258068
rect 121460 258052 121512 258058
rect 121460 257994 121512 258000
rect 121472 257145 121500 257994
rect 121550 257816 121606 257825
rect 121550 257751 121606 257760
rect 121458 257136 121514 257145
rect 121458 257071 121514 257080
rect 121564 256766 121592 257751
rect 121552 256760 121604 256766
rect 121552 256702 121604 256708
rect 121460 256692 121512 256698
rect 121460 256634 121512 256640
rect 121472 256465 121500 256634
rect 121552 256624 121604 256630
rect 121552 256566 121604 256572
rect 121458 256456 121514 256465
rect 121458 256391 121514 256400
rect 121564 255785 121592 256566
rect 121550 255776 121606 255785
rect 121550 255711 121606 255720
rect 121458 255096 121514 255105
rect 121458 255031 121514 255040
rect 121472 253978 121500 255031
rect 122102 254416 122158 254425
rect 122102 254351 122158 254360
rect 121460 253972 121512 253978
rect 121460 253914 121512 253920
rect 121458 253736 121514 253745
rect 121458 253671 121514 253680
rect 121472 252686 121500 253671
rect 121550 253056 121606 253065
rect 121550 252991 121606 253000
rect 121460 252680 121512 252686
rect 121460 252622 121512 252628
rect 121564 252618 121592 252991
rect 121552 252612 121604 252618
rect 121552 252554 121604 252560
rect 121460 252544 121512 252550
rect 121460 252486 121512 252492
rect 121472 252385 121500 252486
rect 121458 252376 121514 252385
rect 121458 252311 121514 252320
rect 121458 251696 121514 251705
rect 121458 251631 121514 251640
rect 121472 251258 121500 251631
rect 121460 251252 121512 251258
rect 121460 251194 121512 251200
rect 121458 250336 121514 250345
rect 121458 250271 121514 250280
rect 121472 249830 121500 250271
rect 121460 249824 121512 249830
rect 121460 249766 121512 249772
rect 121552 249756 121604 249762
rect 121552 249698 121604 249704
rect 121564 248985 121592 249698
rect 121550 248976 121606 248985
rect 121550 248911 121606 248920
rect 121552 248396 121604 248402
rect 121552 248338 121604 248344
rect 121458 248296 121514 248305
rect 121458 248231 121514 248240
rect 121472 247994 121500 248231
rect 121460 247988 121512 247994
rect 121460 247930 121512 247936
rect 121564 247625 121592 248338
rect 121550 247616 121606 247625
rect 121550 247551 121606 247560
rect 121550 246936 121606 246945
rect 121550 246871 121606 246880
rect 121458 246256 121514 246265
rect 121458 246191 121514 246200
rect 121472 245682 121500 246191
rect 121564 245818 121592 246871
rect 121552 245812 121604 245818
rect 121552 245754 121604 245760
rect 121460 245676 121512 245682
rect 121460 245618 121512 245624
rect 121552 245608 121604 245614
rect 121458 245576 121514 245585
rect 121552 245550 121604 245556
rect 121458 245511 121514 245520
rect 121472 244322 121500 245511
rect 121564 244905 121592 245550
rect 121550 244896 121606 244905
rect 121550 244831 121606 244840
rect 121460 244316 121512 244322
rect 121460 244258 121512 244264
rect 121458 244216 121514 244225
rect 121458 244151 121514 244160
rect 121472 242962 121500 244151
rect 121460 242956 121512 242962
rect 121460 242898 121512 242904
rect 121552 242888 121604 242894
rect 121458 242856 121514 242865
rect 121552 242830 121604 242836
rect 121458 242791 121460 242800
rect 121512 242791 121514 242800
rect 121460 242762 121512 242768
rect 121564 242185 121592 242830
rect 121550 242176 121606 242185
rect 121550 242111 121606 242120
rect 121458 240816 121514 240825
rect 121458 240751 121514 240760
rect 121472 240242 121500 240751
rect 121460 240236 121512 240242
rect 121460 240178 121512 240184
rect 121458 240136 121514 240145
rect 120816 240100 120868 240106
rect 121458 240071 121514 240080
rect 120816 240042 120868 240048
rect 121472 238882 121500 240071
rect 121460 238876 121512 238882
rect 121460 238818 121512 238824
rect 122116 222970 122144 254351
rect 122208 247722 122236 282231
rect 123484 273284 123536 273290
rect 123484 273226 123536 273232
rect 122286 272096 122342 272105
rect 122286 272031 122342 272040
rect 122300 247790 122328 272031
rect 123496 261934 123524 273226
rect 123484 261928 123536 261934
rect 123484 261870 123536 261876
rect 123484 247988 123536 247994
rect 123484 247930 123536 247936
rect 122288 247784 122340 247790
rect 122288 247726 122340 247732
rect 122196 247716 122248 247722
rect 122196 247658 122248 247664
rect 122104 222964 122156 222970
rect 122104 222906 122156 222912
rect 120722 199336 120778 199345
rect 120722 199271 120778 199280
rect 119344 185632 119396 185638
rect 119344 185574 119396 185580
rect 119712 182368 119764 182374
rect 119712 182310 119764 182316
rect 110696 182300 110748 182306
rect 110696 182242 110748 182248
rect 109960 179444 110012 179450
rect 109960 179386 110012 179392
rect 109684 177336 109736 177342
rect 109684 177278 109736 177284
rect 109972 177041 110000 179386
rect 110708 177721 110736 182242
rect 116952 180872 117004 180878
rect 116952 180814 117004 180820
rect 115848 179512 115900 179518
rect 115848 179454 115900 179460
rect 114376 178220 114428 178226
rect 114376 178162 114428 178168
rect 112260 178152 112312 178158
rect 112260 178094 112312 178100
rect 110694 177712 110750 177721
rect 110694 177647 110750 177656
rect 109958 177032 110014 177041
rect 109958 176967 110014 176976
rect 108120 176860 108172 176866
rect 108120 176802 108172 176808
rect 108132 176769 108160 176802
rect 112272 176769 112300 178094
rect 114388 176769 114416 178162
rect 115860 177177 115888 179454
rect 116964 177721 116992 180814
rect 119724 177721 119752 182310
rect 123300 182232 123352 182238
rect 123300 182174 123352 182180
rect 121184 180940 121236 180946
rect 121184 180882 121236 180888
rect 121196 177721 121224 180882
rect 123312 177721 123340 182174
rect 123496 178770 123524 247930
rect 123588 234462 123616 282950
rect 123680 238950 123708 287026
rect 123772 279478 123800 296958
rect 124128 292664 124180 292670
rect 124128 292606 124180 292612
rect 124140 292534 124168 292606
rect 124128 292528 124180 292534
rect 124128 292470 124180 292476
rect 123760 279472 123812 279478
rect 123760 279414 123812 279420
rect 124140 264246 124168 292470
rect 124232 287026 124260 331162
rect 124312 329792 124364 329798
rect 124312 329734 124364 329740
rect 124324 328506 124352 329734
rect 124312 328500 124364 328506
rect 124312 328442 124364 328448
rect 124324 322454 124352 328442
rect 124312 322448 124364 322454
rect 124312 322390 124364 322396
rect 124310 314664 124366 314673
rect 124310 314599 124312 314608
rect 124364 314599 124366 314608
rect 124312 314570 124364 314576
rect 124864 295384 124916 295390
rect 124864 295326 124916 295332
rect 124220 287020 124272 287026
rect 124220 286962 124272 286968
rect 124128 264240 124180 264246
rect 124128 264182 124180 264188
rect 123760 245812 123812 245818
rect 123760 245754 123812 245760
rect 123668 238944 123720 238950
rect 123668 238886 123720 238892
rect 123576 234456 123628 234462
rect 123576 234398 123628 234404
rect 123772 202366 123800 245754
rect 123760 202360 123812 202366
rect 123760 202302 123812 202308
rect 124876 187066 124904 295326
rect 124968 294982 124996 365706
rect 125520 358766 125548 382638
rect 125612 381546 125640 484366
rect 125704 436082 125732 538222
rect 125784 535492 125836 535498
rect 125784 535434 125836 535440
rect 125796 438734 125824 535434
rect 125888 487082 125916 580926
rect 125980 535537 126008 586570
rect 126244 575544 126296 575550
rect 126244 575486 126296 575492
rect 126256 565146 126284 575486
rect 126244 565140 126296 565146
rect 126244 565082 126296 565088
rect 125966 535528 126022 535537
rect 125966 535463 126022 535472
rect 126992 535430 127020 635598
rect 127164 634092 127216 634098
rect 127164 634034 127216 634040
rect 127070 583808 127126 583817
rect 127070 583743 127126 583752
rect 126980 535424 127032 535430
rect 126980 535366 127032 535372
rect 126992 534138 127020 535366
rect 126980 534132 127032 534138
rect 126980 534074 127032 534080
rect 127084 491298 127112 583743
rect 127176 540938 127204 634034
rect 127254 589928 127310 589937
rect 127254 589863 127310 589872
rect 127164 540932 127216 540938
rect 127164 540874 127216 540880
rect 127164 534744 127216 534750
rect 127164 534686 127216 534692
rect 127072 491292 127124 491298
rect 127072 491234 127124 491240
rect 126980 488572 127032 488578
rect 126980 488514 127032 488520
rect 125876 487076 125928 487082
rect 125876 487018 125928 487024
rect 125876 447160 125928 447166
rect 125876 447102 125928 447108
rect 125784 438728 125836 438734
rect 125784 438670 125836 438676
rect 125692 436076 125744 436082
rect 125692 436018 125744 436024
rect 125600 381540 125652 381546
rect 125600 381482 125652 381488
rect 125508 358760 125560 358766
rect 125508 358702 125560 358708
rect 125796 336598 125824 438670
rect 125888 369238 125916 447102
rect 126888 383172 126940 383178
rect 126888 383114 126940 383120
rect 126900 381614 126928 383114
rect 126992 382702 127020 488514
rect 127176 437442 127204 534686
rect 127268 533458 127296 589863
rect 128372 538218 128400 636958
rect 128464 571334 128492 669394
rect 133972 669384 134024 669390
rect 133972 669326 134024 669332
rect 128544 663876 128596 663882
rect 128544 663818 128596 663824
rect 128452 571328 128504 571334
rect 128452 571270 128504 571276
rect 128556 566506 128584 663818
rect 133788 657552 133840 657558
rect 133788 657494 133840 657500
rect 133800 656946 133828 657494
rect 132500 656940 132552 656946
rect 132500 656882 132552 656888
rect 133788 656940 133840 656946
rect 133788 656882 133840 656888
rect 129832 651432 129884 651438
rect 129832 651374 129884 651380
rect 129740 632800 129792 632806
rect 129740 632742 129792 632748
rect 128636 583840 128688 583846
rect 128636 583782 128688 583788
rect 128544 566500 128596 566506
rect 128544 566442 128596 566448
rect 128360 538212 128412 538218
rect 128360 538154 128412 538160
rect 128452 536104 128504 536110
rect 128452 536046 128504 536052
rect 127256 533452 127308 533458
rect 127256 533394 127308 533400
rect 128360 495508 128412 495514
rect 128360 495450 128412 495456
rect 127348 493332 127400 493338
rect 127348 493274 127400 493280
rect 127164 437436 127216 437442
rect 127164 437378 127216 437384
rect 127256 396840 127308 396846
rect 127256 396782 127308 396788
rect 127072 386504 127124 386510
rect 127072 386446 127124 386452
rect 126980 382696 127032 382702
rect 126980 382638 127032 382644
rect 126244 381608 126296 381614
rect 126244 381550 126296 381556
rect 126888 381608 126940 381614
rect 126888 381550 126940 381556
rect 125876 369232 125928 369238
rect 125876 369174 125928 369180
rect 125784 336592 125836 336598
rect 125784 336534 125836 336540
rect 125508 314628 125560 314634
rect 125508 314570 125560 314576
rect 125520 313410 125548 314570
rect 125508 313404 125560 313410
rect 125508 313346 125560 313352
rect 126256 301034 126284 381550
rect 126428 367804 126480 367810
rect 126428 367746 126480 367752
rect 126336 367192 126388 367198
rect 126336 367134 126388 367140
rect 125784 301028 125836 301034
rect 125784 300970 125836 300976
rect 126244 301028 126296 301034
rect 126244 300970 126296 300976
rect 125796 300218 125824 300970
rect 125784 300212 125836 300218
rect 125784 300154 125836 300160
rect 125048 295588 125100 295594
rect 125048 295530 125100 295536
rect 124956 294976 125008 294982
rect 124956 294918 125008 294924
rect 124956 282192 125008 282198
rect 124956 282134 125008 282140
rect 124968 235686 124996 282134
rect 125060 268394 125088 295530
rect 126348 294846 126376 367134
rect 126440 352578 126468 367746
rect 126428 352572 126480 352578
rect 126428 352514 126480 352520
rect 126888 336592 126940 336598
rect 126888 336534 126940 336540
rect 126900 336054 126928 336534
rect 126888 336048 126940 336054
rect 126888 335990 126940 335996
rect 126428 334756 126480 334762
rect 126428 334698 126480 334704
rect 126336 294840 126388 294846
rect 126336 294782 126388 294788
rect 125598 293312 125654 293321
rect 125598 293247 125654 293256
rect 125140 271924 125192 271930
rect 125140 271866 125192 271872
rect 125048 268388 125100 268394
rect 125048 268330 125100 268336
rect 125152 262818 125180 271866
rect 125140 262812 125192 262818
rect 125140 262754 125192 262760
rect 125612 239018 125640 293247
rect 126242 293176 126298 293185
rect 126242 293111 126298 293120
rect 125600 239012 125652 239018
rect 125600 238954 125652 238960
rect 124956 235680 125008 235686
rect 124956 235622 125008 235628
rect 126256 196790 126284 293111
rect 126440 289202 126468 334698
rect 126980 332580 127032 332586
rect 126980 332522 127032 332528
rect 126888 322924 126940 322930
rect 126888 322866 126940 322872
rect 126428 289196 126480 289202
rect 126428 289138 126480 289144
rect 126900 262206 126928 322866
rect 126888 262200 126940 262206
rect 126888 262142 126940 262148
rect 126900 261526 126928 262142
rect 126888 261520 126940 261526
rect 126888 261462 126940 261468
rect 126336 252680 126388 252686
rect 126336 252622 126388 252628
rect 126348 200938 126376 252622
rect 126428 240236 126480 240242
rect 126428 240178 126480 240184
rect 126440 224330 126468 240178
rect 126992 230450 127020 332522
rect 127084 283626 127112 386446
rect 127164 384396 127216 384402
rect 127164 384338 127216 384344
rect 127176 300150 127204 384338
rect 127268 336666 127296 396782
rect 127360 393990 127388 493274
rect 127348 393984 127400 393990
rect 127348 393926 127400 393932
rect 128372 389842 128400 495450
rect 128464 439074 128492 536046
rect 128556 474638 128584 566442
rect 128648 496126 128676 583782
rect 129752 534750 129780 632742
rect 129844 554742 129872 651374
rect 129924 638988 129976 638994
rect 129924 638930 129976 638936
rect 129832 554736 129884 554742
rect 129832 554678 129884 554684
rect 129844 554130 129872 554678
rect 129832 554124 129884 554130
rect 129832 554066 129884 554072
rect 129936 543726 129964 638930
rect 131120 638308 131172 638314
rect 131120 638250 131172 638256
rect 130106 585440 130162 585449
rect 130106 585375 130162 585384
rect 130016 552084 130068 552090
rect 130016 552026 130068 552032
rect 129924 543720 129976 543726
rect 129924 543662 129976 543668
rect 129740 534744 129792 534750
rect 129740 534686 129792 534692
rect 128636 496120 128688 496126
rect 128636 496062 128688 496068
rect 129924 493400 129976 493406
rect 129924 493342 129976 493348
rect 129832 492720 129884 492726
rect 129832 492662 129884 492668
rect 128544 474632 128596 474638
rect 128544 474574 128596 474580
rect 128544 467152 128596 467158
rect 128544 467094 128596 467100
rect 128452 439068 128504 439074
rect 128452 439010 128504 439016
rect 128452 436144 128504 436150
rect 128452 436086 128504 436092
rect 128360 389836 128412 389842
rect 128360 389778 128412 389784
rect 128372 389230 128400 389778
rect 128360 389224 128412 389230
rect 128360 389166 128412 389172
rect 128360 385688 128412 385694
rect 128360 385630 128412 385636
rect 128372 385082 128400 385630
rect 128360 385076 128412 385082
rect 128360 385018 128412 385024
rect 127256 336660 127308 336666
rect 127256 336602 127308 336608
rect 127164 300144 127216 300150
rect 127164 300086 127216 300092
rect 127622 297392 127678 297401
rect 127622 297327 127678 297336
rect 127072 283620 127124 283626
rect 127072 283562 127124 283568
rect 127084 283014 127112 283562
rect 127072 283008 127124 283014
rect 127072 282950 127124 282956
rect 126980 230444 127032 230450
rect 126980 230386 127032 230392
rect 126428 224324 126480 224330
rect 126428 224266 126480 224272
rect 126336 200932 126388 200938
rect 126336 200874 126388 200880
rect 127636 198014 127664 297327
rect 127716 282940 127768 282946
rect 127716 282882 127768 282888
rect 127728 271182 127756 282882
rect 128268 274848 128320 274854
rect 128268 274790 128320 274796
rect 127716 271176 127768 271182
rect 127716 271118 127768 271124
rect 128280 237386 128308 274790
rect 128268 237380 128320 237386
rect 128268 237322 128320 237328
rect 128372 237250 128400 385018
rect 128464 339386 128492 436086
rect 128556 396778 128584 467094
rect 129740 444440 129792 444446
rect 129740 444382 129792 444388
rect 128544 396772 128596 396778
rect 128544 396714 128596 396720
rect 128544 389972 128596 389978
rect 128544 389914 128596 389920
rect 128452 339380 128504 339386
rect 128452 339322 128504 339328
rect 128556 325038 128584 389914
rect 128636 358760 128688 358766
rect 128636 358702 128688 358708
rect 128648 357474 128676 358702
rect 128636 357468 128688 357474
rect 128636 357410 128688 357416
rect 128648 330818 128676 357410
rect 128728 342916 128780 342922
rect 128728 342858 128780 342864
rect 128740 342281 128768 342858
rect 128726 342272 128782 342281
rect 128726 342207 128782 342216
rect 129752 337385 129780 444382
rect 129844 397202 129872 492662
rect 129936 402914 129964 493342
rect 130028 460222 130056 552026
rect 130120 494766 130148 585375
rect 130200 552696 130252 552702
rect 130200 552638 130252 552644
rect 130212 552090 130240 552638
rect 130200 552084 130252 552090
rect 130200 552026 130252 552032
rect 130752 543720 130804 543726
rect 130752 543662 130804 543668
rect 130764 543046 130792 543662
rect 130752 543040 130804 543046
rect 130752 542982 130804 542988
rect 131132 538150 131160 638250
rect 131304 632732 131356 632738
rect 131304 632674 131356 632680
rect 131210 585168 131266 585177
rect 131210 585103 131266 585112
rect 131120 538144 131172 538150
rect 131120 538086 131172 538092
rect 131132 535430 131160 538086
rect 130384 535424 130436 535430
rect 130384 535366 130436 535372
rect 131120 535424 131172 535430
rect 131120 535366 131172 535372
rect 130108 494760 130160 494766
rect 130108 494702 130160 494708
rect 130016 460216 130068 460222
rect 130016 460158 130068 460164
rect 130396 442270 130424 535366
rect 131120 534132 131172 534138
rect 131120 534074 131172 534080
rect 130384 442264 130436 442270
rect 130384 442206 130436 442212
rect 131132 439006 131160 534074
rect 131224 492250 131252 585103
rect 131316 559638 131344 632674
rect 131764 629944 131816 629950
rect 131764 629886 131816 629892
rect 131304 559632 131356 559638
rect 131304 559574 131356 559580
rect 131304 540932 131356 540938
rect 131304 540874 131356 540880
rect 131212 492244 131264 492250
rect 131212 492186 131264 492192
rect 131120 439000 131172 439006
rect 131120 438942 131172 438948
rect 129936 402886 130240 402914
rect 129844 397174 130148 397202
rect 129832 396908 129884 396914
rect 129832 396850 129884 396856
rect 129844 396166 129872 396850
rect 129832 396160 129884 396166
rect 129832 396102 129884 396108
rect 130016 396160 130068 396166
rect 130016 396102 130068 396108
rect 129922 378720 129978 378729
rect 129922 378655 129978 378664
rect 129832 378208 129884 378214
rect 129832 378150 129884 378156
rect 129844 374678 129872 378150
rect 129832 374672 129884 374678
rect 129832 374614 129884 374620
rect 129832 370524 129884 370530
rect 129832 370466 129884 370472
rect 129738 337376 129794 337385
rect 129738 337311 129794 337320
rect 129752 334626 129780 337311
rect 129740 334620 129792 334626
rect 129740 334562 129792 334568
rect 128636 330812 128688 330818
rect 128636 330754 128688 330760
rect 129740 330744 129792 330750
rect 129740 330686 129792 330692
rect 129752 329866 129780 330686
rect 129740 329860 129792 329866
rect 129740 329802 129792 329808
rect 128544 325032 128596 325038
rect 128544 324974 128596 324980
rect 129188 313336 129240 313342
rect 129188 313278 129240 313284
rect 129004 307080 129056 307086
rect 129004 307022 129056 307028
rect 128360 237244 128412 237250
rect 128360 237186 128412 237192
rect 127624 198008 127676 198014
rect 127624 197950 127676 197956
rect 126244 196784 126296 196790
rect 126244 196726 126296 196732
rect 129016 193866 129044 307022
rect 129096 304360 129148 304366
rect 129096 304302 129148 304308
rect 129108 195566 129136 304302
rect 129200 249762 129228 313278
rect 129188 249756 129240 249762
rect 129188 249698 129240 249704
rect 129752 235618 129780 329802
rect 129844 292534 129872 370466
rect 129936 318073 129964 378655
rect 130028 340814 130056 396102
rect 130120 394126 130148 397174
rect 130212 395350 130240 402886
rect 130200 395344 130252 395350
rect 130200 395286 130252 395292
rect 130108 394120 130160 394126
rect 130108 394062 130160 394068
rect 131224 392698 131252 492186
rect 131316 447166 131344 540874
rect 131776 539510 131804 629886
rect 132512 559570 132540 656882
rect 132868 644564 132920 644570
rect 132868 644506 132920 644512
rect 132684 634160 132736 634166
rect 132684 634102 132736 634108
rect 132592 567860 132644 567866
rect 132592 567802 132644 567808
rect 132500 559564 132552 559570
rect 132500 559506 132552 559512
rect 131764 539504 131816 539510
rect 131764 539446 131816 539452
rect 132500 496120 132552 496126
rect 132500 496062 132552 496068
rect 131304 447160 131356 447166
rect 131304 447102 131356 447108
rect 131488 439068 131540 439074
rect 131488 439010 131540 439016
rect 131304 405068 131356 405074
rect 131304 405010 131356 405016
rect 131212 392692 131264 392698
rect 131212 392634 131264 392640
rect 130384 389224 130436 389230
rect 130384 389166 130436 389172
rect 130396 378826 130424 389166
rect 130384 378820 130436 378826
rect 130384 378762 130436 378768
rect 131316 341630 131344 405010
rect 131396 394052 131448 394058
rect 131396 393994 131448 394000
rect 131408 393446 131436 393994
rect 131396 393440 131448 393446
rect 131396 393382 131448 393388
rect 131304 341624 131356 341630
rect 131304 341566 131356 341572
rect 130016 340808 130068 340814
rect 130016 340750 130068 340756
rect 131212 337408 131264 337414
rect 131212 337350 131264 337356
rect 131120 322312 131172 322318
rect 131120 322254 131172 322260
rect 131132 321638 131160 322254
rect 131120 321632 131172 321638
rect 131120 321574 131172 321580
rect 129922 318064 129978 318073
rect 129922 317999 129978 318008
rect 129924 317416 129976 317422
rect 129922 317384 129924 317393
rect 129976 317384 129978 317393
rect 129922 317319 129978 317328
rect 130384 316736 130436 316742
rect 130384 316678 130436 316684
rect 130290 316160 130346 316169
rect 130290 316095 130346 316104
rect 130304 316062 130332 316095
rect 130292 316056 130344 316062
rect 130292 315998 130344 316004
rect 129924 298784 129976 298790
rect 129924 298726 129976 298732
rect 129832 292528 129884 292534
rect 129832 292470 129884 292476
rect 129936 274854 129964 298726
rect 130396 280158 130424 316678
rect 130474 292088 130530 292097
rect 130474 292023 130530 292032
rect 130384 280152 130436 280158
rect 130384 280094 130436 280100
rect 129924 274848 129976 274854
rect 129924 274790 129976 274796
rect 130384 269136 130436 269142
rect 130384 269078 130436 269084
rect 129740 235612 129792 235618
rect 129740 235554 129792 235560
rect 129096 195560 129148 195566
rect 129096 195502 129148 195508
rect 129004 193860 129056 193866
rect 129004 193802 129056 193808
rect 130396 192642 130424 269078
rect 130488 215937 130516 292023
rect 131132 277370 131160 321574
rect 131120 277364 131172 277370
rect 131120 277306 131172 277312
rect 130568 276072 130620 276078
rect 130568 276014 130620 276020
rect 130580 240038 130608 276014
rect 130568 240032 130620 240038
rect 130568 239974 130620 239980
rect 131224 238814 131252 337350
rect 131408 333946 131436 393382
rect 131500 334762 131528 439010
rect 132512 385014 132540 496062
rect 132604 475386 132632 567802
rect 132696 539442 132724 634102
rect 132776 559564 132828 559570
rect 132776 559506 132828 559512
rect 132684 539436 132736 539442
rect 132684 539378 132736 539384
rect 132592 475380 132644 475386
rect 132592 475322 132644 475328
rect 132500 385008 132552 385014
rect 132500 384950 132552 384956
rect 132604 383654 132632 475322
rect 132788 467838 132816 559506
rect 132880 549234 132908 644506
rect 133880 635520 133932 635526
rect 133880 635462 133932 635468
rect 133892 634846 133920 635462
rect 133880 634840 133932 634846
rect 133880 634782 133932 634788
rect 132868 549228 132920 549234
rect 132868 549170 132920 549176
rect 133788 549228 133840 549234
rect 133788 549170 133840 549176
rect 133800 548622 133828 549170
rect 133788 548616 133840 548622
rect 133788 548558 133840 548564
rect 132868 539640 132920 539646
rect 132868 539582 132920 539588
rect 132776 467832 132828 467838
rect 132776 467774 132828 467780
rect 132880 442377 132908 539582
rect 133892 535362 133920 634782
rect 133984 572014 134012 669326
rect 142160 663808 142212 663814
rect 142160 663750 142212 663756
rect 136732 659796 136784 659802
rect 136732 659738 136784 659744
rect 135260 644496 135312 644502
rect 135260 644438 135312 644444
rect 134064 643748 134116 643754
rect 134064 643690 134116 643696
rect 135168 643748 135220 643754
rect 135168 643690 135220 643696
rect 133972 572008 134024 572014
rect 133972 571950 134024 571956
rect 134076 557534 134104 643690
rect 135180 643142 135208 643690
rect 135168 643136 135220 643142
rect 135168 643078 135220 643084
rect 134156 572008 134208 572014
rect 134156 571950 134208 571956
rect 133984 557506 134104 557534
rect 133984 554062 134012 557506
rect 133972 554056 134024 554062
rect 133972 553998 134024 554004
rect 133880 535356 133932 535362
rect 133880 535298 133932 535304
rect 133880 472048 133932 472054
rect 133880 471990 133932 471996
rect 132866 442368 132922 442377
rect 132866 442303 132922 442312
rect 132684 439136 132736 439142
rect 132684 439078 132736 439084
rect 132512 383626 132632 383654
rect 132512 369850 132540 383626
rect 132592 375420 132644 375426
rect 132592 375362 132644 375368
rect 132500 369844 132552 369850
rect 132500 369786 132552 369792
rect 132604 354674 132632 375362
rect 132512 354646 132632 354674
rect 131762 342272 131818 342281
rect 131762 342207 131818 342216
rect 131488 334756 131540 334762
rect 131488 334698 131540 334704
rect 131396 333940 131448 333946
rect 131396 333882 131448 333888
rect 131776 257378 131804 342207
rect 132512 326534 132540 354646
rect 132590 347712 132646 347721
rect 132590 347647 132646 347656
rect 132604 347070 132632 347647
rect 132592 347064 132644 347070
rect 132592 347006 132644 347012
rect 132696 337890 132724 439078
rect 133144 390720 133196 390726
rect 133144 390662 133196 390668
rect 133156 360330 133184 390662
rect 133788 376032 133840 376038
rect 133788 375974 133840 375980
rect 133800 375426 133828 375974
rect 133788 375420 133840 375426
rect 133788 375362 133840 375368
rect 133892 365702 133920 471990
rect 133984 462330 134012 553998
rect 134064 494760 134116 494766
rect 134064 494702 134116 494708
rect 133972 462324 134024 462330
rect 133972 462266 134024 462272
rect 133972 440292 134024 440298
rect 133972 440234 134024 440240
rect 133880 365696 133932 365702
rect 133880 365638 133932 365644
rect 133144 360324 133196 360330
rect 133144 360266 133196 360272
rect 132776 350600 132828 350606
rect 132776 350542 132828 350548
rect 132684 337884 132736 337890
rect 132684 337826 132736 337832
rect 132500 326528 132552 326534
rect 132500 326470 132552 326476
rect 132498 320240 132554 320249
rect 132498 320175 132554 320184
rect 131856 274780 131908 274786
rect 131856 274722 131908 274728
rect 131764 257372 131816 257378
rect 131764 257314 131816 257320
rect 131212 238808 131264 238814
rect 131212 238750 131264 238756
rect 131776 235754 131804 257314
rect 131764 235748 131816 235754
rect 131764 235690 131816 235696
rect 131868 217598 131896 274722
rect 132512 237318 132540 320175
rect 132592 301504 132644 301510
rect 132592 301446 132644 301452
rect 132604 242826 132632 301446
rect 132788 300830 132816 350542
rect 133156 315314 133184 360266
rect 133880 354068 133932 354074
rect 133880 354010 133932 354016
rect 133892 353433 133920 354010
rect 133878 353424 133934 353433
rect 133878 353359 133934 353368
rect 133788 347064 133840 347070
rect 133788 347006 133840 347012
rect 133800 346526 133828 347006
rect 133788 346520 133840 346526
rect 133788 346462 133840 346468
rect 133880 337476 133932 337482
rect 133880 337418 133932 337424
rect 133144 315308 133196 315314
rect 133144 315250 133196 315256
rect 133144 308576 133196 308582
rect 133144 308518 133196 308524
rect 132776 300824 132828 300830
rect 132776 300766 132828 300772
rect 132592 242820 132644 242826
rect 132592 242762 132644 242768
rect 132500 237312 132552 237318
rect 132500 237254 132552 237260
rect 131856 217592 131908 217598
rect 131856 217534 131908 217540
rect 130474 215928 130530 215937
rect 130474 215863 130530 215872
rect 130384 192636 130436 192642
rect 130384 192578 130436 192584
rect 133156 190126 133184 308518
rect 133788 300824 133840 300830
rect 133788 300766 133840 300772
rect 133800 300218 133828 300766
rect 133788 300212 133840 300218
rect 133788 300154 133840 300160
rect 133236 295656 133288 295662
rect 133236 295598 133288 295604
rect 133248 209302 133276 295598
rect 133892 273222 133920 337418
rect 133984 336734 134012 440234
rect 134076 391270 134104 494702
rect 134168 480214 134196 571950
rect 135168 566500 135220 566506
rect 135168 566442 135220 566448
rect 135180 565894 135208 566442
rect 134524 565888 134576 565894
rect 134524 565830 134576 565836
rect 135168 565888 135220 565894
rect 135168 565830 135220 565836
rect 134156 480208 134208 480214
rect 134156 480150 134208 480156
rect 134168 478922 134196 480150
rect 134156 478916 134208 478922
rect 134156 478858 134208 478864
rect 134536 474706 134564 565830
rect 135272 547194 135300 644438
rect 136640 636880 136692 636886
rect 136640 636822 136692 636828
rect 135904 561672 135956 561678
rect 135904 561614 135956 561620
rect 135916 560998 135944 561614
rect 135904 560992 135956 560998
rect 135904 560934 135956 560940
rect 135260 547188 135312 547194
rect 135260 547130 135312 547136
rect 134524 474700 134576 474706
rect 134524 474642 134576 474648
rect 135272 458930 135300 547130
rect 135444 474700 135496 474706
rect 135444 474642 135496 474648
rect 135260 458924 135312 458930
rect 135260 458866 135312 458872
rect 135272 458250 135300 458866
rect 135260 458244 135312 458250
rect 135260 458186 135312 458192
rect 135352 445800 135404 445806
rect 135352 445742 135404 445748
rect 135260 392216 135312 392222
rect 135260 392158 135312 392164
rect 134064 391264 134116 391270
rect 134064 391206 134116 391212
rect 134064 390652 134116 390658
rect 134064 390594 134116 390600
rect 133972 336728 134024 336734
rect 133972 336670 134024 336676
rect 134076 322930 134104 390594
rect 134156 385756 134208 385762
rect 134156 385698 134208 385704
rect 134168 338065 134196 385698
rect 134522 359272 134578 359281
rect 134522 359207 134578 359216
rect 134154 338056 134210 338065
rect 134154 337991 134210 338000
rect 134536 337414 134564 359207
rect 135168 354680 135220 354686
rect 135168 354622 135220 354628
rect 135180 354074 135208 354622
rect 135168 354068 135220 354074
rect 135168 354010 135220 354016
rect 135166 338056 135222 338065
rect 135166 337991 135222 338000
rect 134524 337408 134576 337414
rect 135180 337385 135208 337991
rect 134524 337350 134576 337356
rect 135166 337376 135222 337385
rect 135166 337311 135222 337320
rect 134064 322924 134116 322930
rect 134064 322866 134116 322872
rect 133972 313404 134024 313410
rect 133972 313346 134024 313352
rect 133880 273216 133932 273222
rect 133880 273158 133932 273164
rect 133984 258074 134012 313346
rect 134616 298376 134668 298382
rect 134616 298318 134668 298324
rect 133892 258046 134012 258074
rect 133892 256630 133920 258046
rect 134524 256760 134576 256766
rect 134524 256702 134576 256708
rect 133880 256624 133932 256630
rect 133880 256566 133932 256572
rect 133788 242820 133840 242826
rect 133788 242762 133840 242768
rect 133800 242185 133828 242762
rect 133786 242176 133842 242185
rect 133786 242111 133842 242120
rect 133236 209296 133288 209302
rect 133236 209238 133288 209244
rect 134536 191214 134564 256702
rect 134628 247926 134656 298318
rect 134708 263628 134760 263634
rect 134708 263570 134760 263576
rect 134616 247920 134668 247926
rect 134616 247862 134668 247868
rect 134720 218890 134748 263570
rect 135168 256624 135220 256630
rect 135168 256566 135220 256572
rect 135180 256018 135208 256566
rect 135168 256012 135220 256018
rect 135168 255954 135220 255960
rect 135272 246362 135300 392158
rect 135364 338026 135392 445742
rect 135456 371890 135484 474642
rect 135916 471306 135944 560934
rect 136652 534070 136680 636822
rect 136744 561678 136772 659738
rect 139400 655580 139452 655586
rect 139400 655522 139452 655528
rect 138020 648644 138072 648650
rect 138020 648586 138072 648592
rect 136824 586560 136876 586566
rect 136824 586502 136876 586508
rect 136732 561672 136784 561678
rect 136732 561614 136784 561620
rect 136732 554124 136784 554130
rect 136732 554066 136784 554072
rect 136640 534064 136692 534070
rect 136640 534006 136692 534012
rect 135904 471300 135956 471306
rect 135904 471242 135956 471248
rect 136652 445058 136680 534006
rect 136744 463010 136772 554066
rect 136836 491201 136864 586502
rect 136914 570752 136970 570761
rect 136914 570687 136970 570696
rect 136822 491192 136878 491201
rect 136822 491127 136878 491136
rect 136928 477494 136956 570687
rect 138032 552702 138060 648586
rect 138110 565040 138166 565049
rect 138110 564975 138166 564984
rect 138020 552696 138072 552702
rect 138020 552638 138072 552644
rect 138124 480254 138152 564975
rect 139412 558890 139440 655522
rect 140780 641776 140832 641782
rect 140780 641718 140832 641724
rect 139490 570616 139546 570625
rect 139490 570551 139546 570560
rect 139400 558884 139452 558890
rect 139400 558826 139452 558832
rect 138664 548548 138716 548554
rect 138664 548490 138716 548496
rect 138032 480226 138152 480254
rect 136916 477488 136968 477494
rect 136916 477430 136968 477436
rect 138032 471986 138060 480226
rect 138020 471980 138072 471986
rect 138020 471922 138072 471928
rect 138032 471374 138060 471922
rect 138020 471368 138072 471374
rect 138020 471310 138072 471316
rect 137008 467832 137060 467838
rect 137008 467774 137060 467780
rect 136732 463004 136784 463010
rect 136732 462946 136784 462952
rect 136916 458244 136968 458250
rect 136916 458186 136968 458192
rect 136640 445052 136692 445058
rect 136640 444994 136692 445000
rect 136824 438932 136876 438938
rect 136824 438874 136876 438880
rect 135444 371884 135496 371890
rect 135444 371826 135496 371832
rect 135904 371340 135956 371346
rect 135904 371282 135956 371288
rect 135916 340882 135944 371282
rect 135904 340876 135956 340882
rect 135904 340818 135956 340824
rect 136836 338026 136864 438874
rect 136928 346390 136956 458186
rect 137020 359514 137048 467774
rect 138676 458862 138704 548490
rect 139400 543040 139452 543046
rect 139400 542982 139452 542988
rect 139308 470552 139360 470558
rect 139308 470494 139360 470500
rect 138664 458856 138716 458862
rect 138664 458798 138716 458804
rect 138664 449948 138716 449954
rect 138664 449890 138716 449896
rect 138112 394120 138164 394126
rect 138112 394062 138164 394068
rect 137284 381540 137336 381546
rect 137284 381482 137336 381488
rect 137008 359508 137060 359514
rect 137008 359450 137060 359456
rect 136916 346384 136968 346390
rect 136916 346326 136968 346332
rect 137192 346384 137244 346390
rect 137192 346326 137244 346332
rect 137204 345710 137232 346326
rect 137192 345704 137244 345710
rect 137192 345646 137244 345652
rect 135352 338020 135404 338026
rect 135352 337962 135404 337968
rect 135628 338020 135680 338026
rect 135628 337962 135680 337968
rect 136640 338020 136692 338026
rect 136640 337962 136692 337968
rect 136824 338020 136876 338026
rect 136824 337962 136876 337968
rect 135640 337414 135668 337962
rect 136652 337482 136680 337962
rect 136640 337476 136692 337482
rect 136640 337418 136692 337424
rect 135628 337408 135680 337414
rect 135628 337350 135680 337356
rect 136732 336048 136784 336054
rect 136732 335990 136784 335996
rect 136640 333260 136692 333266
rect 136640 333202 136692 333208
rect 135904 319524 135956 319530
rect 135904 319466 135956 319472
rect 135260 246356 135312 246362
rect 135260 246298 135312 246304
rect 134708 218884 134760 218890
rect 134708 218826 134760 218832
rect 135916 207738 135944 319466
rect 135996 299736 136048 299742
rect 135996 299678 136048 299684
rect 135904 207732 135956 207738
rect 135904 207674 135956 207680
rect 136008 192681 136036 299678
rect 136652 231674 136680 333202
rect 136744 263566 136772 335990
rect 136732 263560 136784 263566
rect 136732 263502 136784 263508
rect 137100 263560 137152 263566
rect 137100 263502 137152 263508
rect 137112 262886 137140 263502
rect 137100 262880 137152 262886
rect 137100 262822 137152 262828
rect 137296 243030 137324 381482
rect 138020 372020 138072 372026
rect 138020 371962 138072 371968
rect 138032 339318 138060 371962
rect 138020 339312 138072 339318
rect 138020 339254 138072 339260
rect 138124 306374 138152 394062
rect 138676 375358 138704 449890
rect 138664 375352 138716 375358
rect 138664 375294 138716 375300
rect 139032 372020 139084 372026
rect 139032 371962 139084 371968
rect 139044 371414 139072 371962
rect 139032 371408 139084 371414
rect 139032 371350 139084 371356
rect 139320 364274 139348 470494
rect 139412 451314 139440 542982
rect 139504 476066 139532 570551
rect 139584 544400 139636 544406
rect 139584 544342 139636 544348
rect 139596 543794 139624 544342
rect 140792 543794 140820 641718
rect 140872 578264 140924 578270
rect 140872 578206 140924 578212
rect 139584 543788 139636 543794
rect 139584 543730 139636 543736
rect 140780 543788 140832 543794
rect 140780 543730 140832 543736
rect 139492 476060 139544 476066
rect 139492 476002 139544 476008
rect 139596 454102 139624 543730
rect 140884 489914 140912 578206
rect 140964 573368 141016 573374
rect 140964 573310 141016 573316
rect 140792 489886 140912 489914
rect 140792 487150 140820 489886
rect 140780 487144 140832 487150
rect 140780 487086 140832 487092
rect 140792 486470 140820 487086
rect 140780 486464 140832 486470
rect 140780 486406 140832 486412
rect 140976 483041 141004 573310
rect 142172 566506 142200 663750
rect 146300 659728 146352 659734
rect 146300 659670 146352 659676
rect 143632 650072 143684 650078
rect 143632 650014 143684 650020
rect 143540 647284 143592 647290
rect 143540 647226 143592 647232
rect 142252 576156 142304 576162
rect 142252 576098 142304 576104
rect 142160 566500 142212 566506
rect 142160 566442 142212 566448
rect 142160 562352 142212 562358
rect 142160 562294 142212 562300
rect 141056 556844 141108 556850
rect 141056 556786 141108 556792
rect 140962 483032 141018 483041
rect 140962 482967 141018 482976
rect 140872 478916 140924 478922
rect 140872 478858 140924 478864
rect 139584 454096 139636 454102
rect 139584 454038 139636 454044
rect 139400 451308 139452 451314
rect 139452 451256 139532 451274
rect 139400 451250 139532 451256
rect 139412 451246 139532 451250
rect 139504 371890 139532 451246
rect 139492 371884 139544 371890
rect 139492 371826 139544 371832
rect 139504 371346 139532 371826
rect 139492 371340 139544 371346
rect 139492 371282 139544 371288
rect 139308 364268 139360 364274
rect 139308 364210 139360 364216
rect 139320 363633 139348 364210
rect 139306 363624 139362 363633
rect 139306 363559 139362 363568
rect 139596 343602 139624 454038
rect 140044 392148 140096 392154
rect 140044 392090 140096 392096
rect 139584 343596 139636 343602
rect 139584 343538 139636 343544
rect 139596 342922 139624 343538
rect 139584 342916 139636 342922
rect 139584 342858 139636 342864
rect 138204 341556 138256 341562
rect 138204 341498 138256 341504
rect 138216 340950 138244 341498
rect 138204 340944 138256 340950
rect 138204 340886 138256 340892
rect 138032 306346 138152 306374
rect 137376 304428 137428 304434
rect 137376 304370 137428 304376
rect 137284 243024 137336 243030
rect 137284 242966 137336 242972
rect 137296 242894 137324 242966
rect 137284 242888 137336 242894
rect 137284 242830 137336 242836
rect 136640 231668 136692 231674
rect 136640 231610 136692 231616
rect 135994 192672 136050 192681
rect 135994 192607 136050 192616
rect 137388 192506 137416 304370
rect 138032 300150 138060 306346
rect 138020 300144 138072 300150
rect 138018 300112 138020 300121
rect 138072 300112 138074 300121
rect 138018 300047 138074 300056
rect 137468 249824 137520 249830
rect 137468 249766 137520 249772
rect 137376 192500 137428 192506
rect 137376 192442 137428 192448
rect 134524 191208 134576 191214
rect 134524 191150 134576 191156
rect 133144 190120 133196 190126
rect 133144 190062 133196 190068
rect 124864 187060 124916 187066
rect 124864 187002 124916 187008
rect 128268 183660 128320 183666
rect 128268 183602 128320 183608
rect 126060 179580 126112 179586
rect 126060 179522 126112 179528
rect 123484 178764 123536 178770
rect 123484 178706 123536 178712
rect 116950 177712 117006 177721
rect 116950 177647 117006 177656
rect 119710 177712 119766 177721
rect 119710 177647 119766 177656
rect 121182 177712 121238 177721
rect 121182 177647 121238 177656
rect 123298 177712 123354 177721
rect 123298 177647 123354 177656
rect 126072 177177 126100 179522
rect 128280 177721 128308 183602
rect 132408 182504 132460 182510
rect 132408 182446 132460 182452
rect 130936 181076 130988 181082
rect 130936 181018 130988 181024
rect 129464 181008 129516 181014
rect 129464 180950 129516 180956
rect 129476 177721 129504 180950
rect 130948 177721 130976 181018
rect 132420 177721 132448 182446
rect 137480 181558 137508 249766
rect 138216 245614 138244 340886
rect 138664 308508 138716 308514
rect 138664 308450 138716 308456
rect 138204 245608 138256 245614
rect 138204 245550 138256 245556
rect 138676 195362 138704 308450
rect 138756 302388 138808 302394
rect 138756 302330 138808 302336
rect 138768 218822 138796 302330
rect 140056 260914 140084 392090
rect 140780 391264 140832 391270
rect 140780 391206 140832 391212
rect 140136 352572 140188 352578
rect 140136 352514 140188 352520
rect 140148 334762 140176 352514
rect 140688 335232 140740 335238
rect 140688 335174 140740 335180
rect 140700 334762 140728 335174
rect 140136 334756 140188 334762
rect 140136 334698 140188 334704
rect 140688 334756 140740 334762
rect 140688 334698 140740 334704
rect 140136 308440 140188 308446
rect 140136 308382 140188 308388
rect 140044 260908 140096 260914
rect 140044 260850 140096 260856
rect 139584 260840 139636 260846
rect 139584 260782 139636 260788
rect 139596 259554 139624 260782
rect 139584 259548 139636 259554
rect 139584 259490 139636 259496
rect 140056 234394 140084 260850
rect 140044 234388 140096 234394
rect 140044 234330 140096 234336
rect 138756 218816 138808 218822
rect 138756 218758 138808 218764
rect 138664 195356 138716 195362
rect 138664 195298 138716 195304
rect 140148 184346 140176 308382
rect 140700 260846 140728 334698
rect 140688 260840 140740 260846
rect 140688 260782 140740 260788
rect 140792 227730 140820 391206
rect 140884 373998 140912 478858
rect 140976 378146 141004 482967
rect 141068 465730 141096 556786
rect 142172 470558 142200 562294
rect 142264 485081 142292 576098
rect 142344 548616 142396 548622
rect 142344 548558 142396 548564
rect 142250 485072 142306 485081
rect 142250 485007 142306 485016
rect 142252 472660 142304 472666
rect 142252 472602 142304 472608
rect 142160 470552 142212 470558
rect 142160 470494 142212 470500
rect 141056 465724 141108 465730
rect 141056 465666 141108 465672
rect 141056 462324 141108 462330
rect 141056 462266 141108 462272
rect 140964 378140 141016 378146
rect 140964 378082 141016 378088
rect 140872 373992 140924 373998
rect 140872 373934 140924 373940
rect 140884 373318 140912 373934
rect 140872 373312 140924 373318
rect 140872 373254 140924 373260
rect 141068 371958 141096 462266
rect 142160 445052 142212 445058
rect 142160 444994 142212 445000
rect 141240 378140 141292 378146
rect 141240 378082 141292 378088
rect 141252 377466 141280 378082
rect 141240 377460 141292 377466
rect 141240 377402 141292 377408
rect 141148 375352 141200 375358
rect 141148 375294 141200 375300
rect 141160 374134 141188 375294
rect 141148 374128 141200 374134
rect 141148 374070 141200 374076
rect 141056 371952 141108 371958
rect 141056 371894 141108 371900
rect 141068 371385 141096 371894
rect 141054 371376 141110 371385
rect 141054 371311 141110 371320
rect 140870 345672 140926 345681
rect 140870 345607 140926 345616
rect 140884 345098 140912 345607
rect 140872 345092 140924 345098
rect 140872 345034 140924 345040
rect 140884 335354 140912 345034
rect 140884 335326 141004 335354
rect 140872 334620 140924 334626
rect 140872 334562 140924 334568
rect 140884 238649 140912 334562
rect 140976 251190 141004 335326
rect 141160 335306 141188 374070
rect 141424 369844 141476 369850
rect 141424 369786 141476 369792
rect 141436 350606 141464 369786
rect 141424 350600 141476 350606
rect 141424 350542 141476 350548
rect 141148 335300 141200 335306
rect 141148 335242 141200 335248
rect 142172 313274 142200 444994
rect 142264 367062 142292 472602
rect 142356 457502 142384 548558
rect 143552 548554 143580 647226
rect 143644 552022 143672 650014
rect 146312 562358 146340 659670
rect 201512 657558 201540 703258
rect 218992 700398 219020 703520
rect 218980 700392 219032 700398
rect 218980 700334 219032 700340
rect 235184 700330 235212 703520
rect 267660 703254 267688 703520
rect 267648 703248 267700 703254
rect 267648 703190 267700 703196
rect 283852 700330 283880 703520
rect 235172 700324 235224 700330
rect 235172 700266 235224 700272
rect 238024 700324 238076 700330
rect 238024 700266 238076 700272
rect 283840 700324 283892 700330
rect 283840 700266 283892 700272
rect 238036 685166 238064 700266
rect 238024 685160 238076 685166
rect 238024 685102 238076 685108
rect 201500 657552 201552 657558
rect 201500 657494 201552 657500
rect 299492 639606 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703186 332548 703520
rect 332508 703180 332560 703186
rect 332508 703122 332560 703128
rect 348804 703118 348832 703520
rect 348792 703112 348844 703118
rect 348792 703054 348844 703060
rect 364996 703050 365024 703520
rect 364340 703044 364392 703050
rect 364340 702986 364392 702992
rect 364984 703044 365036 703050
rect 364984 702986 365036 702992
rect 364352 700754 364380 702986
rect 397472 702681 397500 703520
rect 413664 702982 413692 703520
rect 413652 702976 413704 702982
rect 413652 702918 413704 702924
rect 429856 702846 429884 703520
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 429200 702840 429252 702846
rect 429200 702782 429252 702788
rect 429844 702840 429896 702846
rect 429844 702782 429896 702788
rect 397458 702672 397514 702681
rect 397458 702607 397514 702616
rect 364260 700726 364380 700754
rect 299480 639600 299532 639606
rect 299480 639542 299532 639548
rect 146300 562352 146352 562358
rect 146300 562294 146352 562300
rect 143632 552016 143684 552022
rect 143632 551958 143684 551964
rect 143540 548548 143592 548554
rect 143540 548490 143592 548496
rect 142436 537532 142488 537538
rect 142436 537474 142488 537480
rect 142448 536858 142476 537474
rect 142436 536852 142488 536858
rect 142436 536794 142488 536800
rect 142448 472666 142476 536794
rect 147772 487212 147824 487218
rect 147772 487154 147824 487160
rect 143724 481772 143776 481778
rect 143724 481714 143776 481720
rect 143540 481704 143592 481710
rect 143540 481646 143592 481652
rect 142436 472660 142488 472666
rect 142436 472602 142488 472608
rect 142528 458856 142580 458862
rect 142528 458798 142580 458804
rect 142344 457496 142396 457502
rect 142344 457438 142396 457444
rect 142252 367056 142304 367062
rect 142252 366998 142304 367004
rect 142540 354674 142568 458798
rect 143552 376718 143580 481646
rect 143632 392080 143684 392086
rect 143632 392022 143684 392028
rect 143540 376712 143592 376718
rect 143540 376654 143592 376660
rect 143538 371376 143594 371385
rect 143538 371311 143594 371320
rect 142356 354646 142568 354674
rect 142252 354000 142304 354006
rect 142252 353942 142304 353948
rect 142160 313268 142212 313274
rect 142160 313210 142212 313216
rect 141422 296032 141478 296041
rect 141422 295967 141478 295976
rect 140964 251184 141016 251190
rect 140964 251126 141016 251132
rect 140870 238640 140926 238649
rect 140870 238575 140926 238584
rect 140884 237425 140912 238575
rect 140870 237416 140926 237425
rect 140870 237351 140926 237360
rect 140780 227724 140832 227730
rect 140780 227666 140832 227672
rect 141436 185706 141464 295967
rect 141514 237416 141570 237425
rect 141514 237351 141570 237360
rect 141528 224806 141556 237351
rect 142264 235890 142292 353942
rect 142356 349042 142384 354646
rect 142436 350600 142488 350606
rect 142436 350542 142488 350548
rect 142344 349036 142396 349042
rect 142344 348978 142396 348984
rect 142448 315382 142476 350542
rect 143448 349036 143500 349042
rect 143448 348978 143500 348984
rect 143460 348537 143488 348978
rect 143446 348528 143502 348537
rect 143446 348463 143502 348472
rect 142988 316804 143040 316810
rect 142988 316746 143040 316752
rect 142436 315376 142488 315382
rect 142436 315318 142488 315324
rect 142804 309800 142856 309806
rect 142804 309742 142856 309748
rect 142252 235884 142304 235890
rect 142252 235826 142304 235832
rect 141516 224800 141568 224806
rect 141516 224742 141568 224748
rect 142816 188494 142844 309742
rect 142896 302320 142948 302326
rect 142896 302262 142948 302268
rect 142908 196722 142936 302262
rect 143000 254862 143028 316746
rect 143448 313268 143500 313274
rect 143448 313210 143500 313216
rect 143460 312662 143488 313210
rect 143448 312656 143500 312662
rect 143448 312598 143500 312604
rect 143448 255264 143500 255270
rect 143448 255206 143500 255212
rect 143460 254862 143488 255206
rect 142988 254856 143040 254862
rect 142988 254798 143040 254804
rect 143448 254856 143500 254862
rect 143448 254798 143500 254804
rect 143460 229022 143488 254798
rect 143552 238610 143580 371311
rect 143644 259418 143672 392022
rect 143736 376038 143764 481714
rect 145104 469260 145156 469266
rect 145104 469202 145156 469208
rect 143816 464364 143868 464370
rect 143816 464306 143868 464312
rect 143724 376032 143776 376038
rect 143724 375974 143776 375980
rect 143724 361616 143776 361622
rect 143724 361558 143776 361564
rect 143632 259412 143684 259418
rect 143632 259354 143684 259360
rect 143736 253201 143764 361558
rect 143828 356046 143856 464306
rect 145012 459604 145064 459610
rect 145012 459546 145064 459552
rect 144920 367056 144972 367062
rect 144920 366998 144972 367004
rect 144276 362228 144328 362234
rect 144276 362170 144328 362176
rect 144288 361622 144316 362170
rect 144276 361616 144328 361622
rect 144276 361558 144328 361564
rect 143816 356040 143868 356046
rect 143816 355982 143868 355988
rect 144828 356040 144880 356046
rect 144828 355982 144880 355988
rect 144840 355366 144868 355982
rect 144828 355360 144880 355366
rect 144828 355302 144880 355308
rect 144184 259548 144236 259554
rect 144184 259490 144236 259496
rect 143722 253192 143778 253201
rect 143722 253127 143778 253136
rect 143540 238604 143592 238610
rect 143540 238546 143592 238552
rect 143448 229016 143500 229022
rect 143448 228958 143500 228964
rect 143460 228410 143488 228958
rect 143448 228404 143500 228410
rect 143448 228346 143500 228352
rect 144196 200802 144224 259490
rect 144828 259412 144880 259418
rect 144828 259354 144880 259360
rect 144840 258738 144868 259354
rect 144828 258732 144880 258738
rect 144828 258674 144880 258680
rect 144932 238649 144960 366998
rect 145024 349110 145052 459546
rect 145116 361554 145144 469202
rect 146484 467900 146536 467906
rect 146484 467842 146536 467848
rect 146392 463004 146444 463010
rect 146392 462946 146444 462952
rect 145196 405000 145248 405006
rect 145196 404942 145248 404948
rect 145104 361548 145156 361554
rect 145104 361490 145156 361496
rect 145116 360874 145144 361490
rect 145104 360868 145156 360874
rect 145104 360810 145156 360816
rect 145208 351830 145236 404942
rect 146300 392624 146352 392630
rect 146300 392566 146352 392572
rect 145196 351824 145248 351830
rect 145196 351766 145248 351772
rect 145208 351121 145236 351766
rect 145194 351112 145250 351121
rect 145194 351047 145250 351056
rect 145012 349104 145064 349110
rect 145012 349046 145064 349052
rect 146208 349104 146260 349110
rect 146208 349046 146260 349052
rect 146220 348401 146248 349046
rect 146206 348392 146262 348401
rect 146206 348327 146262 348336
rect 145656 307148 145708 307154
rect 145656 307090 145708 307096
rect 145564 296948 145616 296954
rect 145564 296890 145616 296896
rect 144918 238640 144974 238649
rect 144918 238575 144974 238584
rect 144932 238542 144960 238575
rect 144920 238536 144972 238542
rect 144920 238478 144972 238484
rect 144184 200796 144236 200802
rect 144184 200738 144236 200744
rect 142896 196716 142948 196722
rect 142896 196658 142948 196664
rect 142804 188488 142856 188494
rect 142804 188430 142856 188436
rect 141424 185700 141476 185706
rect 141424 185642 141476 185648
rect 145576 184414 145604 296890
rect 145668 199646 145696 307090
rect 146312 248402 146340 392566
rect 146404 354686 146432 462946
rect 146496 360194 146524 467842
rect 147680 460964 147732 460970
rect 147680 460906 147732 460912
rect 146944 393508 146996 393514
rect 146944 393450 146996 393456
rect 146956 365838 146984 393450
rect 146944 365832 146996 365838
rect 146944 365774 146996 365780
rect 146956 364334 146984 365774
rect 146956 364306 147168 364334
rect 146484 360188 146536 360194
rect 146484 360130 146536 360136
rect 146496 359417 146524 360130
rect 146482 359408 146538 359417
rect 146482 359343 146538 359352
rect 146944 358080 146996 358086
rect 146944 358022 146996 358028
rect 146392 354680 146444 354686
rect 146392 354622 146444 354628
rect 146300 248396 146352 248402
rect 146300 248338 146352 248344
rect 146312 247858 146340 248338
rect 146300 247852 146352 247858
rect 146300 247794 146352 247800
rect 146956 204270 146984 358022
rect 147036 301572 147088 301578
rect 147036 301514 147088 301520
rect 146944 204264 146996 204270
rect 146944 204206 146996 204212
rect 146956 203590 146984 204206
rect 146944 203584 146996 203590
rect 146944 203526 146996 203532
rect 145656 199640 145708 199646
rect 145656 199582 145708 199588
rect 147048 187202 147076 301514
rect 147140 284306 147168 364306
rect 147692 351898 147720 460906
rect 147784 383178 147812 487154
rect 152096 486464 152148 486470
rect 152096 486406 152148 486412
rect 148968 471368 149020 471374
rect 148968 471310 149020 471316
rect 148980 470626 149008 471310
rect 149244 471300 149296 471306
rect 149244 471242 149296 471248
rect 148968 470620 149020 470626
rect 148968 470562 149020 470568
rect 147864 389904 147916 389910
rect 147864 389846 147916 389852
rect 147772 383172 147824 383178
rect 147772 383114 147824 383120
rect 147772 383036 147824 383042
rect 147772 382978 147824 382984
rect 147784 382294 147812 382978
rect 147772 382288 147824 382294
rect 147772 382230 147824 382236
rect 147680 351892 147732 351898
rect 147680 351834 147732 351840
rect 147692 351218 147720 351834
rect 147680 351212 147732 351218
rect 147680 351154 147732 351160
rect 147784 294778 147812 382230
rect 147876 297430 147904 389846
rect 148980 364410 149008 470562
rect 149152 395344 149204 395350
rect 149152 395286 149204 395292
rect 149060 376712 149112 376718
rect 149060 376654 149112 376660
rect 148968 364404 149020 364410
rect 148968 364346 149020 364352
rect 148416 305652 148468 305658
rect 148416 305594 148468 305600
rect 147864 297424 147916 297430
rect 147864 297366 147916 297372
rect 148140 297424 148192 297430
rect 148140 297366 148192 297372
rect 148152 296954 148180 297366
rect 148140 296948 148192 296954
rect 148140 296890 148192 296896
rect 147772 294772 147824 294778
rect 147772 294714 147824 294720
rect 148324 293276 148376 293282
rect 148324 293218 148376 293224
rect 147128 284300 147180 284306
rect 147128 284242 147180 284248
rect 147220 266484 147272 266490
rect 147220 266426 147272 266432
rect 147128 247920 147180 247926
rect 147128 247862 147180 247868
rect 147140 218754 147168 247862
rect 147232 240825 147260 266426
rect 147218 240816 147274 240825
rect 147218 240751 147274 240760
rect 147128 218748 147180 218754
rect 147128 218690 147180 218696
rect 147036 187196 147088 187202
rect 147036 187138 147088 187144
rect 148336 185842 148364 293218
rect 148428 291174 148456 305594
rect 148508 300280 148560 300286
rect 148508 300222 148560 300228
rect 148416 291168 148468 291174
rect 148416 291110 148468 291116
rect 148416 280220 148468 280226
rect 148416 280162 148468 280168
rect 148428 189689 148456 280162
rect 148520 223446 148548 300222
rect 148600 291168 148652 291174
rect 148600 291110 148652 291116
rect 148612 290018 148640 291110
rect 148600 290012 148652 290018
rect 148600 289954 148652 289960
rect 148612 256698 148640 289954
rect 148600 256692 148652 256698
rect 148600 256634 148652 256640
rect 149072 238746 149100 376654
rect 149164 269074 149192 395286
rect 149256 362914 149284 471242
rect 151912 465724 151964 465730
rect 151912 465666 151964 465672
rect 150532 457496 150584 457502
rect 150532 457438 150584 457444
rect 150440 456816 150492 456822
rect 150440 456758 150492 456764
rect 149244 362908 149296 362914
rect 149244 362850 149296 362856
rect 149256 362302 149284 362850
rect 149244 362296 149296 362302
rect 149244 362238 149296 362244
rect 150452 345030 150480 456758
rect 150544 346361 150572 457438
rect 151820 394732 151872 394738
rect 151820 394674 151872 394680
rect 150624 357400 150676 357406
rect 150624 357342 150676 357348
rect 150636 356114 150664 357342
rect 150624 356108 150676 356114
rect 150624 356050 150676 356056
rect 150530 346352 150586 346361
rect 150530 346287 150586 346296
rect 150544 345681 150572 346287
rect 150530 345672 150586 345681
rect 150530 345607 150586 345616
rect 150440 345024 150492 345030
rect 150440 344966 150492 344972
rect 150452 344350 150480 344966
rect 150440 344344 150492 344350
rect 150440 344286 150492 344292
rect 149704 312588 149756 312594
rect 149704 312530 149756 312536
rect 149152 269068 149204 269074
rect 149152 269010 149204 269016
rect 149336 269068 149388 269074
rect 149336 269010 149388 269016
rect 149348 268462 149376 269010
rect 149336 268456 149388 268462
rect 149336 268398 149388 268404
rect 149060 238740 149112 238746
rect 149060 238682 149112 238688
rect 148508 223440 148560 223446
rect 148508 223382 148560 223388
rect 149716 203726 149744 312530
rect 150636 282198 150664 356050
rect 151084 330608 151136 330614
rect 151084 330550 151136 330556
rect 150624 282192 150676 282198
rect 150624 282134 150676 282140
rect 149796 266416 149848 266422
rect 149796 266358 149848 266364
rect 149808 235890 149836 266358
rect 149796 235884 149848 235890
rect 149796 235826 149848 235832
rect 149704 203720 149756 203726
rect 149704 203662 149756 203668
rect 151096 194002 151124 330550
rect 151360 292732 151412 292738
rect 151360 292674 151412 292680
rect 151176 291916 151228 291922
rect 151176 291858 151228 291864
rect 151084 193996 151136 194002
rect 151084 193938 151136 193944
rect 148414 189680 148470 189689
rect 148414 189615 148470 189624
rect 151188 188562 151216 291858
rect 151268 245676 151320 245682
rect 151268 245618 151320 245624
rect 151176 188556 151228 188562
rect 151176 188498 151228 188504
rect 148324 185836 148376 185842
rect 148324 185778 148376 185784
rect 145564 184408 145616 184414
rect 145564 184350 145616 184356
rect 140136 184340 140188 184346
rect 140136 184282 140188 184288
rect 137468 181552 137520 181558
rect 137468 181494 137520 181500
rect 151280 180334 151308 245618
rect 151372 234462 151400 292674
rect 151832 279449 151860 394674
rect 151924 357406 151952 465666
rect 152004 393984 152056 393990
rect 152004 393926 152056 393932
rect 151912 357400 151964 357406
rect 151912 357342 151964 357348
rect 152016 288318 152044 393926
rect 152108 382226 152136 486406
rect 286324 484424 286376 484430
rect 286324 484366 286376 484372
rect 164884 403096 164936 403102
rect 164884 403038 164936 403044
rect 162124 401668 162176 401674
rect 162124 401610 162176 401616
rect 155222 400344 155278 400353
rect 153844 400308 153896 400314
rect 155222 400279 155278 400288
rect 153844 400250 153896 400256
rect 152096 382220 152148 382226
rect 152096 382162 152148 382168
rect 153108 382220 153160 382226
rect 153108 382162 153160 382168
rect 153120 381546 153148 382162
rect 153108 381540 153160 381546
rect 153108 381482 153160 381488
rect 153200 364404 153252 364410
rect 153200 364346 153252 364352
rect 152556 301028 152608 301034
rect 152556 300970 152608 300976
rect 152464 296948 152516 296954
rect 152464 296890 152516 296896
rect 152004 288312 152056 288318
rect 152004 288254 152056 288260
rect 151818 279440 151874 279449
rect 151818 279375 151874 279384
rect 151360 234456 151412 234462
rect 151360 234398 151412 234404
rect 152476 231606 152504 296890
rect 152568 239873 152596 300970
rect 153108 288312 153160 288318
rect 153108 288254 153160 288260
rect 153120 287706 153148 288254
rect 153108 287700 153160 287706
rect 153108 287642 153160 287648
rect 153212 285598 153240 364346
rect 153476 292664 153528 292670
rect 153476 292606 153528 292612
rect 153488 291990 153516 292606
rect 153476 291984 153528 291990
rect 153476 291926 153528 291932
rect 153200 285592 153252 285598
rect 153200 285534 153252 285540
rect 153212 284889 153240 285534
rect 153198 284880 153254 284889
rect 153198 284815 153254 284824
rect 152648 265056 152700 265062
rect 152648 264998 152700 265004
rect 152554 239864 152610 239873
rect 152554 239799 152610 239808
rect 152464 231600 152516 231606
rect 152464 231542 152516 231548
rect 152660 226273 152688 264998
rect 152646 226264 152702 226273
rect 152646 226199 152702 226208
rect 153856 184249 153884 400250
rect 154672 396772 154724 396778
rect 154672 396714 154724 396720
rect 154580 387184 154632 387190
rect 154580 387126 154632 387132
rect 154592 386510 154620 387126
rect 154580 386504 154632 386510
rect 154580 386446 154632 386452
rect 153936 291984 153988 291990
rect 153936 291926 153988 291932
rect 153948 239426 153976 291926
rect 154120 258120 154172 258126
rect 154120 258062 154172 258068
rect 154028 244316 154080 244322
rect 154028 244258 154080 244264
rect 153936 239420 153988 239426
rect 153936 239362 153988 239368
rect 154040 222154 154068 244258
rect 154132 242214 154160 258062
rect 154592 258058 154620 386446
rect 154684 292670 154712 396714
rect 154672 292664 154724 292670
rect 154672 292606 154724 292612
rect 154580 258052 154632 258058
rect 154580 257994 154632 258000
rect 154120 242208 154172 242214
rect 154120 242150 154172 242156
rect 154028 222148 154080 222154
rect 154028 222090 154080 222096
rect 153842 184240 153898 184249
rect 155236 184210 155264 400279
rect 160744 399492 160796 399498
rect 160744 399434 160796 399440
rect 159364 399016 159416 399022
rect 159364 398958 159416 398964
rect 157984 398132 158036 398138
rect 157984 398074 158036 398080
rect 155960 377460 156012 377466
rect 155960 377402 156012 377408
rect 155972 376854 156000 377402
rect 155960 376848 156012 376854
rect 155960 376790 156012 376796
rect 155316 300212 155368 300218
rect 155316 300154 155368 300160
rect 155328 226234 155356 300154
rect 155408 292800 155460 292806
rect 155408 292742 155460 292748
rect 155420 233034 155448 292742
rect 155500 252612 155552 252618
rect 155500 252554 155552 252560
rect 155512 238066 155540 252554
rect 155972 252550 156000 376790
rect 156696 298444 156748 298450
rect 156696 298386 156748 298392
rect 156604 289944 156656 289950
rect 156604 289886 156656 289892
rect 155960 252544 156012 252550
rect 155960 252486 156012 252492
rect 155500 238060 155552 238066
rect 155500 238002 155552 238008
rect 155408 233028 155460 233034
rect 155408 232970 155460 232976
rect 155316 226228 155368 226234
rect 155316 226170 155368 226176
rect 156616 203794 156644 289886
rect 156708 220794 156736 298386
rect 156696 220788 156748 220794
rect 156696 220730 156748 220736
rect 157996 214606 158024 398074
rect 158076 302456 158128 302462
rect 158076 302398 158128 302404
rect 158088 221950 158116 302398
rect 158168 264988 158220 264994
rect 158168 264930 158220 264936
rect 158180 240786 158208 264930
rect 158168 240780 158220 240786
rect 158168 240722 158220 240728
rect 158076 221944 158128 221950
rect 158076 221886 158128 221892
rect 157984 214600 158036 214606
rect 157984 214542 158036 214548
rect 156604 203788 156656 203794
rect 156604 203730 156656 203736
rect 153842 184175 153898 184184
rect 155224 184204 155276 184210
rect 155224 184146 155276 184152
rect 159376 181626 159404 398958
rect 159456 388544 159508 388550
rect 159456 388486 159508 388492
rect 159364 181620 159416 181626
rect 159364 181562 159416 181568
rect 151268 180328 151320 180334
rect 151268 180270 151320 180276
rect 134708 179648 134760 179654
rect 134708 179590 134760 179596
rect 128266 177712 128322 177721
rect 128266 177647 128322 177656
rect 129462 177712 129518 177721
rect 129462 177647 129518 177656
rect 130934 177712 130990 177721
rect 130934 177647 130990 177656
rect 132406 177712 132462 177721
rect 132406 177647 132462 177656
rect 134720 177177 134748 179590
rect 148232 178288 148284 178294
rect 148232 178230 148284 178236
rect 115846 177168 115902 177177
rect 115846 177103 115902 177112
rect 126058 177168 126114 177177
rect 126058 177103 126114 177112
rect 134706 177168 134762 177177
rect 134706 177103 134762 177112
rect 128176 177064 128228 177070
rect 128176 177006 128228 177012
rect 124496 176996 124548 177002
rect 124496 176938 124548 176944
rect 124508 176769 124536 176938
rect 128188 176769 128216 177006
rect 136088 176792 136140 176798
rect 97814 176760 97870 176769
rect 97814 176695 97870 176704
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 108118 176760 108174 176769
rect 108118 176695 108174 176704
rect 112258 176760 112314 176769
rect 112258 176695 112314 176704
rect 114374 176760 114430 176769
rect 114374 176695 114430 176704
rect 124494 176760 124550 176769
rect 124494 176695 124550 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 133142 176760 133198 176769
rect 133142 176695 133144 176704
rect 133196 176695 133198 176704
rect 136086 176760 136088 176769
rect 148244 176769 148272 178230
rect 159468 177449 159496 388486
rect 159640 298308 159692 298314
rect 159640 298250 159692 298256
rect 159548 296880 159600 296886
rect 159548 296822 159600 296828
rect 159560 202162 159588 296822
rect 159652 238134 159680 298250
rect 159640 238128 159692 238134
rect 159640 238070 159692 238076
rect 159548 202156 159600 202162
rect 159548 202098 159600 202104
rect 160756 180130 160784 399434
rect 160836 368620 160888 368626
rect 160836 368562 160888 368568
rect 160848 323678 160876 368562
rect 160836 323672 160888 323678
rect 160836 323614 160888 323620
rect 160836 296812 160888 296818
rect 160836 296754 160888 296760
rect 160848 267034 160876 296754
rect 160836 267028 160888 267034
rect 160836 266970 160888 266976
rect 160928 261520 160980 261526
rect 160928 261462 160980 261468
rect 160836 247784 160888 247790
rect 160836 247726 160888 247732
rect 160744 180124 160796 180130
rect 160744 180066 160796 180072
rect 159454 177440 159510 177449
rect 159454 177375 159510 177384
rect 160100 177064 160152 177070
rect 160100 177006 160152 177012
rect 158904 176928 158956 176934
rect 158904 176870 158956 176876
rect 158916 176769 158944 176870
rect 136140 176760 136142 176769
rect 136086 176695 136142 176704
rect 148230 176760 148286 176769
rect 148230 176695 148286 176704
rect 158902 176760 158958 176769
rect 158902 176695 158958 176704
rect 133144 176666 133196 176672
rect 118424 176316 118476 176322
rect 118424 176258 118476 176264
rect 102048 176112 102100 176118
rect 102048 176054 102100 176060
rect 98368 176044 98420 176050
rect 98368 175986 98420 175992
rect 98380 175409 98408 175986
rect 102060 175409 102088 176054
rect 118436 175409 118464 176258
rect 160112 176186 160140 177006
rect 160100 176180 160152 176186
rect 160100 176122 160152 176128
rect 121920 175976 121972 175982
rect 160848 175953 160876 247726
rect 160940 196654 160968 261462
rect 161020 253972 161072 253978
rect 161020 253914 161072 253920
rect 161032 233170 161060 253914
rect 161020 233164 161072 233170
rect 161020 233106 161072 233112
rect 160928 196648 160980 196654
rect 160928 196590 160980 196596
rect 162136 178702 162164 401610
rect 163504 378820 163556 378826
rect 163504 378762 163556 378768
rect 162216 365968 162268 365974
rect 162216 365910 162268 365916
rect 162228 327962 162256 365910
rect 162216 327956 162268 327962
rect 162216 327898 162268 327904
rect 162216 324964 162268 324970
rect 162216 324906 162268 324912
rect 162228 228818 162256 324906
rect 162306 298208 162362 298217
rect 162306 298143 162362 298152
rect 162320 231713 162348 298143
rect 162400 274712 162452 274718
rect 162400 274654 162452 274660
rect 162412 237318 162440 274654
rect 162400 237312 162452 237318
rect 162400 237254 162452 237260
rect 162306 231704 162362 231713
rect 162306 231639 162362 231648
rect 162216 228812 162268 228818
rect 162216 228754 162268 228760
rect 162216 222896 162268 222902
rect 162216 222838 162268 222844
rect 162228 198218 162256 222838
rect 162216 198212 162268 198218
rect 162216 198154 162268 198160
rect 162124 178696 162176 178702
rect 162124 178638 162176 178644
rect 163516 176254 163544 378762
rect 163596 300144 163648 300150
rect 163596 300086 163648 300092
rect 163608 234433 163636 300086
rect 163688 279472 163740 279478
rect 163688 279414 163740 279420
rect 163594 234424 163650 234433
rect 163594 234359 163650 234368
rect 163700 220250 163728 279414
rect 163688 220244 163740 220250
rect 163688 220186 163740 220192
rect 164896 181665 164924 403038
rect 228364 398948 228416 398954
rect 228364 398890 228416 398896
rect 220084 392012 220136 392018
rect 220084 391954 220136 391960
rect 169022 390824 169078 390833
rect 169022 390759 169078 390768
rect 167644 386572 167696 386578
rect 167644 386514 167696 386520
rect 166264 367328 166316 367334
rect 166264 367270 166316 367276
rect 166276 333266 166304 367270
rect 166356 362228 166408 362234
rect 166356 362170 166408 362176
rect 166264 333260 166316 333266
rect 166264 333202 166316 333208
rect 165528 331288 165580 331294
rect 165528 331230 165580 331236
rect 165068 287700 165120 287706
rect 165068 287642 165120 287648
rect 164976 247716 165028 247722
rect 164976 247658 165028 247664
rect 164988 190058 165016 247658
rect 165080 235754 165108 287642
rect 165068 235748 165120 235754
rect 165068 235690 165120 235696
rect 165540 207942 165568 331230
rect 166264 300892 166316 300898
rect 166264 300834 166316 300840
rect 166276 214810 166304 300834
rect 166368 288386 166396 362170
rect 166448 299532 166500 299538
rect 166448 299474 166500 299480
rect 166356 288380 166408 288386
rect 166356 288322 166408 288328
rect 166356 256012 166408 256018
rect 166356 255954 166408 255960
rect 166368 230489 166396 255954
rect 166460 250481 166488 299474
rect 166540 258732 166592 258738
rect 166540 258674 166592 258680
rect 166446 250472 166502 250481
rect 166446 250407 166502 250416
rect 166552 237250 166580 258674
rect 166540 237244 166592 237250
rect 166540 237186 166592 237192
rect 166354 230480 166410 230489
rect 166354 230415 166410 230424
rect 166356 228472 166408 228478
rect 166356 228414 166408 228420
rect 166264 214804 166316 214810
rect 166264 214746 166316 214752
rect 165528 207936 165580 207942
rect 165528 207878 165580 207884
rect 164976 190052 165028 190058
rect 164976 189994 165028 190000
rect 164976 182504 165028 182510
rect 164976 182446 165028 182452
rect 164882 181656 164938 181665
rect 164882 181591 164938 181600
rect 163504 176248 163556 176254
rect 163504 176190 163556 176196
rect 121920 175918 121972 175924
rect 160834 175944 160890 175953
rect 121932 175409 121960 175918
rect 160834 175879 160890 175888
rect 98366 175400 98422 175409
rect 98366 175335 98422 175344
rect 102046 175400 102102 175409
rect 102046 175335 102102 175344
rect 118422 175400 118478 175409
rect 118422 175335 118478 175344
rect 121918 175400 121974 175409
rect 121918 175335 121974 175344
rect 164988 173874 165016 182446
rect 165436 179648 165488 179654
rect 165436 179590 165488 179596
rect 165252 176996 165304 177002
rect 165252 176938 165304 176944
rect 165264 174554 165292 176938
rect 165448 175234 165476 179590
rect 166264 179512 166316 179518
rect 166264 179454 166316 179460
rect 165436 175228 165488 175234
rect 165436 175170 165488 175176
rect 165252 174548 165304 174554
rect 165252 174490 165304 174496
rect 164976 173868 165028 173874
rect 164976 173810 165028 173816
rect 166276 165578 166304 179454
rect 166368 178838 166396 228414
rect 167656 204921 167684 386514
rect 167736 358896 167788 358902
rect 167736 358838 167788 358844
rect 167748 316742 167776 358838
rect 167736 316736 167788 316742
rect 167736 316678 167788 316684
rect 167736 304292 167788 304298
rect 167736 304234 167788 304240
rect 167748 220182 167776 304234
rect 168288 289196 168340 289202
rect 168288 289138 168340 289144
rect 168300 288454 168328 289138
rect 168288 288448 168340 288454
rect 168288 288390 168340 288396
rect 167736 220176 167788 220182
rect 167736 220118 167788 220124
rect 167642 204912 167698 204921
rect 167642 204847 167698 204856
rect 168300 181762 168328 288390
rect 169036 222873 169064 390759
rect 177302 387968 177358 387977
rect 177302 387903 177358 387912
rect 184204 387932 184256 387938
rect 171784 376916 171836 376922
rect 171784 376858 171836 376864
rect 170404 372836 170456 372842
rect 170404 372778 170456 372784
rect 169116 370116 169168 370122
rect 169116 370058 169168 370064
rect 169128 327758 169156 370058
rect 169208 365900 169260 365906
rect 169208 365842 169260 365848
rect 169220 330750 169248 365842
rect 170416 336025 170444 372778
rect 170496 339516 170548 339522
rect 170496 339458 170548 339464
rect 170402 336016 170458 336025
rect 170402 335951 170458 335960
rect 169208 330744 169260 330750
rect 169208 330686 169260 330692
rect 169668 328500 169720 328506
rect 169668 328442 169720 328448
rect 169116 327752 169168 327758
rect 169116 327694 169168 327700
rect 169116 305040 169168 305046
rect 169116 304982 169168 304988
rect 169022 222864 169078 222873
rect 169022 222799 169078 222808
rect 169024 185020 169076 185026
rect 169024 184962 169076 184968
rect 168288 181756 168340 181762
rect 168288 181698 168340 181704
rect 166540 181076 166592 181082
rect 166540 181018 166592 181024
rect 166356 178832 166408 178838
rect 166356 178774 166408 178780
rect 166448 178220 166500 178226
rect 166448 178162 166500 178168
rect 166356 176316 166408 176322
rect 166356 176258 166408 176264
rect 166368 167006 166396 176258
rect 166356 167000 166408 167006
rect 166356 166942 166408 166948
rect 166264 165572 166316 165578
rect 166264 165514 166316 165520
rect 166460 165510 166488 178162
rect 166552 173806 166580 181018
rect 167920 181008 167972 181014
rect 167920 180950 167972 180956
rect 167828 180940 167880 180946
rect 167828 180882 167880 180888
rect 167734 177032 167790 177041
rect 167734 176967 167790 176976
rect 166540 173800 166592 173806
rect 166540 173742 166592 173748
rect 167642 171592 167698 171601
rect 167642 171527 167698 171536
rect 166448 165504 166500 165510
rect 166448 165446 166500 165452
rect 167656 153882 167684 171527
rect 167748 160070 167776 176967
rect 167840 168366 167868 180882
rect 167932 172514 167960 180950
rect 168012 179580 168064 179586
rect 168012 179522 168064 179528
rect 167920 172508 167972 172514
rect 167920 172450 167972 172456
rect 168024 171086 168052 179522
rect 168012 171080 168064 171086
rect 168012 171022 168064 171028
rect 167828 168360 167880 168366
rect 167828 168302 167880 168308
rect 167736 160064 167788 160070
rect 167736 160006 167788 160012
rect 169036 157350 169064 184962
rect 169128 180033 169156 304982
rect 169208 289876 169260 289882
rect 169208 289818 169260 289824
rect 169220 180402 169248 289818
rect 169680 209166 169708 328442
rect 170508 321638 170536 339458
rect 171796 327826 171824 376858
rect 174636 370048 174688 370054
rect 174636 369990 174688 369996
rect 171876 364540 171928 364546
rect 171876 364482 171928 364488
rect 171784 327820 171836 327826
rect 171784 327762 171836 327768
rect 171888 326466 171916 364482
rect 173254 359408 173310 359417
rect 173254 359343 173310 359352
rect 173164 335368 173216 335374
rect 173164 335310 173216 335316
rect 171968 327956 172020 327962
rect 171968 327898 172020 327904
rect 171876 326460 171928 326466
rect 171876 326402 171928 326408
rect 170588 325712 170640 325718
rect 170588 325654 170640 325660
rect 170496 321632 170548 321638
rect 170496 321574 170548 321580
rect 170404 281580 170456 281586
rect 170404 281522 170456 281528
rect 169668 209160 169720 209166
rect 169668 209102 169720 209108
rect 169208 180396 169260 180402
rect 169208 180338 169260 180344
rect 169114 180024 169170 180033
rect 169114 179959 169170 179968
rect 169300 179444 169352 179450
rect 169300 179386 169352 179392
rect 169116 176860 169168 176866
rect 169116 176802 169168 176808
rect 169128 161430 169156 176802
rect 169312 162858 169340 179386
rect 170416 178974 170444 281522
rect 170508 227730 170536 321574
rect 170600 234530 170628 325654
rect 171784 306468 171836 306474
rect 171784 306410 171836 306416
rect 171796 306374 171824 306410
rect 171980 306374 172008 327898
rect 173176 325718 173204 335310
rect 173164 325712 173216 325718
rect 173164 325654 173216 325660
rect 172426 320240 172482 320249
rect 172426 320175 172428 320184
rect 172480 320175 172482 320184
rect 172428 320146 172480 320152
rect 171796 306346 172008 306374
rect 170680 259480 170732 259486
rect 170680 259422 170732 259428
rect 170588 234524 170640 234530
rect 170588 234466 170640 234472
rect 170496 227724 170548 227730
rect 170496 227666 170548 227672
rect 170404 178968 170456 178974
rect 170404 178910 170456 178916
rect 170496 178288 170548 178294
rect 170496 178230 170548 178236
rect 170404 176044 170456 176050
rect 170404 175986 170456 175992
rect 169300 162852 169352 162858
rect 169300 162794 169352 162800
rect 169116 161424 169168 161430
rect 169116 161366 169168 161372
rect 169024 157344 169076 157350
rect 169024 157286 169076 157292
rect 170416 155922 170444 175986
rect 170404 155916 170456 155922
rect 170404 155858 170456 155864
rect 167644 153876 167696 153882
rect 167644 153818 167696 153824
rect 170508 150414 170536 178230
rect 170600 177313 170628 234466
rect 170692 181694 170720 259422
rect 171796 184278 171824 306346
rect 171968 303680 172020 303686
rect 171968 303622 172020 303628
rect 171876 273352 171928 273358
rect 171876 273294 171928 273300
rect 171784 184272 171836 184278
rect 171784 184214 171836 184220
rect 170772 182436 170824 182442
rect 170772 182378 170824 182384
rect 170680 181688 170732 181694
rect 170680 181630 170732 181636
rect 170586 177304 170642 177313
rect 170586 177239 170642 177248
rect 170784 160002 170812 182378
rect 170864 180872 170916 180878
rect 170864 180814 170916 180820
rect 170876 166938 170904 180814
rect 171784 176112 171836 176118
rect 171784 176054 171836 176060
rect 170864 166932 170916 166938
rect 170864 166874 170916 166880
rect 170772 159996 170824 160002
rect 170772 159938 170824 159944
rect 171796 158710 171824 176054
rect 171888 176050 171916 273294
rect 171980 233986 172008 303622
rect 171968 233980 172020 233986
rect 171968 233922 172020 233928
rect 172440 218958 172468 320146
rect 173164 318096 173216 318102
rect 173164 318038 173216 318044
rect 173176 221513 173204 318038
rect 173268 294710 173296 359343
rect 174542 337376 174598 337385
rect 174542 337311 174598 337320
rect 173256 294704 173308 294710
rect 173256 294646 173308 294652
rect 173348 281580 173400 281586
rect 173348 281522 173400 281528
rect 173256 270564 173308 270570
rect 173256 270506 173308 270512
rect 173162 221504 173218 221513
rect 173162 221439 173218 221448
rect 172428 218952 172480 218958
rect 172428 218894 172480 218900
rect 173268 187270 173296 270506
rect 173360 235958 173388 281522
rect 173440 247852 173492 247858
rect 173440 247794 173492 247800
rect 173348 235952 173400 235958
rect 173348 235894 173400 235900
rect 173256 187264 173308 187270
rect 173256 187206 173308 187212
rect 173360 186998 173388 235894
rect 173452 229022 173480 247794
rect 173440 229016 173492 229022
rect 173440 228958 173492 228964
rect 173348 186992 173400 186998
rect 173348 186934 173400 186940
rect 173164 184952 173216 184958
rect 173164 184894 173216 184900
rect 171968 178152 172020 178158
rect 171968 178094 172020 178100
rect 171876 176044 171928 176050
rect 171876 175986 171928 175992
rect 171980 164218 172008 178094
rect 171968 164212 172020 164218
rect 171968 164154 172020 164160
rect 171784 158704 171836 158710
rect 171784 158646 171836 158652
rect 173176 157282 173204 184894
rect 173164 157276 173216 157282
rect 173164 157218 173216 157224
rect 173164 153264 173216 153270
rect 173164 153206 173216 153212
rect 170496 150408 170548 150414
rect 170496 150350 170548 150356
rect 171784 146328 171836 146334
rect 171784 146270 171836 146276
rect 166264 144968 166316 144974
rect 166264 144910 166316 144916
rect 67638 126304 67694 126313
rect 67638 126239 67694 126248
rect 67652 91089 67680 126239
rect 68284 100768 68336 100774
rect 68284 100710 68336 100716
rect 67638 91080 67694 91089
rect 67638 91015 67694 91024
rect 68296 80034 68324 100710
rect 165252 98048 165304 98054
rect 165252 97990 165304 97996
rect 164882 95160 164938 95169
rect 164882 95095 164938 95104
rect 85578 94752 85634 94761
rect 85578 94687 85634 94696
rect 112350 94752 112406 94761
rect 112350 94687 112406 94696
rect 125414 94752 125470 94761
rect 125414 94687 125470 94696
rect 85592 93906 85620 94687
rect 112364 93974 112392 94687
rect 125428 94042 125456 94687
rect 161480 94580 161532 94586
rect 161480 94522 161532 94528
rect 130384 94512 130436 94518
rect 130384 94454 130436 94460
rect 125416 94036 125468 94042
rect 125416 93978 125468 93984
rect 112352 93968 112404 93974
rect 112352 93910 112404 93916
rect 85580 93900 85632 93906
rect 85580 93842 85632 93848
rect 118238 93664 118294 93673
rect 118238 93599 118294 93608
rect 98550 93528 98606 93537
rect 98550 93463 98606 93472
rect 98564 93158 98592 93463
rect 118252 93362 118280 93599
rect 129462 93528 129518 93537
rect 129462 93463 129518 93472
rect 118240 93356 118292 93362
rect 118240 93298 118292 93304
rect 103334 93256 103390 93265
rect 103334 93191 103390 93200
rect 110142 93256 110198 93265
rect 129476 93226 129504 93463
rect 110142 93191 110198 93200
rect 129464 93220 129516 93226
rect 98552 93152 98604 93158
rect 98552 93094 98604 93100
rect 85118 92440 85174 92449
rect 85118 92375 85174 92384
rect 86774 92440 86830 92449
rect 86774 92375 86830 92384
rect 88982 92440 89038 92449
rect 88982 92375 89038 92384
rect 75366 91216 75422 91225
rect 75366 91151 75422 91160
rect 75380 86970 75408 91151
rect 85132 91118 85160 92375
rect 86788 92206 86816 92375
rect 88996 92274 89024 92375
rect 88984 92268 89036 92274
rect 88984 92210 89036 92216
rect 86776 92200 86828 92206
rect 86776 92142 86828 92148
rect 90546 91760 90602 91769
rect 90546 91695 90602 91704
rect 95054 91760 95110 91769
rect 95054 91695 95110 91704
rect 88062 91216 88118 91225
rect 88062 91151 88118 91160
rect 85120 91112 85172 91118
rect 85120 91054 85172 91060
rect 75368 86964 75420 86970
rect 75368 86906 75420 86912
rect 88076 85542 88104 91151
rect 90560 89690 90588 91695
rect 92386 91216 92442 91225
rect 92386 91151 92442 91160
rect 93766 91216 93822 91225
rect 93766 91151 93822 91160
rect 90548 89684 90600 89690
rect 90548 89626 90600 89632
rect 88064 85536 88116 85542
rect 88064 85478 88116 85484
rect 92400 83978 92428 91151
rect 92388 83972 92440 83978
rect 92388 83914 92440 83920
rect 68284 80028 68336 80034
rect 68284 79970 68336 79976
rect 93780 79966 93808 91151
rect 95068 89622 95096 91695
rect 101862 91488 101918 91497
rect 101862 91423 101918 91432
rect 97906 91352 97962 91361
rect 97906 91287 97962 91296
rect 99194 91352 99250 91361
rect 99194 91287 99250 91296
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97814 91216 97870 91225
rect 97814 91151 97870 91160
rect 95056 89616 95108 89622
rect 95056 89558 95108 89564
rect 93768 79960 93820 79966
rect 93768 79902 93820 79908
rect 95160 78606 95188 91151
rect 96540 84046 96568 91151
rect 96528 84040 96580 84046
rect 96528 83982 96580 83988
rect 97828 81190 97856 91151
rect 97816 81184 97868 81190
rect 97816 81126 97868 81132
rect 97920 79762 97948 91287
rect 99208 81394 99236 91287
rect 99286 91216 99342 91225
rect 99286 91151 99342 91160
rect 100206 91216 100262 91225
rect 100206 91151 100262 91160
rect 100574 91216 100630 91225
rect 100574 91151 100630 91160
rect 99196 81388 99248 81394
rect 99196 81330 99248 81336
rect 97908 79756 97960 79762
rect 97908 79698 97960 79704
rect 95148 78600 95200 78606
rect 99300 78577 99328 91151
rect 100220 86766 100248 91151
rect 100588 88330 100616 91151
rect 100576 88324 100628 88330
rect 100576 88266 100628 88272
rect 100208 86760 100260 86766
rect 100208 86702 100260 86708
rect 101876 85338 101904 91423
rect 102046 91352 102102 91361
rect 102046 91287 102102 91296
rect 101954 91216 102010 91225
rect 101954 91151 102010 91160
rect 101864 85332 101916 85338
rect 101864 85274 101916 85280
rect 101968 82686 101996 91151
rect 101956 82680 102008 82686
rect 101956 82622 102008 82628
rect 102060 79830 102088 91287
rect 103348 89554 103376 93191
rect 110156 92478 110184 93191
rect 129464 93162 129516 93168
rect 110144 92472 110196 92478
rect 107750 92440 107806 92449
rect 110144 92414 110196 92420
rect 114374 92440 114430 92449
rect 107750 92375 107806 92384
rect 114374 92375 114430 92384
rect 115478 92440 115534 92449
rect 115478 92375 115534 92384
rect 120354 92440 120410 92449
rect 120354 92375 120356 92384
rect 107290 91352 107346 91361
rect 107290 91287 107346 91296
rect 103426 91216 103482 91225
rect 103426 91151 103482 91160
rect 104438 91216 104494 91225
rect 104438 91151 104494 91160
rect 104806 91216 104862 91225
rect 104806 91151 104862 91160
rect 105542 91216 105598 91225
rect 105542 91151 105598 91160
rect 106094 91216 106150 91225
rect 106094 91151 106150 91160
rect 103336 89548 103388 89554
rect 103336 89490 103388 89496
rect 103440 84114 103468 91151
rect 104452 88262 104480 91151
rect 104440 88256 104492 88262
rect 104440 88198 104492 88204
rect 103428 84108 103480 84114
rect 103428 84050 103480 84056
rect 104820 81433 104848 91151
rect 105556 86902 105584 91151
rect 105544 86896 105596 86902
rect 105544 86838 105596 86844
rect 106108 86834 106136 91151
rect 107304 88126 107332 91287
rect 107566 91216 107622 91225
rect 107566 91151 107622 91160
rect 107292 88120 107344 88126
rect 107292 88062 107344 88068
rect 106096 86828 106148 86834
rect 106096 86770 106148 86776
rect 107580 82754 107608 91151
rect 107764 90914 107792 92375
rect 110234 91352 110290 91361
rect 110234 91287 110290 91296
rect 108946 91216 109002 91225
rect 108946 91151 109002 91160
rect 107752 90908 107804 90914
rect 107752 90850 107804 90856
rect 108960 82822 108988 91151
rect 108948 82816 109000 82822
rect 108948 82758 109000 82764
rect 107568 82748 107620 82754
rect 107568 82690 107620 82696
rect 104806 81424 104862 81433
rect 104806 81359 104862 81368
rect 110248 81258 110276 91287
rect 110326 91216 110382 91225
rect 110326 91151 110382 91160
rect 111246 91216 111302 91225
rect 111246 91151 111302 91160
rect 112442 91216 112498 91225
rect 112442 91151 112498 91160
rect 110236 81252 110288 81258
rect 110236 81194 110288 81200
rect 102048 79824 102100 79830
rect 102048 79766 102100 79772
rect 95148 78542 95200 78548
rect 99286 78568 99342 78577
rect 110340 78538 110368 91151
rect 111260 85270 111288 91151
rect 112456 85513 112484 91151
rect 114388 90982 114416 92375
rect 115492 92342 115520 92375
rect 120408 92375 120410 92384
rect 122102 92440 122158 92449
rect 122102 92375 122158 92384
rect 120356 92346 120408 92352
rect 115480 92336 115532 92342
rect 115480 92278 115532 92284
rect 117134 91352 117190 91361
rect 117134 91287 117190 91296
rect 119894 91352 119950 91361
rect 119894 91287 119950 91296
rect 114466 91216 114522 91225
rect 114466 91151 114522 91160
rect 114926 91216 114982 91225
rect 114926 91151 114982 91160
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 114376 90976 114428 90982
rect 114376 90918 114428 90924
rect 112442 85504 112498 85513
rect 112442 85439 112498 85448
rect 111248 85264 111300 85270
rect 111248 85206 111300 85212
rect 114480 78674 114508 91151
rect 114940 87990 114968 91151
rect 114928 87984 114980 87990
rect 114928 87926 114980 87932
rect 115860 86630 115888 91151
rect 115848 86624 115900 86630
rect 115848 86566 115900 86572
rect 117148 83910 117176 91287
rect 117226 91216 117282 91225
rect 117226 91151 117282 91160
rect 117136 83904 117188 83910
rect 117136 83846 117188 83852
rect 117240 82618 117268 91151
rect 117228 82612 117280 82618
rect 117228 82554 117280 82560
rect 119908 82550 119936 91287
rect 119986 91216 120042 91225
rect 119986 91151 120042 91160
rect 120630 91216 120686 91225
rect 120630 91151 120686 91160
rect 119896 82544 119948 82550
rect 119896 82486 119948 82492
rect 120000 81326 120028 91151
rect 120644 85406 120672 91151
rect 120724 91112 120776 91118
rect 120724 91054 120776 91060
rect 120632 85400 120684 85406
rect 120632 85342 120684 85348
rect 119988 81320 120040 81326
rect 119988 81262 120040 81268
rect 114468 78668 114520 78674
rect 114468 78610 114520 78616
rect 99286 78503 99342 78512
rect 110328 78532 110380 78538
rect 110328 78474 110380 78480
rect 120736 77246 120764 91054
rect 122116 90846 122144 92375
rect 130396 92206 130424 94454
rect 133142 93528 133198 93537
rect 133142 93463 133198 93472
rect 151726 93528 151782 93537
rect 151726 93463 151782 93472
rect 133156 93294 133184 93463
rect 151740 93430 151768 93463
rect 151728 93424 151780 93430
rect 151728 93366 151780 93372
rect 133144 93288 133196 93294
rect 133144 93230 133196 93236
rect 130750 92440 130806 92449
rect 130750 92375 130806 92384
rect 135166 92440 135222 92449
rect 135166 92375 135222 92384
rect 136086 92440 136142 92449
rect 136086 92375 136142 92384
rect 151634 92440 151690 92449
rect 151634 92375 151690 92384
rect 130764 92206 130792 92375
rect 130384 92200 130436 92206
rect 130384 92142 130436 92148
rect 130752 92200 130804 92206
rect 130752 92142 130804 92148
rect 126518 91760 126574 91769
rect 126518 91695 126574 91704
rect 122838 91488 122894 91497
rect 122838 91423 122894 91432
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 122104 90840 122156 90846
rect 122104 90782 122156 90788
rect 122760 82482 122788 91151
rect 122852 89418 122880 91423
rect 123298 91216 123354 91225
rect 123298 91151 123354 91160
rect 123942 91216 123998 91225
rect 123942 91151 123998 91160
rect 124770 91216 124826 91225
rect 124770 91151 124826 91160
rect 122840 89412 122892 89418
rect 122840 89354 122892 89360
rect 123312 86698 123340 91151
rect 123300 86692 123352 86698
rect 123300 86634 123352 86640
rect 122748 82476 122800 82482
rect 122748 82418 122800 82424
rect 120724 77240 120776 77246
rect 120724 77182 120776 77188
rect 123956 77178 123984 91151
rect 124784 88194 124812 91151
rect 126532 89486 126560 91695
rect 126886 91216 126942 91225
rect 126886 91151 126942 91160
rect 127622 91216 127678 91225
rect 127622 91151 127678 91160
rect 132406 91216 132462 91225
rect 132406 91151 132462 91160
rect 126520 89480 126572 89486
rect 126520 89422 126572 89428
rect 124772 88188 124824 88194
rect 124772 88130 124824 88136
rect 126900 79898 126928 91151
rect 127636 85474 127664 91151
rect 127624 85468 127676 85474
rect 127624 85410 127676 85416
rect 132420 83842 132448 91151
rect 135180 90710 135208 92375
rect 136100 92138 136128 92375
rect 136088 92132 136140 92138
rect 136088 92074 136140 92080
rect 151450 91216 151506 91225
rect 151450 91151 151506 91160
rect 135168 90704 135220 90710
rect 135168 90646 135220 90652
rect 151464 88058 151492 91151
rect 151648 90778 151676 92375
rect 153014 91488 153070 91497
rect 153014 91423 153070 91432
rect 151636 90772 151688 90778
rect 151636 90714 151688 90720
rect 153028 89350 153056 91423
rect 161492 90914 161520 94522
rect 161480 90908 161532 90914
rect 161480 90850 161532 90856
rect 153016 89344 153068 89350
rect 153016 89286 153068 89292
rect 151452 88052 151504 88058
rect 151452 87994 151504 88000
rect 132408 83836 132460 83842
rect 132408 83778 132460 83784
rect 126888 79892 126940 79898
rect 126888 79834 126940 79840
rect 128360 77988 128412 77994
rect 128360 77930 128412 77936
rect 123944 77172 123996 77178
rect 123944 77114 123996 77120
rect 102140 76560 102192 76566
rect 102140 76502 102192 76508
rect 93860 75268 93912 75274
rect 93860 75210 93912 75216
rect 86960 73908 87012 73914
rect 86960 73850 87012 73856
rect 80060 71120 80112 71126
rect 80060 71062 80112 71068
rect 73160 64184 73212 64190
rect 73160 64126 73212 64132
rect 67640 54596 67692 54602
rect 67640 54538 67692 54544
rect 67548 21412 67600 21418
rect 67548 21354 67600 21360
rect 63512 16546 64368 16574
rect 66272 16546 66760 16574
rect 63132 5500 63184 5506
rect 63132 5442 63184 5448
rect 63052 3454 63264 3482
rect 63236 480 63264 3454
rect 64340 480 64368 16546
rect 65524 9036 65576 9042
rect 65524 8978 65576 8984
rect 65536 480 65564 8978
rect 66732 480 66760 16546
rect 61998 354 62110 480
rect 61580 326 62110 354
rect 61998 -960 62110 326
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 54538
rect 70400 51808 70452 51814
rect 70400 51750 70452 51756
rect 69020 21548 69072 21554
rect 69020 21490 69072 21496
rect 69032 6914 69060 21490
rect 69112 17332 69164 17338
rect 69112 17274 69164 17280
rect 69124 16574 69152 17274
rect 70412 16574 70440 51750
rect 71780 50516 71832 50522
rect 71780 50458 71832 50464
rect 71792 16574 71820 50458
rect 73172 16574 73200 64126
rect 74540 53236 74592 53242
rect 74540 53178 74592 53184
rect 74552 16574 74580 53178
rect 79322 51776 79378 51785
rect 79322 51711 79378 51720
rect 77300 22908 77352 22914
rect 77300 22850 77352 22856
rect 75920 17468 75972 17474
rect 75920 17410 75972 17416
rect 69124 16546 69888 16574
rect 70412 16546 71544 16574
rect 71792 16546 72648 16574
rect 73172 16546 73384 16574
rect 74552 16546 75040 16574
rect 69032 6886 69152 6914
rect 69124 480 69152 6886
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 16546
rect 71516 480 71544 16546
rect 72620 480 72648 16546
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 16546
rect 75012 480 75040 16546
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 75932 354 75960 17410
rect 77312 16574 77340 22850
rect 77312 16546 77432 16574
rect 77404 480 77432 16546
rect 79232 15904 79284 15910
rect 79232 15846 79284 15852
rect 78588 3664 78640 3670
rect 78588 3606 78640 3612
rect 78600 480 78628 3606
rect 76166 354 76278 480
rect 75932 326 76278 354
rect 76166 -960 76278 326
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 15846
rect 79336 3602 79364 51711
rect 80072 16574 80100 71062
rect 84200 58812 84252 58818
rect 84200 58754 84252 58760
rect 82820 29640 82872 29646
rect 82820 29582 82872 29588
rect 81438 26888 81494 26897
rect 81438 26823 81494 26832
rect 81452 16574 81480 26823
rect 82832 16574 82860 29582
rect 80072 16546 80928 16574
rect 81452 16546 81664 16574
rect 82832 16546 83320 16574
rect 79324 3596 79376 3602
rect 79324 3538 79376 3544
rect 80900 480 80928 16546
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 81636 354 81664 16546
rect 83292 480 83320 16546
rect 82054 354 82166 480
rect 81636 326 82166 354
rect 82054 -960 82166 326
rect 83250 -960 83362 480
rect 84212 354 84240 58754
rect 85580 31204 85632 31210
rect 85580 31146 85632 31152
rect 85592 3602 85620 31146
rect 86972 16574 87000 73850
rect 88340 49088 88392 49094
rect 88340 49030 88392 49036
rect 88352 16574 88380 49030
rect 89720 43444 89772 43450
rect 89720 43386 89772 43392
rect 89732 16574 89760 43386
rect 92480 38004 92532 38010
rect 92480 37946 92532 37952
rect 91100 21480 91152 21486
rect 91100 21422 91152 21428
rect 91112 16574 91140 21422
rect 86972 16546 87552 16574
rect 88352 16546 89208 16574
rect 89732 16546 89944 16574
rect 91112 16546 91600 16574
rect 85672 15972 85724 15978
rect 85672 15914 85724 15920
rect 85580 3596 85632 3602
rect 85580 3538 85632 3544
rect 85684 480 85712 15914
rect 86500 3596 86552 3602
rect 86500 3538 86552 3544
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86512 354 86540 3538
rect 86838 354 86950 480
rect 86512 326 86950 354
rect 87524 354 87552 16546
rect 89180 480 89208 16546
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 16546
rect 91572 480 91600 16546
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92492 354 92520 37946
rect 93872 3602 93900 75210
rect 98000 62892 98052 62898
rect 98000 62834 98052 62840
rect 93952 40724 94004 40730
rect 93952 40666 94004 40672
rect 93860 3596 93912 3602
rect 93860 3538 93912 3544
rect 93964 480 93992 40666
rect 95240 32428 95292 32434
rect 95240 32370 95292 32376
rect 95252 16574 95280 32370
rect 96620 24268 96672 24274
rect 96620 24210 96672 24216
rect 96632 16574 96660 24210
rect 98012 16574 98040 62834
rect 99380 47660 99432 47666
rect 99380 47602 99432 47608
rect 99392 16574 99420 47602
rect 100760 31136 100812 31142
rect 100760 31078 100812 31084
rect 95252 16546 95832 16574
rect 96632 16546 97488 16574
rect 98012 16546 98224 16574
rect 99392 16546 99880 16574
rect 94780 3596 94832 3602
rect 94780 3538 94832 3544
rect 92726 354 92838 480
rect 92492 326 92838 354
rect 92726 -960 92838 326
rect 93922 -960 94034 480
rect 94792 354 94820 3538
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95804 354 95832 16546
rect 97460 480 97488 16546
rect 96222 354 96334 480
rect 95804 326 96334 354
rect 95118 -960 95230 326
rect 96222 -960 96334 326
rect 97418 -960 97530 480
rect 98196 354 98224 16546
rect 99852 480 99880 16546
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 31078
rect 102152 16574 102180 76502
rect 121460 73840 121512 73846
rect 121460 73782 121512 73788
rect 107660 72548 107712 72554
rect 107660 72490 107712 72496
rect 104900 68400 104952 68406
rect 104900 68342 104952 68348
rect 104164 18760 104216 18766
rect 104164 18702 104216 18708
rect 102152 16546 102272 16574
rect 102244 480 102272 16546
rect 104176 3670 104204 18702
rect 104912 16574 104940 68342
rect 106278 25528 106334 25537
rect 106278 25463 106334 25472
rect 106292 16574 106320 25463
rect 107672 16574 107700 72490
rect 114560 67040 114612 67046
rect 114560 66982 114612 66988
rect 110420 47592 110472 47598
rect 110420 47534 110472 47540
rect 104912 16546 105768 16574
rect 106292 16546 106504 16574
rect 107672 16546 108160 16574
rect 104532 6248 104584 6254
rect 104532 6190 104584 6196
rect 104164 3664 104216 3670
rect 104164 3606 104216 3612
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103348 480 103376 3538
rect 104544 480 104572 6190
rect 105740 480 105768 16546
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106476 354 106504 16546
rect 108132 480 108160 16546
rect 109316 3664 109368 3670
rect 109316 3606 109368 3612
rect 109328 480 109356 3606
rect 110432 3398 110460 47534
rect 113180 43512 113232 43518
rect 113180 43454 113232 43460
rect 111800 35284 111852 35290
rect 111800 35226 111852 35232
rect 110512 29708 110564 29714
rect 110512 29650 110564 29656
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 29650
rect 111812 16574 111840 35226
rect 113192 16574 113220 43454
rect 114572 16574 114600 66982
rect 118700 61464 118752 61470
rect 118700 61406 118752 61412
rect 115940 46368 115992 46374
rect 115940 46310 115992 46316
rect 115952 16574 115980 46310
rect 117320 39432 117372 39438
rect 117320 39374 117372 39380
rect 111812 16546 112392 16574
rect 113192 16546 114048 16574
rect 114572 16546 114784 16574
rect 115952 16546 116440 16574
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 106894 354 107006 480
rect 106476 326 107006 354
rect 106894 -960 107006 326
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 16546
rect 114020 480 114048 16546
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 16546
rect 116412 480 116440 16546
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117332 354 117360 39374
rect 118712 3398 118740 61406
rect 120080 40792 120132 40798
rect 120080 40734 120132 40740
rect 118792 32496 118844 32502
rect 118792 32438 118844 32444
rect 118700 3392 118752 3398
rect 118700 3334 118752 3340
rect 118804 480 118832 32438
rect 120092 16574 120120 40734
rect 121472 16574 121500 73782
rect 122840 56024 122892 56030
rect 122840 55966 122892 55972
rect 122852 16574 122880 55966
rect 124220 54528 124272 54534
rect 124220 54470 124272 54476
rect 124232 16574 124260 54470
rect 128372 16574 128400 77930
rect 132500 40860 132552 40866
rect 132500 40802 132552 40808
rect 132512 16574 132540 40802
rect 120092 16546 120672 16574
rect 121472 16546 122328 16574
rect 122852 16546 123064 16574
rect 124232 16546 124720 16574
rect 128372 16546 128952 16574
rect 132512 16546 133000 16574
rect 119896 3392 119948 3398
rect 119896 3334 119948 3340
rect 119908 480 119936 3334
rect 117566 354 117678 480
rect 117332 326 117678 354
rect 117566 -960 117678 326
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120644 354 120672 16546
rect 122300 480 122328 16546
rect 121062 354 121174 480
rect 120644 326 121174 354
rect 121062 -960 121174 326
rect 122258 -960 122370 480
rect 123036 354 123064 16546
rect 124692 480 124720 16546
rect 125876 3732 125928 3738
rect 125876 3674 125928 3680
rect 125888 480 125916 3674
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 128924 354 128952 16546
rect 132972 480 133000 16546
rect 164424 14476 164476 14482
rect 164424 14418 164476 14424
rect 136456 6316 136508 6322
rect 136456 6258 136508 6264
rect 136468 480 136496 6258
rect 150624 3528 150676 3534
rect 150624 3470 150676 3476
rect 150636 480 150664 3470
rect 129342 354 129454 480
rect 128924 326 129454 354
rect 129342 -960 129454 326
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 14418
rect 164896 3738 164924 95095
rect 165264 93906 165292 97990
rect 165252 93900 165304 93906
rect 165252 93842 165304 93848
rect 166276 83842 166304 144910
rect 167736 144220 167788 144226
rect 167736 144162 167788 144168
rect 167644 142180 167696 142186
rect 167644 142122 167696 142128
rect 166356 139460 166408 139466
rect 166356 139402 166408 139408
rect 166264 83836 166316 83842
rect 166264 83778 166316 83784
rect 166368 82482 166396 139402
rect 166448 121508 166500 121514
rect 166448 121450 166500 121456
rect 166460 93362 166488 121450
rect 166540 110492 166592 110498
rect 166540 110434 166592 110440
rect 166448 93356 166500 93362
rect 166448 93298 166500 93304
rect 166552 86766 166580 110434
rect 167656 93945 167684 142122
rect 167748 110129 167776 144162
rect 170404 138032 170456 138038
rect 170404 137974 170456 137980
rect 169116 125656 169168 125662
rect 169116 125598 169168 125604
rect 169024 120148 169076 120154
rect 169024 120090 169076 120096
rect 167920 111784 167972 111790
rect 167918 111752 167920 111761
rect 167972 111752 167974 111761
rect 167918 111687 167974 111696
rect 167734 110120 167790 110129
rect 167734 110055 167790 110064
rect 167828 109064 167880 109070
rect 167828 109006 167880 109012
rect 167736 99408 167788 99414
rect 167736 99350 167788 99356
rect 167642 93936 167698 93945
rect 167642 93871 167698 93880
rect 166540 86760 166592 86766
rect 166540 86702 166592 86708
rect 167748 85542 167776 99350
rect 167736 85536 167788 85542
rect 167736 85478 167788 85484
rect 166356 82476 166408 82482
rect 166356 82418 166408 82424
rect 167840 81190 167868 109006
rect 168104 108996 168156 109002
rect 168104 108938 168156 108944
rect 168116 108769 168144 108938
rect 168102 108760 168158 108769
rect 168102 108695 168158 108704
rect 168288 95940 168340 95946
rect 168288 95882 168340 95888
rect 168300 92138 168328 95882
rect 168288 92132 168340 92138
rect 168288 92074 168340 92080
rect 169036 86630 169064 120090
rect 169128 94042 169156 125598
rect 169208 107704 169260 107710
rect 169208 107646 169260 107652
rect 169116 94036 169168 94042
rect 169116 93978 169168 93984
rect 169220 89622 169248 107646
rect 169300 98660 169352 98666
rect 169300 98602 169352 98608
rect 169312 92274 169340 98602
rect 169300 92268 169352 92274
rect 169300 92210 169352 92216
rect 169208 89616 169260 89622
rect 169208 89558 169260 89564
rect 169024 86624 169076 86630
rect 169024 86566 169076 86572
rect 170416 82550 170444 137974
rect 170496 122868 170548 122874
rect 170496 122810 170548 122816
rect 170508 90846 170536 122810
rect 170588 118856 170640 118862
rect 170588 118798 170640 118804
rect 170496 90840 170548 90846
rect 170496 90782 170548 90788
rect 170600 87990 170628 118798
rect 170680 106344 170732 106350
rect 170680 106286 170732 106292
rect 170588 87984 170640 87990
rect 170588 87926 170640 87932
rect 170692 83978 170720 106286
rect 171796 90710 171824 146270
rect 171968 132524 172020 132530
rect 171968 132466 172020 132472
rect 171876 124228 171928 124234
rect 171876 124170 171928 124176
rect 171784 90704 171836 90710
rect 171784 90646 171836 90652
rect 171784 89004 171836 89010
rect 171784 88946 171836 88952
rect 170680 83972 170732 83978
rect 170680 83914 170732 83920
rect 170404 82544 170456 82550
rect 170404 82486 170456 82492
rect 167828 81184 167880 81190
rect 167828 81126 167880 81132
rect 164884 3732 164936 3738
rect 164884 3674 164936 3680
rect 171796 3670 171824 88946
rect 171888 77178 171916 124170
rect 171980 88126 172008 132466
rect 172060 104916 172112 104922
rect 172060 104858 172112 104864
rect 172072 89690 172100 104858
rect 173176 93430 173204 153206
rect 173348 129804 173400 129810
rect 173348 129746 173400 129752
rect 173256 127016 173308 127022
rect 173256 126958 173308 126964
rect 173164 93424 173216 93430
rect 173164 93366 173216 93372
rect 172060 89684 172112 89690
rect 172060 89626 172112 89632
rect 171968 88120 172020 88126
rect 171968 88062 172020 88068
rect 173268 79762 173296 126958
rect 173360 89554 173388 129746
rect 173440 117360 173492 117366
rect 173440 117302 173492 117308
rect 173348 89548 173400 89554
rect 173348 89490 173400 89496
rect 173452 85270 173480 117302
rect 173440 85264 173492 85270
rect 173440 85206 173492 85212
rect 173256 79756 173308 79762
rect 173256 79698 173308 79704
rect 171876 77172 171928 77178
rect 171876 77114 171928 77120
rect 174556 6866 174584 337311
rect 174648 322250 174676 369990
rect 176108 366036 176160 366042
rect 176108 365978 176160 365984
rect 175924 362296 175976 362302
rect 175924 362238 175976 362244
rect 174636 322244 174688 322250
rect 174636 322186 174688 322192
rect 175188 314696 175240 314702
rect 175188 314638 175240 314644
rect 175096 301504 175148 301510
rect 175096 301446 175148 301452
rect 175108 300966 175136 301446
rect 175096 300960 175148 300966
rect 175096 300902 175148 300908
rect 175108 215966 175136 300902
rect 175096 215960 175148 215966
rect 175096 215902 175148 215908
rect 175200 181393 175228 314638
rect 175186 181384 175242 181393
rect 175186 181319 175242 181328
rect 174636 140072 174688 140078
rect 174636 140014 174688 140020
rect 174648 92206 174676 140014
rect 174728 111852 174780 111858
rect 174728 111794 174780 111800
rect 174636 92200 174688 92206
rect 174636 92142 174688 92148
rect 174740 85338 174768 111794
rect 174820 109132 174872 109138
rect 174820 109074 174872 109080
rect 174728 85332 174780 85338
rect 174728 85274 174780 85280
rect 174832 84046 174860 109074
rect 175936 87718 175964 362238
rect 176016 314016 176068 314022
rect 176016 313958 176068 313964
rect 176028 213450 176056 313958
rect 176120 311166 176148 365978
rect 176108 311160 176160 311166
rect 176108 311102 176160 311108
rect 176660 267028 176712 267034
rect 176660 266970 176712 266976
rect 176672 266422 176700 266970
rect 176660 266416 176712 266422
rect 176660 266358 176712 266364
rect 176108 255332 176160 255338
rect 176108 255274 176160 255280
rect 176120 233102 176148 255274
rect 176200 248464 176252 248470
rect 176200 248406 176252 248412
rect 176108 233096 176160 233102
rect 176212 233073 176240 248406
rect 176108 233038 176160 233044
rect 176198 233064 176254 233073
rect 176016 213444 176068 213450
rect 176016 213386 176068 213392
rect 176120 192574 176148 233038
rect 176198 232999 176254 233008
rect 176108 192568 176160 192574
rect 176108 192510 176160 192516
rect 176016 129872 176068 129878
rect 176016 129814 176068 129820
rect 175924 87712 175976 87718
rect 175924 87654 175976 87660
rect 174820 84040 174872 84046
rect 174820 83982 174872 83988
rect 176028 82686 176056 129814
rect 176200 110560 176252 110566
rect 176200 110502 176252 110508
rect 176108 106412 176160 106418
rect 176108 106354 176160 106360
rect 176016 82680 176068 82686
rect 176016 82622 176068 82628
rect 176120 79966 176148 106354
rect 176212 93158 176240 110502
rect 176200 93152 176252 93158
rect 176200 93094 176252 93100
rect 177316 86358 177344 387903
rect 184204 387874 184256 387880
rect 181444 381540 181496 381546
rect 181444 381482 181496 381488
rect 178684 351212 178736 351218
rect 178684 351154 178736 351160
rect 177948 319524 178000 319530
rect 177948 319466 178000 319472
rect 177960 318850 177988 319466
rect 177948 318844 178000 318850
rect 177948 318786 178000 318792
rect 177396 291848 177448 291854
rect 177396 291790 177448 291796
rect 177408 223038 177436 291790
rect 177856 266416 177908 266422
rect 177856 266358 177908 266364
rect 177396 223032 177448 223038
rect 177396 222974 177448 222980
rect 177868 217326 177896 266358
rect 177856 217320 177908 217326
rect 177856 217262 177908 217268
rect 177960 185774 177988 318786
rect 177948 185768 178000 185774
rect 177948 185710 178000 185716
rect 177396 178084 177448 178090
rect 177396 178026 177448 178032
rect 177408 155854 177436 178026
rect 177396 155848 177448 155854
rect 177396 155790 177448 155796
rect 177396 133952 177448 133958
rect 177396 133894 177448 133900
rect 177304 86352 177356 86358
rect 177304 86294 177356 86300
rect 176108 79960 176160 79966
rect 176108 79902 176160 79908
rect 177408 78538 177436 133894
rect 177488 128376 177540 128382
rect 177488 128318 177540 128324
rect 177500 79830 177528 128318
rect 177488 79824 177540 79830
rect 177488 79766 177540 79772
rect 177396 78532 177448 78538
rect 177396 78474 177448 78480
rect 178696 69834 178724 351154
rect 180064 346520 180116 346526
rect 180064 346462 180116 346468
rect 179328 346452 179380 346458
rect 179328 346394 179380 346400
rect 179236 290012 179288 290018
rect 179236 289954 179288 289960
rect 178776 262880 178828 262886
rect 178776 262822 178828 262828
rect 178788 255406 178816 262822
rect 178776 255400 178828 255406
rect 178776 255342 178828 255348
rect 179248 210458 179276 289954
rect 179236 210452 179288 210458
rect 179236 210394 179288 210400
rect 179340 209710 179368 346394
rect 179420 283620 179472 283626
rect 179420 283562 179472 283568
rect 179432 282946 179460 283562
rect 179420 282940 179472 282946
rect 179420 282882 179472 282888
rect 179880 259480 179932 259486
rect 179880 259422 179932 259428
rect 179892 255338 179920 259422
rect 179880 255332 179932 255338
rect 179880 255274 179932 255280
rect 179328 209704 179380 209710
rect 179328 209646 179380 209652
rect 179340 209234 179368 209646
rect 179328 209228 179380 209234
rect 179328 209170 179380 209176
rect 178776 140820 178828 140826
rect 178776 140762 178828 140768
rect 178788 86698 178816 140762
rect 178868 118788 178920 118794
rect 178868 118730 178920 118736
rect 178880 93974 178908 118730
rect 178868 93968 178920 93974
rect 178868 93910 178920 93916
rect 178776 86692 178828 86698
rect 178776 86634 178828 86640
rect 178684 69828 178736 69834
rect 178684 69770 178736 69776
rect 174544 6860 174596 6866
rect 174544 6802 174596 6808
rect 180076 4962 180104 346462
rect 180156 345704 180208 345710
rect 180156 345646 180208 345652
rect 180168 77994 180196 345646
rect 180708 282940 180760 282946
rect 180708 282882 180760 282888
rect 180616 255400 180668 255406
rect 180616 255342 180668 255348
rect 180248 183660 180300 183666
rect 180248 183602 180300 183608
rect 180260 171018 180288 183602
rect 180628 181490 180656 255342
rect 180720 206310 180748 282882
rect 180708 206304 180760 206310
rect 180708 206246 180760 206252
rect 180616 181484 180668 181490
rect 180616 181426 180668 181432
rect 180248 171012 180300 171018
rect 180248 170954 180300 170960
rect 180248 145580 180300 145586
rect 180248 145522 180300 145528
rect 180260 109002 180288 145522
rect 180340 124296 180392 124302
rect 180340 124238 180392 124244
rect 180248 108996 180300 109002
rect 180248 108938 180300 108944
rect 180352 89418 180380 124238
rect 180432 107772 180484 107778
rect 180432 107714 180484 107720
rect 180340 89412 180392 89418
rect 180340 89354 180392 89360
rect 180444 78606 180472 107714
rect 180432 78600 180484 78606
rect 180432 78542 180484 78548
rect 180156 77988 180208 77994
rect 180156 77930 180208 77936
rect 181456 8294 181484 381482
rect 182916 367260 182968 367266
rect 182916 367202 182968 367208
rect 181536 364676 181588 364682
rect 181536 364618 181588 364624
rect 181548 319462 181576 364618
rect 182824 355360 182876 355366
rect 182824 355302 182876 355308
rect 181536 319456 181588 319462
rect 181536 319398 181588 319404
rect 181536 316056 181588 316062
rect 181536 315998 181588 316004
rect 181548 198286 181576 315998
rect 182180 306400 182232 306406
rect 182180 306342 182232 306348
rect 182192 300830 182220 306342
rect 182180 300824 182232 300830
rect 182180 300766 182232 300772
rect 182088 285796 182140 285802
rect 182088 285738 182140 285744
rect 181628 268456 181680 268462
rect 181628 268398 181680 268404
rect 181640 237114 181668 268398
rect 181628 237108 181680 237114
rect 181628 237050 181680 237056
rect 182100 222018 182128 285738
rect 182088 222012 182140 222018
rect 182088 221954 182140 221960
rect 182100 221542 182128 221954
rect 182088 221536 182140 221542
rect 182088 221478 182140 221484
rect 181536 198280 181588 198286
rect 181536 198222 181588 198228
rect 181536 136672 181588 136678
rect 181536 136614 181588 136620
rect 181548 83910 181576 136614
rect 181628 116000 181680 116006
rect 181628 115942 181680 115948
rect 181536 83904 181588 83910
rect 181536 83846 181588 83852
rect 181640 81258 181668 115942
rect 181628 81252 181680 81258
rect 181628 81194 181680 81200
rect 182836 45558 182864 355302
rect 182928 330682 182956 367202
rect 182916 330676 182968 330682
rect 182916 330618 182968 330624
rect 183468 300824 183520 300830
rect 183468 300766 183520 300772
rect 183480 300150 183508 300766
rect 183468 300144 183520 300150
rect 183468 300086 183520 300092
rect 182916 296744 182968 296750
rect 182916 296686 182968 296692
rect 182928 231538 182956 296686
rect 183376 268388 183428 268394
rect 183376 268330 183428 268336
rect 183388 267850 183416 268330
rect 183376 267844 183428 267850
rect 183376 267786 183428 267792
rect 183388 232626 183416 267786
rect 183376 232620 183428 232626
rect 183376 232562 183428 232568
rect 182916 231532 182968 231538
rect 182916 231474 182968 231480
rect 183480 189786 183508 300086
rect 183468 189780 183520 189786
rect 183468 189722 183520 189728
rect 182914 181656 182970 181665
rect 182914 181591 182970 181600
rect 182928 93158 182956 181591
rect 183008 120216 183060 120222
rect 183008 120158 183060 120164
rect 182916 93152 182968 93158
rect 182916 93094 182968 93100
rect 183020 82618 183048 120158
rect 183008 82612 183060 82618
rect 183008 82554 183060 82560
rect 184216 80714 184244 387874
rect 209780 382288 209832 382294
rect 209780 382230 209832 382236
rect 189724 380180 189776 380186
rect 189724 380122 189776 380128
rect 185584 373312 185636 373318
rect 185584 373254 185636 373260
rect 184848 361684 184900 361690
rect 184848 361626 184900 361632
rect 184296 299668 184348 299674
rect 184296 299610 184348 299616
rect 184308 211954 184336 299610
rect 184756 281648 184808 281654
rect 184756 281590 184808 281596
rect 184388 243024 184440 243030
rect 184388 242966 184440 242972
rect 184400 238513 184428 242966
rect 184386 238504 184442 238513
rect 184386 238439 184442 238448
rect 184768 214742 184796 281590
rect 184860 278730 184888 361626
rect 184848 278724 184900 278730
rect 184848 278666 184900 278672
rect 184860 278254 184888 278666
rect 184848 278248 184900 278254
rect 184848 278190 184900 278196
rect 184756 214736 184808 214742
rect 184756 214678 184808 214684
rect 184296 211948 184348 211954
rect 184296 211890 184348 211896
rect 184296 196784 184348 196790
rect 184296 196726 184348 196732
rect 184308 96014 184336 196726
rect 184388 127084 184440 127090
rect 184388 127026 184440 127032
rect 184296 96008 184348 96014
rect 184296 95950 184348 95956
rect 184400 81394 184428 127026
rect 184388 81388 184440 81394
rect 184388 81330 184440 81336
rect 184204 80708 184256 80714
rect 184204 80650 184256 80656
rect 182824 45552 182876 45558
rect 182824 45494 182876 45500
rect 185596 39506 185624 373254
rect 187056 363248 187108 363254
rect 187056 363190 187108 363196
rect 186964 356788 187016 356794
rect 186964 356730 187016 356736
rect 185676 337408 185728 337414
rect 185676 337350 185728 337356
rect 185688 83502 185716 337350
rect 185768 289128 185820 289134
rect 185768 289070 185820 289076
rect 185780 235278 185808 289070
rect 185860 242956 185912 242962
rect 185860 242898 185912 242904
rect 185768 235272 185820 235278
rect 185768 235214 185820 235220
rect 185872 228886 185900 242898
rect 185860 228880 185912 228886
rect 185860 228822 185912 228828
rect 185676 83496 185728 83502
rect 185676 83438 185728 83444
rect 185584 39500 185636 39506
rect 185584 39442 185636 39448
rect 186976 9654 187004 356730
rect 187068 289814 187096 363190
rect 188344 344344 188396 344350
rect 188344 344286 188396 344292
rect 187240 303680 187292 303686
rect 187240 303622 187292 303628
rect 187252 298178 187280 303622
rect 187240 298172 187292 298178
rect 187240 298114 187292 298120
rect 187056 289808 187108 289814
rect 187056 289750 187108 289756
rect 187056 278248 187108 278254
rect 187056 278190 187108 278196
rect 187068 180266 187096 278190
rect 187148 274712 187200 274718
rect 187148 274654 187200 274660
rect 187160 271930 187188 274654
rect 187148 271924 187200 271930
rect 187148 271866 187200 271872
rect 187056 180260 187108 180266
rect 187056 180202 187108 180208
rect 187160 180198 187188 271866
rect 187252 239494 187280 298114
rect 187240 239488 187292 239494
rect 187240 239430 187292 239436
rect 187148 180192 187200 180198
rect 187148 180134 187200 180140
rect 187054 177440 187110 177449
rect 187054 177375 187110 177384
rect 187068 82249 187096 177375
rect 187054 82240 187110 82249
rect 187054 82175 187110 82184
rect 188356 64326 188384 344286
rect 188528 332580 188580 332586
rect 188528 332522 188580 332528
rect 188540 331265 188568 332522
rect 188526 331256 188582 331265
rect 188526 331191 188582 331200
rect 188436 295520 188488 295526
rect 188436 295462 188488 295468
rect 188448 192778 188476 295462
rect 188528 291236 188580 291242
rect 188528 291178 188580 291184
rect 188540 229974 188568 291178
rect 188620 251252 188672 251258
rect 188620 251194 188672 251200
rect 188632 233918 188660 251194
rect 188620 233912 188672 233918
rect 188620 233854 188672 233860
rect 188528 229968 188580 229974
rect 188528 229910 188580 229916
rect 188436 192772 188488 192778
rect 188436 192714 188488 192720
rect 188434 184240 188490 184249
rect 188434 184175 188490 184184
rect 188448 78062 188476 184175
rect 188526 82104 188582 82113
rect 188526 82039 188582 82048
rect 188436 78056 188488 78062
rect 188436 77998 188488 78004
rect 188344 64320 188396 64326
rect 188344 64262 188396 64268
rect 186964 9648 187016 9654
rect 186964 9590 187016 9596
rect 181444 8288 181496 8294
rect 181444 8230 181496 8236
rect 180064 4956 180116 4962
rect 180064 4898 180116 4904
rect 171784 3664 171836 3670
rect 171784 3606 171836 3612
rect 171966 3496 172022 3505
rect 188540 3466 188568 82039
rect 189736 47734 189764 380122
rect 209042 379536 209098 379545
rect 209042 379471 209098 379480
rect 198004 372632 198056 372638
rect 198004 372574 198056 372580
rect 194048 368756 194100 368762
rect 194048 368698 194100 368704
rect 189816 366104 189868 366110
rect 189816 366046 189868 366052
rect 189828 323610 189856 366046
rect 191104 363180 191156 363186
rect 191104 363122 191156 363128
rect 190460 340944 190512 340950
rect 190460 340886 190512 340892
rect 189816 323604 189868 323610
rect 189816 323546 189868 323552
rect 190368 310548 190420 310554
rect 190368 310490 190420 310496
rect 189816 292596 189868 292602
rect 189816 292538 189868 292544
rect 189828 249082 189856 292538
rect 190276 260908 190328 260914
rect 190276 260850 190328 260856
rect 189816 249076 189868 249082
rect 189816 249018 189868 249024
rect 189816 242208 189868 242214
rect 189816 242150 189868 242156
rect 189828 233102 189856 242150
rect 189816 233096 189868 233102
rect 189816 233038 189868 233044
rect 190184 231124 190236 231130
rect 190184 231066 190236 231072
rect 190196 227118 190224 231066
rect 190184 227112 190236 227118
rect 190184 227054 190236 227060
rect 190288 213246 190316 260850
rect 190276 213240 190328 213246
rect 190276 213182 190328 213188
rect 189816 187196 189868 187202
rect 189816 187138 189868 187144
rect 189828 90370 189856 187138
rect 190380 177478 190408 310490
rect 190472 281654 190500 340886
rect 191116 330546 191144 363122
rect 192484 363044 192536 363050
rect 192484 362986 192536 362992
rect 191104 330540 191156 330546
rect 191104 330482 191156 330488
rect 191104 320884 191156 320890
rect 191104 320826 191156 320832
rect 190460 281648 190512 281654
rect 190460 281590 190512 281596
rect 190368 177472 190420 177478
rect 190368 177414 190420 177420
rect 189816 90364 189868 90370
rect 189816 90306 189868 90312
rect 189724 47728 189776 47734
rect 189724 47670 189776 47676
rect 191116 4146 191144 320826
rect 191748 281648 191800 281654
rect 191748 281590 191800 281596
rect 191760 281450 191788 281590
rect 192496 281518 192524 362986
rect 193956 358964 194008 358970
rect 193956 358906 194008 358912
rect 193864 342916 193916 342922
rect 193864 342858 193916 342864
rect 193128 302252 193180 302258
rect 193128 302194 193180 302200
rect 193036 297220 193088 297226
rect 193036 297162 193088 297168
rect 192484 281512 192536 281518
rect 192484 281454 192536 281460
rect 191748 281444 191800 281450
rect 191748 281386 191800 281392
rect 192484 278792 192536 278798
rect 192484 278734 192536 278740
rect 191748 275460 191800 275466
rect 191748 275402 191800 275408
rect 191196 267776 191248 267782
rect 191196 267718 191248 267724
rect 191208 235686 191236 267718
rect 191288 252612 191340 252618
rect 191288 252554 191340 252560
rect 191196 235680 191248 235686
rect 191196 235622 191248 235628
rect 191300 231130 191328 252554
rect 191288 231124 191340 231130
rect 191288 231066 191340 231072
rect 191760 216714 191788 275402
rect 192496 231130 192524 278734
rect 192944 246356 192996 246362
rect 192944 246298 192996 246304
rect 192484 231124 192536 231130
rect 192484 231066 192536 231072
rect 192956 221474 192984 246298
rect 193048 239562 193076 297162
rect 193036 239556 193088 239562
rect 193036 239498 193088 239504
rect 192944 221468 192996 221474
rect 192944 221410 192996 221416
rect 191748 216708 191800 216714
rect 191748 216650 191800 216656
rect 193140 189990 193168 302194
rect 193128 189984 193180 189990
rect 193128 189926 193180 189932
rect 192484 125724 192536 125730
rect 192484 125666 192536 125672
rect 192496 89486 192524 125666
rect 192576 104984 192628 104990
rect 192576 104926 192628 104932
rect 192588 93809 192616 104926
rect 192574 93800 192630 93809
rect 192574 93735 192630 93744
rect 192484 89480 192536 89486
rect 192484 89422 192536 89428
rect 193876 65686 193904 342858
rect 193968 285666 193996 358906
rect 194060 339454 194088 368698
rect 196808 364744 196860 364750
rect 196808 364686 196860 364692
rect 195428 364608 195480 364614
rect 195428 364550 195480 364556
rect 195336 363112 195388 363118
rect 195336 363054 195388 363060
rect 195242 360360 195298 360369
rect 195242 360295 195298 360304
rect 194048 339448 194100 339454
rect 194048 339390 194100 339396
rect 195060 336796 195112 336802
rect 195060 336738 195112 336744
rect 195072 335238 195100 336738
rect 195060 335232 195112 335238
rect 195060 335174 195112 335180
rect 195256 310486 195284 360295
rect 195244 310480 195296 310486
rect 195244 310422 195296 310428
rect 195244 309120 195296 309126
rect 195244 309062 195296 309068
rect 195256 307834 195284 309062
rect 195244 307828 195296 307834
rect 195244 307770 195296 307776
rect 194048 292596 194100 292602
rect 194048 292538 194100 292544
rect 193956 285660 194008 285666
rect 193956 285602 194008 285608
rect 194060 255270 194088 292538
rect 194508 273284 194560 273290
rect 194508 273226 194560 273232
rect 194048 255264 194100 255270
rect 194048 255206 194100 255212
rect 194416 249076 194468 249082
rect 194416 249018 194468 249024
rect 194428 248810 194456 249018
rect 194416 248804 194468 248810
rect 194416 248746 194468 248752
rect 194324 240780 194376 240786
rect 194324 240722 194376 240728
rect 194336 238202 194364 240722
rect 194324 238196 194376 238202
rect 194324 238138 194376 238144
rect 194428 225826 194456 248746
rect 194416 225820 194468 225826
rect 194416 225762 194468 225768
rect 194520 195498 194548 273226
rect 195152 239420 195204 239426
rect 195152 239362 195204 239368
rect 195164 237046 195192 239362
rect 195152 237040 195204 237046
rect 195152 236982 195204 236988
rect 194508 195492 194560 195498
rect 194508 195434 194560 195440
rect 195256 182986 195284 307770
rect 195348 294642 195376 363054
rect 195440 326398 195468 364550
rect 196624 362296 196676 362302
rect 196624 362238 196676 362244
rect 195520 327140 195572 327146
rect 195520 327082 195572 327088
rect 195428 326392 195480 326398
rect 195428 326334 195480 326340
rect 195428 312656 195480 312662
rect 195428 312598 195480 312604
rect 195336 294636 195388 294642
rect 195336 294578 195388 294584
rect 195440 277394 195468 312598
rect 195532 309126 195560 327082
rect 195520 309120 195572 309126
rect 195520 309062 195572 309068
rect 196636 302938 196664 362238
rect 196716 360392 196768 360398
rect 196716 360334 196768 360340
rect 196728 338026 196756 360334
rect 196820 354006 196848 364686
rect 198016 357474 198044 372574
rect 209056 366042 209084 379471
rect 209792 374066 209820 382230
rect 213184 378208 213236 378214
rect 213184 378150 213236 378156
rect 209780 374060 209832 374066
rect 209780 374002 209832 374008
rect 209044 366036 209096 366042
rect 209044 365978 209096 365984
rect 206466 365800 206522 365809
rect 206466 365735 206522 365744
rect 198648 364404 198700 364410
rect 198648 364346 198700 364352
rect 198186 360224 198242 360233
rect 198186 360159 198242 360168
rect 198094 358320 198150 358329
rect 198094 358255 198150 358264
rect 198004 357468 198056 357474
rect 198004 357410 198056 357416
rect 196808 354000 196860 354006
rect 196808 353942 196860 353948
rect 198016 353705 198044 357410
rect 198002 353696 198058 353705
rect 198002 353631 198058 353640
rect 197360 350600 197412 350606
rect 197360 350542 197412 350548
rect 197372 349625 197400 350542
rect 197358 349616 197414 349625
rect 197358 349551 197414 349560
rect 197358 347440 197414 347449
rect 197358 347375 197414 347384
rect 197372 346458 197400 347375
rect 197360 346452 197412 346458
rect 197360 346394 197412 346400
rect 198002 342680 198058 342689
rect 198002 342615 198058 342624
rect 197358 340640 197414 340649
rect 197358 340575 197414 340584
rect 197372 339522 197400 340575
rect 197360 339516 197412 339522
rect 197360 339458 197412 339464
rect 196716 338020 196768 338026
rect 196716 337962 196768 337968
rect 197358 337920 197414 337929
rect 197358 337855 197414 337864
rect 197372 336802 197400 337855
rect 197360 336796 197412 336802
rect 197360 336738 197412 336744
rect 197358 335880 197414 335889
rect 197358 335815 197414 335824
rect 197372 335374 197400 335815
rect 197360 335368 197412 335374
rect 197360 335310 197412 335316
rect 197358 331800 197414 331809
rect 197358 331735 197414 331744
rect 197372 331294 197400 331735
rect 197360 331288 197412 331294
rect 197360 331230 197412 331236
rect 197358 329080 197414 329089
rect 197358 329015 197414 329024
rect 197372 328506 197400 329015
rect 197360 328500 197412 328506
rect 197360 328442 197412 328448
rect 197358 327176 197414 327185
rect 197358 327111 197360 327120
rect 197412 327111 197414 327120
rect 197360 327082 197412 327088
rect 197360 322924 197412 322930
rect 197360 322866 197412 322872
rect 197372 322425 197400 322866
rect 197358 322416 197414 322425
rect 197358 322351 197414 322360
rect 197358 320240 197414 320249
rect 197358 320175 197360 320184
rect 197412 320175 197414 320184
rect 197360 320146 197412 320152
rect 197176 317484 197228 317490
rect 197176 317426 197228 317432
rect 196806 309360 196862 309369
rect 196806 309295 196862 309304
rect 196820 306374 196848 309295
rect 196728 306346 196848 306374
rect 196624 302932 196676 302938
rect 196624 302874 196676 302880
rect 196728 301594 196756 306346
rect 196636 301566 196756 301594
rect 196636 295730 196664 301566
rect 196716 298240 196768 298246
rect 196716 298182 196768 298188
rect 196624 295724 196676 295730
rect 196624 295666 196676 295672
rect 195888 295452 195940 295458
rect 195888 295394 195940 295400
rect 195796 277500 195848 277506
rect 195796 277442 195848 277448
rect 195808 277394 195836 277442
rect 195440 277366 195836 277394
rect 195704 264240 195756 264246
rect 195704 264182 195756 264188
rect 195716 235958 195744 264182
rect 195704 235952 195756 235958
rect 195704 235894 195756 235900
rect 195808 222902 195836 277366
rect 195900 239698 195928 295394
rect 195888 239692 195940 239698
rect 195888 239634 195940 239640
rect 196636 229906 196664 295666
rect 196728 234054 196756 298182
rect 196808 285728 196860 285734
rect 196808 285670 196860 285676
rect 196820 242554 196848 285670
rect 196808 242548 196860 242554
rect 196808 242490 196860 242496
rect 196808 239488 196860 239494
rect 197188 239465 197216 317426
rect 197358 315480 197414 315489
rect 197358 315415 197414 315424
rect 197372 314702 197400 315415
rect 197360 314696 197412 314702
rect 197360 314638 197412 314644
rect 197358 313440 197414 313449
rect 197358 313375 197414 313384
rect 197372 313342 197400 313375
rect 197360 313336 197412 313342
rect 197360 313278 197412 313284
rect 197358 311400 197414 311409
rect 197358 311335 197414 311344
rect 197372 310554 197400 311335
rect 197360 310548 197412 310554
rect 197360 310490 197412 310496
rect 197266 306640 197322 306649
rect 197266 306575 197322 306584
rect 197280 301510 197308 306575
rect 197358 304600 197414 304609
rect 197358 304535 197414 304544
rect 197372 303686 197400 304535
rect 197360 303680 197412 303686
rect 197360 303622 197412 303628
rect 197358 302560 197414 302569
rect 197358 302495 197414 302504
rect 197372 302258 197400 302495
rect 197360 302252 197412 302258
rect 197360 302194 197412 302200
rect 197268 301504 197320 301510
rect 197268 301446 197320 301452
rect 198016 301345 198044 342615
rect 198108 332586 198136 358255
rect 198200 354686 198228 360159
rect 198660 356726 198688 364346
rect 206480 363254 206508 365735
rect 206468 363248 206520 363254
rect 206468 363190 206520 363196
rect 199384 362364 199436 362370
rect 199384 362306 199436 362312
rect 198832 360256 198884 360262
rect 198832 360198 198884 360204
rect 198844 358086 198872 360198
rect 198832 358080 198884 358086
rect 198832 358022 198884 358028
rect 198280 356720 198332 356726
rect 198280 356662 198332 356668
rect 198648 356720 198700 356726
rect 198648 356662 198700 356668
rect 198292 356425 198320 356662
rect 198278 356416 198334 356425
rect 198278 356351 198334 356360
rect 198188 354680 198240 354686
rect 198188 354622 198240 354628
rect 198278 351520 198334 351529
rect 198278 351455 198334 351464
rect 198186 344720 198242 344729
rect 198186 344655 198242 344664
rect 198096 332580 198148 332586
rect 198096 332522 198148 332528
rect 198094 325000 198150 325009
rect 198094 324935 198150 324944
rect 198108 309194 198136 324935
rect 198200 319530 198228 344655
rect 198292 327962 198320 351455
rect 199014 333840 199070 333849
rect 199014 333775 199070 333784
rect 199028 332654 199056 333775
rect 198832 332648 198884 332654
rect 198832 332590 198884 332596
rect 199016 332648 199068 332654
rect 199016 332590 199068 332596
rect 198280 327956 198332 327962
rect 198280 327898 198332 327904
rect 198188 319524 198240 319530
rect 198188 319466 198240 319472
rect 198646 318200 198702 318209
rect 198646 318135 198702 318144
rect 198660 317490 198688 318135
rect 198648 317484 198700 317490
rect 198648 317426 198700 317432
rect 198096 309188 198148 309194
rect 198096 309130 198148 309136
rect 197450 301336 197506 301345
rect 197450 301271 197506 301280
rect 198002 301336 198058 301345
rect 198002 301271 198058 301280
rect 197464 300937 197492 301271
rect 197450 300928 197506 300937
rect 197450 300863 197506 300872
rect 197360 300144 197412 300150
rect 197360 300086 197412 300092
rect 197372 299985 197400 300086
rect 197358 299976 197414 299985
rect 197358 299911 197414 299920
rect 197358 297800 197414 297809
rect 197358 297735 197414 297744
rect 197372 297226 197400 297735
rect 197360 297220 197412 297226
rect 197360 297162 197412 297168
rect 197464 296714 197492 300863
rect 197372 296686 197492 296714
rect 197372 275466 197400 296686
rect 197450 295760 197506 295769
rect 197450 295695 197506 295704
rect 197464 295458 197492 295695
rect 197452 295452 197504 295458
rect 197452 295394 197504 295400
rect 197450 293720 197506 293729
rect 197450 293655 197506 293664
rect 197464 292602 197492 293655
rect 197452 292596 197504 292602
rect 197452 292538 197504 292544
rect 197450 291000 197506 291009
rect 197450 290935 197506 290944
rect 197464 289882 197492 290935
rect 197452 289876 197504 289882
rect 197452 289818 197504 289824
rect 197450 288960 197506 288969
rect 197450 288895 197506 288904
rect 197464 288454 197492 288895
rect 197452 288448 197504 288454
rect 197452 288390 197504 288396
rect 197450 286920 197506 286929
rect 197450 286855 197506 286864
rect 197464 285802 197492 286855
rect 197452 285796 197504 285802
rect 197452 285738 197504 285744
rect 197450 284200 197506 284209
rect 197450 284135 197506 284144
rect 197464 282946 197492 284135
rect 197452 282940 197504 282946
rect 197452 282882 197504 282888
rect 197450 282160 197506 282169
rect 197450 282095 197506 282104
rect 197464 281586 197492 282095
rect 197452 281580 197504 281586
rect 197452 281522 197504 281528
rect 197452 281444 197504 281450
rect 197452 281386 197504 281392
rect 197464 280265 197492 281386
rect 197450 280256 197506 280265
rect 197450 280191 197506 280200
rect 197450 277536 197506 277545
rect 197450 277471 197452 277480
rect 197504 277471 197506 277480
rect 197452 277442 197504 277448
rect 197360 275460 197412 275466
rect 197360 275402 197412 275408
rect 197358 275360 197414 275369
rect 197358 275295 197414 275304
rect 197372 274718 197400 275295
rect 197360 274712 197412 274718
rect 197360 274654 197412 274660
rect 197358 273320 197414 273329
rect 197358 273255 197360 273264
rect 197412 273255 197414 273264
rect 197360 273226 197412 273232
rect 197358 271280 197414 271289
rect 197358 271215 197414 271224
rect 197372 271182 197400 271215
rect 197360 271176 197412 271182
rect 197360 271118 197412 271124
rect 197358 268560 197414 268569
rect 197358 268495 197414 268504
rect 197372 267850 197400 268495
rect 197360 267844 197412 267850
rect 197360 267786 197412 267792
rect 197358 266520 197414 266529
rect 197358 266455 197414 266464
rect 197372 266422 197400 266455
rect 197360 266416 197412 266422
rect 197360 266358 197412 266364
rect 197358 264480 197414 264489
rect 197358 264415 197414 264424
rect 197372 264246 197400 264415
rect 197360 264240 197412 264246
rect 197360 264182 197412 264188
rect 197358 261760 197414 261769
rect 197358 261695 197414 261704
rect 197372 260914 197400 261695
rect 197360 260908 197412 260914
rect 197360 260850 197412 260856
rect 197358 259720 197414 259729
rect 197358 259655 197414 259664
rect 197372 259486 197400 259655
rect 197360 259480 197412 259486
rect 197360 259422 197412 259428
rect 197358 257680 197414 257689
rect 197358 257615 197414 257624
rect 197372 257378 197400 257615
rect 197360 257372 197412 257378
rect 197360 257314 197412 257320
rect 197358 255640 197414 255649
rect 197358 255575 197414 255584
rect 197372 255338 197400 255575
rect 197360 255332 197412 255338
rect 197360 255274 197412 255280
rect 197358 252920 197414 252929
rect 197358 252855 197414 252864
rect 197372 252618 197400 252855
rect 197360 252612 197412 252618
rect 197360 252554 197412 252560
rect 197358 248840 197414 248849
rect 197358 248775 197360 248784
rect 197412 248775 197414 248784
rect 197360 248746 197412 248752
rect 197360 246356 197412 246362
rect 197360 246298 197412 246304
rect 197372 246265 197400 246298
rect 197358 246256 197414 246265
rect 197358 246191 197414 246200
rect 197268 242548 197320 242554
rect 197268 242490 197320 242496
rect 196808 239430 196860 239436
rect 197174 239456 197230 239465
rect 196716 234048 196768 234054
rect 196716 233990 196768 233996
rect 196624 229900 196676 229906
rect 196624 229842 196676 229848
rect 196820 225758 196848 239430
rect 197174 239391 197230 239400
rect 196808 225752 196860 225758
rect 196808 225694 196860 225700
rect 195796 222896 195848 222902
rect 195796 222838 195848 222844
rect 197280 208010 197308 242490
rect 197268 208004 197320 208010
rect 197268 207946 197320 207952
rect 195336 198008 195388 198014
rect 195336 197950 195388 197956
rect 195244 182980 195296 182986
rect 195244 182922 195296 182928
rect 195244 180124 195296 180130
rect 195244 180066 195296 180072
rect 195256 79422 195284 180066
rect 195348 84930 195376 197950
rect 196624 188488 196676 188494
rect 196624 188430 196676 188436
rect 195428 175976 195480 175982
rect 195428 175918 195480 175924
rect 195440 168298 195468 175918
rect 195428 168292 195480 168298
rect 195428 168234 195480 168240
rect 195520 114572 195572 114578
rect 195520 114514 195572 114520
rect 195336 84924 195388 84930
rect 195336 84866 195388 84872
rect 195428 84856 195480 84862
rect 195428 84798 195480 84804
rect 195244 79416 195296 79422
rect 195244 79358 195296 79364
rect 193864 65680 193916 65686
rect 193864 65622 193916 65628
rect 191104 4140 191156 4146
rect 191104 4082 191156 4088
rect 195440 3602 195468 84798
rect 195532 82754 195560 114514
rect 195520 82748 195572 82754
rect 195520 82690 195572 82696
rect 196636 51066 196664 188430
rect 196716 183592 196768 183598
rect 196716 183534 196768 183540
rect 196728 161362 196756 183534
rect 196808 182300 196860 182306
rect 196808 182242 196860 182248
rect 196820 162790 196848 182242
rect 198004 178696 198056 178702
rect 198004 178638 198056 178644
rect 196808 162784 196860 162790
rect 196808 162726 196860 162732
rect 196716 161356 196768 161362
rect 196716 161298 196768 161304
rect 196716 135312 196768 135318
rect 196716 135254 196768 135260
rect 196728 90982 196756 135254
rect 196808 122936 196860 122942
rect 196808 122878 196860 122884
rect 196716 90976 196768 90982
rect 196716 90918 196768 90924
rect 196820 85406 196848 122878
rect 196900 113212 196952 113218
rect 196900 113154 196952 113160
rect 196808 85400 196860 85406
rect 196808 85342 196860 85348
rect 196912 84114 196940 113154
rect 196900 84108 196952 84114
rect 196900 84050 196952 84056
rect 196624 51060 196676 51066
rect 196624 51002 196676 51008
rect 198016 26994 198044 178638
rect 198108 177449 198136 309130
rect 198646 271280 198702 271289
rect 198646 271215 198702 271224
rect 198464 242548 198516 242554
rect 198464 242490 198516 242496
rect 198476 242185 198504 242490
rect 198462 242176 198518 242185
rect 198462 242111 198518 242120
rect 198188 216708 198240 216714
rect 198188 216650 198240 216656
rect 198094 177440 198150 177449
rect 198094 177375 198150 177384
rect 198096 143608 198148 143614
rect 198096 143550 198148 143556
rect 198108 93226 198136 143550
rect 198200 95198 198228 216650
rect 198660 216034 198688 271215
rect 198844 232558 198872 332590
rect 199396 329118 199424 362306
rect 202604 361684 202656 361690
rect 202604 361626 202656 361632
rect 199476 360460 199528 360466
rect 199476 360402 199528 360408
rect 199488 338094 199516 360402
rect 202616 359924 202644 361626
rect 204536 360256 204588 360262
rect 204536 360198 204588 360204
rect 204548 359924 204576 360198
rect 206480 359924 206508 363190
rect 209056 359924 209084 365978
rect 209792 364334 209820 374002
rect 212908 369980 212960 369986
rect 212908 369922 212960 369928
rect 209792 364306 210648 364334
rect 210620 359938 210648 364306
rect 212920 362954 212948 369922
rect 213196 362982 213224 378150
rect 217968 375420 218020 375426
rect 217968 375362 218020 375368
rect 216588 364744 216640 364750
rect 216588 364686 216640 364692
rect 216600 362982 216628 364686
rect 213184 362976 213236 362982
rect 212920 362926 213040 362954
rect 210620 359910 211002 359938
rect 213012 359530 213040 362926
rect 213184 362918 213236 362924
rect 216588 362976 216640 362982
rect 216588 362918 216640 362924
rect 213196 362166 213224 362918
rect 217416 362908 217468 362914
rect 217416 362850 217468 362856
rect 213184 362160 213236 362166
rect 213184 362102 213236 362108
rect 214840 362160 214892 362166
rect 214840 362102 214892 362108
rect 214852 359924 214880 362102
rect 217428 359924 217456 362850
rect 217980 362409 218008 375362
rect 220096 373046 220124 391954
rect 220084 373040 220136 373046
rect 220084 372982 220136 372988
rect 220728 373040 220780 373046
rect 220728 372982 220780 372988
rect 220740 372706 220768 372982
rect 220728 372700 220780 372706
rect 220728 372642 220780 372648
rect 217966 362400 218022 362409
rect 217966 362335 218022 362344
rect 217980 362098 218008 362335
rect 217968 362092 218020 362098
rect 217968 362034 218020 362040
rect 219348 362092 219400 362098
rect 219348 362034 219400 362040
rect 219360 359924 219388 362034
rect 220740 361706 220768 372642
rect 223488 369912 223540 369918
rect 223488 369854 223540 369860
rect 223500 362273 223528 369854
rect 227720 364608 227772 364614
rect 227720 364550 227772 364556
rect 225788 363180 225840 363186
rect 225788 363122 225840 363128
rect 223486 362264 223542 362273
rect 223486 362199 223542 362208
rect 223500 362080 223528 362199
rect 223500 362052 223620 362080
rect 220740 361678 220952 361706
rect 220924 359938 220952 361678
rect 223592 359938 223620 362052
rect 225800 361758 225828 363122
rect 227732 363089 227760 364550
rect 227718 363080 227774 363089
rect 227718 363015 227774 363024
rect 225788 361752 225840 361758
rect 225788 361694 225840 361700
rect 220924 359910 221306 359938
rect 223592 359910 223882 359938
rect 225800 359924 225828 361694
rect 227732 359924 227760 363015
rect 228376 362914 228404 398890
rect 268384 397520 268436 397526
rect 268384 397462 268436 397468
rect 231858 394768 231914 394777
rect 231858 394703 231914 394712
rect 228364 362908 228416 362914
rect 228364 362850 228416 362856
rect 229652 362908 229704 362914
rect 229652 362850 229704 362856
rect 229664 359924 229692 362850
rect 231872 359938 231900 394703
rect 253202 389328 253258 389337
rect 253202 389263 253258 389272
rect 244924 387864 244976 387870
rect 244924 387806 244976 387812
rect 233884 375488 233936 375494
rect 233884 375430 233936 375436
rect 233896 363050 233924 375430
rect 244936 366042 244964 387806
rect 253216 374202 253244 389263
rect 263600 385144 263652 385150
rect 263600 385086 263652 385092
rect 263612 376786 263640 385086
rect 263600 376780 263652 376786
rect 263600 376722 263652 376728
rect 253204 374196 253256 374202
rect 253204 374138 253256 374144
rect 253216 373994 253244 374138
rect 253124 373966 253244 373994
rect 249708 370184 249760 370190
rect 249708 370126 249760 370132
rect 247040 366104 247092 366110
rect 247040 366046 247092 366052
rect 244924 366036 244976 366042
rect 244924 365978 244976 365984
rect 238668 365900 238720 365906
rect 238668 365842 238720 365848
rect 236092 364540 236144 364546
rect 236092 364482 236144 364488
rect 233884 363044 233936 363050
rect 233884 362986 233936 362992
rect 233896 359938 233924 362986
rect 231872 359910 232254 359938
rect 233896 359910 234186 359938
rect 236104 359924 236132 364482
rect 238680 359924 238708 365842
rect 242256 364676 242308 364682
rect 242256 364618 242308 364624
rect 242268 363186 242296 364618
rect 242256 363180 242308 363186
rect 242256 363122 242308 363128
rect 240600 361616 240652 361622
rect 240600 361558 240652 361564
rect 240612 359924 240640 361558
rect 242268 359938 242296 363122
rect 244936 359938 244964 365978
rect 247052 364449 247080 366046
rect 247038 364440 247094 364449
rect 247038 364375 247094 364384
rect 242268 359910 242558 359938
rect 244936 359910 245134 359938
rect 247052 359924 247080 364375
rect 249720 362370 249748 370126
rect 249708 362364 249760 362370
rect 249708 362306 249760 362312
rect 250904 362364 250956 362370
rect 250904 362306 250956 362312
rect 248970 361720 249026 361729
rect 248970 361655 249026 361664
rect 249706 361720 249762 361729
rect 249706 361655 249708 361664
rect 248984 359924 249012 361655
rect 249760 361655 249762 361664
rect 249708 361626 249760 361632
rect 250916 359924 250944 362306
rect 253124 359938 253152 373966
rect 255320 369164 255372 369170
rect 255320 369106 255372 369112
rect 255332 368558 255360 369106
rect 258724 368824 258776 368830
rect 258724 368766 258776 368772
rect 255320 368552 255372 368558
rect 255320 368494 255372 368500
rect 255332 364334 255360 368494
rect 257344 364540 257396 364546
rect 257344 364482 257396 364488
rect 255332 364306 255452 364334
rect 253124 359910 253506 359938
rect 255424 359924 255452 364306
rect 257356 360398 257384 364482
rect 258736 364478 258764 368766
rect 261850 364576 261906 364585
rect 261850 364511 261906 364520
rect 258724 364472 258776 364478
rect 258724 364414 258776 364420
rect 258736 361962 258764 364414
rect 258724 361956 258776 361962
rect 258724 361898 258776 361904
rect 259920 361956 259972 361962
rect 259920 361898 259972 361904
rect 257344 360392 257396 360398
rect 257344 360334 257396 360340
rect 257356 359924 257384 360334
rect 259932 359924 259960 361898
rect 261864 359924 261892 364511
rect 263612 359938 263640 376722
rect 265624 374672 265676 374678
rect 265624 374614 265676 374620
rect 265636 364478 265664 374614
rect 265624 364472 265676 364478
rect 265624 364414 265676 364420
rect 265636 364334 265664 364414
rect 265636 364306 265756 364334
rect 263612 359910 263810 359938
rect 265728 359924 265756 364306
rect 268396 363050 268424 397462
rect 286336 396098 286364 484366
rect 323584 418192 323636 418198
rect 323584 418134 323636 418140
rect 320272 400240 320324 400246
rect 320272 400182 320324 400188
rect 289084 396160 289136 396166
rect 289084 396102 289136 396108
rect 286324 396092 286376 396098
rect 286324 396034 286376 396040
rect 278044 393372 278096 393378
rect 278044 393314 278096 393320
rect 278056 383654 278084 393314
rect 278056 383626 278176 383654
rect 270224 368688 270276 368694
rect 270224 368630 270276 368636
rect 270236 367470 270264 368630
rect 269856 367464 269908 367470
rect 269856 367406 269908 367412
rect 270224 367464 270276 367470
rect 270224 367406 270276 367412
rect 268384 363044 268436 363050
rect 268384 362986 268436 362992
rect 268396 359938 268424 362986
rect 268318 359910 268424 359938
rect 269868 359938 269896 367406
rect 275928 366104 275980 366110
rect 275928 366046 275980 366052
rect 275940 362302 275968 366046
rect 275928 362296 275980 362302
rect 275928 362238 275980 362244
rect 276664 362296 276716 362302
rect 276664 362238 276716 362244
rect 274730 361992 274786 362001
rect 274730 361927 274786 361936
rect 274744 361593 274772 361927
rect 274730 361584 274786 361593
rect 274730 361519 274786 361528
rect 272156 360392 272208 360398
rect 272156 360334 272208 360340
rect 272168 359938 272196 360334
rect 269868 359910 270250 359938
rect 271984 359924 272196 359938
rect 274744 359924 274772 361519
rect 276676 359924 276704 362238
rect 278148 360534 278176 383626
rect 284300 372768 284352 372774
rect 284300 372710 284352 372716
rect 284312 370530 284340 372710
rect 284300 370524 284352 370530
rect 284300 370466 284352 370472
rect 282920 370116 282972 370122
rect 282920 370058 282972 370064
rect 282932 368694 282960 370058
rect 282920 368688 282972 368694
rect 282920 368630 282972 368636
rect 281172 361888 281224 361894
rect 281172 361830 281224 361836
rect 281184 361622 281212 361830
rect 281172 361616 281224 361622
rect 281172 361558 281224 361564
rect 278136 360528 278188 360534
rect 278136 360470 278188 360476
rect 278596 360528 278648 360534
rect 278596 360470 278648 360476
rect 278608 359924 278636 360470
rect 281184 359924 281212 361558
rect 282932 359938 282960 368630
rect 286336 367402 286364 396034
rect 286324 367396 286376 367402
rect 286324 367338 286376 367344
rect 286600 367396 286652 367402
rect 286600 367338 286652 367344
rect 285034 363216 285090 363225
rect 285034 363151 285090 363160
rect 271984 359910 272182 359924
rect 282932 359910 283130 359938
rect 285048 359924 285076 363151
rect 286612 359938 286640 367338
rect 289096 364334 289124 396102
rect 291844 394800 291896 394806
rect 291844 394742 291896 394748
rect 289096 364306 289216 364334
rect 289188 361962 289216 364306
rect 289176 361956 289228 361962
rect 289176 361898 289228 361904
rect 289188 359938 289216 361898
rect 291474 360224 291530 360233
rect 291474 360159 291530 360168
rect 291488 359938 291516 360159
rect 291856 359938 291884 394742
rect 304264 394732 304316 394738
rect 304264 394674 304316 394680
rect 301504 385076 301556 385082
rect 301504 385018 301556 385024
rect 297364 376100 297416 376106
rect 297364 376042 297416 376048
rect 295340 370048 295392 370054
rect 295340 369990 295392 369996
rect 295352 367198 295380 369990
rect 293224 367192 293276 367198
rect 293224 367134 293276 367140
rect 295340 367192 295392 367198
rect 295340 367134 295392 367140
rect 295616 367192 295668 367198
rect 295616 367134 295668 367140
rect 293236 360505 293264 367134
rect 293222 360496 293278 360505
rect 293222 360431 293278 360440
rect 286612 359910 286994 359938
rect 289188 359910 289570 359938
rect 291488 359924 291884 359938
rect 291502 359910 291884 359924
rect 293236 359938 293264 360431
rect 295628 359938 295656 367134
rect 297376 365906 297404 376042
rect 300124 367328 300176 367334
rect 300124 367270 300176 367276
rect 297364 365900 297416 365906
rect 297364 365842 297416 365848
rect 297376 364334 297404 365842
rect 297376 364306 297496 364334
rect 297468 359938 297496 364306
rect 300136 361865 300164 367270
rect 300122 361856 300178 361865
rect 300122 361791 300178 361800
rect 300136 359938 300164 361791
rect 301516 361622 301544 385018
rect 304276 364334 304304 394674
rect 316684 393440 316736 393446
rect 316684 393382 316736 393388
rect 309140 388476 309192 388482
rect 309140 388418 309192 388424
rect 305644 376916 305696 376922
rect 305644 376858 305696 376864
rect 304276 364306 304396 364334
rect 301504 361616 301556 361622
rect 301504 361558 301556 361564
rect 293236 359910 293434 359938
rect 295628 359910 296010 359938
rect 297468 359910 297942 359938
rect 299874 359910 300164 359938
rect 301516 359938 301544 361558
rect 304368 360233 304396 364306
rect 305656 363254 305684 376858
rect 305644 363248 305696 363254
rect 305644 363190 305696 363196
rect 306288 363248 306340 363254
rect 306288 363190 306340 363196
rect 304354 360224 304410 360233
rect 304354 360159 304410 360168
rect 301516 359910 301806 359938
rect 304368 359924 304396 360159
rect 306300 359924 306328 363190
rect 309152 360874 309180 388418
rect 313280 376848 313332 376854
rect 313280 376790 313332 376796
rect 313292 376106 313320 376790
rect 313280 376100 313332 376106
rect 313280 376042 313332 376048
rect 312728 365764 312780 365770
rect 312728 365706 312780 365712
rect 309968 364676 310020 364682
rect 309968 364618 310020 364624
rect 309980 362234 310008 364618
rect 309968 362228 310020 362234
rect 309968 362170 310020 362176
rect 310796 361820 310848 361826
rect 310796 361762 310848 361768
rect 308496 360868 308548 360874
rect 308496 360810 308548 360816
rect 309140 360868 309192 360874
rect 309140 360810 309192 360816
rect 308508 359938 308536 360810
rect 310808 360466 310836 361762
rect 310796 360460 310848 360466
rect 310796 360402 310848 360408
rect 308246 359910 308536 359938
rect 310808 359924 310836 360402
rect 312740 360262 312768 365706
rect 316696 362506 316724 393382
rect 318800 376100 318852 376106
rect 318800 376042 318852 376048
rect 316684 362500 316736 362506
rect 316684 362442 316736 362448
rect 317328 362500 317380 362506
rect 317328 362442 317380 362448
rect 317052 361752 317104 361758
rect 317052 361694 317104 361700
rect 314660 360596 314712 360602
rect 314660 360538 314712 360544
rect 312728 360256 312780 360262
rect 312728 360198 312780 360204
rect 312740 359924 312768 360198
rect 314672 359938 314700 360538
rect 314672 359924 314884 359938
rect 314686 359910 314884 359924
rect 271984 359553 272012 359910
rect 212552 359502 213040 359530
rect 271970 359544 272026 359553
rect 212552 359446 212580 359502
rect 271970 359479 272026 359488
rect 314856 359446 314884 359910
rect 317064 359553 317092 361694
rect 317340 359666 317368 362442
rect 318812 359938 318840 376042
rect 320180 366104 320232 366110
rect 320180 366046 320232 366052
rect 319444 361956 319496 361962
rect 319444 361898 319496 361904
rect 318812 359910 319300 359938
rect 317262 359650 317552 359666
rect 317262 359644 317564 359650
rect 317262 359638 317512 359644
rect 317512 359586 317564 359592
rect 317050 359544 317106 359553
rect 317050 359479 317106 359488
rect 212540 359440 212592 359446
rect 212540 359382 212592 359388
rect 314844 359440 314896 359446
rect 314844 359382 314896 359388
rect 319272 359258 319300 359910
rect 199672 359230 200054 359258
rect 319194 359230 319392 359258
rect 199672 358873 199700 359230
rect 199844 358964 199896 358970
rect 199844 358906 199896 358912
rect 199658 358864 199714 358873
rect 199658 358799 199714 358808
rect 199856 357406 199884 358906
rect 319364 358873 319392 359230
rect 319350 358864 319406 358873
rect 319350 358799 319406 358808
rect 199844 357400 199896 357406
rect 199844 357342 199896 357348
rect 319350 356416 319406 356425
rect 319350 356351 319406 356360
rect 199476 338088 199528 338094
rect 199476 338030 199528 338036
rect 319364 335354 319392 356351
rect 319456 351218 319484 361898
rect 319902 361856 319958 361865
rect 319902 361791 319958 361800
rect 319536 359644 319588 359650
rect 319536 359586 319588 359592
rect 319548 358086 319576 359586
rect 319536 358080 319588 358086
rect 319536 358022 319588 358028
rect 319916 355366 319944 361791
rect 319904 355360 319956 355366
rect 319904 355302 319956 355308
rect 319444 351212 319496 351218
rect 319444 351154 319496 351160
rect 319272 335326 319392 335354
rect 199384 329112 199436 329118
rect 199384 329054 199436 329060
rect 198922 313440 198978 313449
rect 198922 313375 198978 313384
rect 198832 232552 198884 232558
rect 198832 232494 198884 232500
rect 198648 216028 198700 216034
rect 198648 215970 198700 215976
rect 198280 134020 198332 134026
rect 198280 133962 198332 133968
rect 198188 95192 198240 95198
rect 198188 95134 198240 95140
rect 198096 93220 198148 93226
rect 198096 93162 198148 93168
rect 198292 91633 198320 133962
rect 198936 93770 198964 313375
rect 199672 240230 200054 240258
rect 199672 240174 199700 240230
rect 199660 240168 199712 240174
rect 199660 240110 199712 240116
rect 199856 238754 199884 240230
rect 318523 240094 318564 240122
rect 201408 239964 201460 239970
rect 201408 239906 201460 239912
rect 201420 239873 201448 239906
rect 201406 239864 201462 239873
rect 201926 239850 201954 240040
rect 203858 239850 203886 240040
rect 201406 239799 201462 239808
rect 201512 239822 201954 239850
rect 202892 239822 203886 239850
rect 200856 239692 200908 239698
rect 200856 239634 200908 239640
rect 199856 238726 199976 238754
rect 199948 237454 199976 238726
rect 199936 237448 199988 237454
rect 199936 237390 199988 237396
rect 200764 190120 200816 190126
rect 200764 190062 200816 190068
rect 199384 151836 199436 151842
rect 199384 151778 199436 151784
rect 198924 93764 198976 93770
rect 198924 93706 198976 93712
rect 198278 91624 198334 91633
rect 198278 91559 198334 91568
rect 199396 90778 199424 151778
rect 199476 103556 199528 103562
rect 199476 103498 199528 103504
rect 199384 90772 199436 90778
rect 199384 90714 199436 90720
rect 199488 80034 199516 103498
rect 199476 80028 199528 80034
rect 199476 79970 199528 79976
rect 200776 79354 200804 190062
rect 200868 182918 200896 239634
rect 201408 238128 201460 238134
rect 201408 238070 201460 238076
rect 201420 237182 201448 238070
rect 201408 237176 201460 237182
rect 201408 237118 201460 237124
rect 201512 223514 201540 239822
rect 201592 239556 201644 239562
rect 201592 239498 201644 239504
rect 201604 226166 201632 239498
rect 202328 237448 202380 237454
rect 202328 237390 202380 237396
rect 202236 227112 202288 227118
rect 202236 227054 202288 227060
rect 201592 226160 201644 226166
rect 201592 226102 201644 226108
rect 201500 223508 201552 223514
rect 201500 223450 201552 223456
rect 202144 184204 202196 184210
rect 202144 184146 202196 184152
rect 200856 182912 200908 182918
rect 200856 182854 200908 182860
rect 201592 176792 201644 176798
rect 201592 176734 201644 176740
rect 201604 176662 201632 176734
rect 201592 176656 201644 176662
rect 201592 176598 201644 176604
rect 200856 146396 200908 146402
rect 200856 146338 200908 146344
rect 200868 93294 200896 146338
rect 200948 113280 201000 113286
rect 200948 113222 201000 113228
rect 200856 93288 200908 93294
rect 200856 93230 200908 93236
rect 200960 88262 200988 113222
rect 200948 88256 201000 88262
rect 200948 88198 201000 88204
rect 200764 79348 200816 79354
rect 200764 79290 200816 79296
rect 198004 26988 198056 26994
rect 198004 26930 198056 26936
rect 202156 11830 202184 184146
rect 202248 95130 202276 227054
rect 202340 178702 202368 237390
rect 202892 230382 202920 239822
rect 204902 239456 204958 239465
rect 204902 239391 204958 239400
rect 204168 238196 204220 238202
rect 204168 238138 204220 238144
rect 204180 231674 204208 238138
rect 204168 231668 204220 231674
rect 204168 231610 204220 231616
rect 202880 230376 202932 230382
rect 202880 230318 202932 230324
rect 203524 230376 203576 230382
rect 203524 230318 203576 230324
rect 202788 226160 202840 226166
rect 202788 226102 202840 226108
rect 202800 225690 202828 226102
rect 202788 225684 202840 225690
rect 202788 225626 202840 225632
rect 202420 223508 202472 223514
rect 202420 223450 202472 223456
rect 202328 178696 202380 178702
rect 202328 178638 202380 178644
rect 202432 177410 202460 223450
rect 202420 177404 202472 177410
rect 202420 177346 202472 177352
rect 203536 177342 203564 230318
rect 203524 177336 203576 177342
rect 203524 177278 203576 177284
rect 202420 136740 202472 136746
rect 202420 136682 202472 136688
rect 202328 131164 202380 131170
rect 202328 131106 202380 131112
rect 202236 95124 202288 95130
rect 202236 95066 202288 95072
rect 202340 86834 202368 131106
rect 202432 92342 202460 136682
rect 203524 121576 203576 121582
rect 203524 121518 203576 121524
rect 202420 92336 202472 92342
rect 202420 92278 202472 92284
rect 202328 86828 202380 86834
rect 202328 86770 202380 86776
rect 203536 81326 203564 121518
rect 203616 117428 203668 117434
rect 203616 117370 203668 117376
rect 203628 92478 203656 117370
rect 204916 95062 204944 239391
rect 204996 238060 205048 238066
rect 204996 238002 205048 238008
rect 205008 227526 205036 238002
rect 205836 233306 205864 240040
rect 207662 237960 207718 237969
rect 207662 237895 207718 237904
rect 205640 233300 205692 233306
rect 205640 233242 205692 233248
rect 205824 233300 205876 233306
rect 205824 233242 205876 233248
rect 205652 231742 205680 233242
rect 206468 232620 206520 232626
rect 206468 232562 206520 232568
rect 205640 231736 205692 231742
rect 205640 231678 205692 231684
rect 204996 227520 205048 227526
rect 204996 227462 205048 227468
rect 204996 182368 205048 182374
rect 204996 182310 205048 182316
rect 205008 166870 205036 182310
rect 206480 181529 206508 232562
rect 206282 181520 206338 181529
rect 206282 181455 206338 181464
rect 206466 181520 206522 181529
rect 206466 181455 206522 181464
rect 205640 176724 205692 176730
rect 205640 176666 205692 176672
rect 205652 175166 205680 176666
rect 205640 175160 205692 175166
rect 205640 175102 205692 175108
rect 204996 166864 205048 166870
rect 204996 166806 205048 166812
rect 205088 150476 205140 150482
rect 205088 150418 205140 150424
rect 204996 140888 205048 140894
rect 204996 140830 205048 140836
rect 204904 95056 204956 95062
rect 204904 94998 204956 95004
rect 203616 92472 203668 92478
rect 203616 92414 203668 92420
rect 205008 88194 205036 140830
rect 205100 111790 205128 150418
rect 205180 111920 205232 111926
rect 205180 111862 205232 111868
rect 205088 111784 205140 111790
rect 205088 111726 205140 111732
rect 205088 100768 205140 100774
rect 205088 100710 205140 100716
rect 204996 88188 205048 88194
rect 204996 88130 205048 88136
rect 203524 81320 203576 81326
rect 203524 81262 203576 81268
rect 205100 77246 205128 100710
rect 205192 88330 205220 111862
rect 205180 88324 205232 88330
rect 205180 88266 205232 88272
rect 205088 77240 205140 77246
rect 205088 77182 205140 77188
rect 206296 35358 206324 181455
rect 206376 151904 206428 151910
rect 206376 151846 206428 151852
rect 206388 89350 206416 151846
rect 206468 143676 206520 143682
rect 206468 143618 206520 143624
rect 206376 89344 206428 89350
rect 206376 89286 206428 89292
rect 206480 85474 206508 143618
rect 207676 93809 207704 237895
rect 208412 215218 208440 240040
rect 210364 239850 210392 240040
rect 210364 239822 210464 239850
rect 210436 237046 210464 239822
rect 210424 237040 210476 237046
rect 210424 236982 210476 236988
rect 210436 225622 210464 236982
rect 211618 235240 211674 235249
rect 211618 235175 211674 235184
rect 211632 230382 211660 235175
rect 212276 234462 212304 240040
rect 214806 239850 214834 240040
rect 216738 239850 216766 240040
rect 213932 239822 214834 239850
rect 216692 239822 216766 239850
rect 218736 239850 218764 240040
rect 218736 239822 218836 239850
rect 211804 234456 211856 234462
rect 211804 234398 211856 234404
rect 212264 234456 212316 234462
rect 212264 234398 212316 234404
rect 211620 230376 211672 230382
rect 211620 230318 211672 230324
rect 210424 225616 210476 225622
rect 210424 225558 210476 225564
rect 208400 215212 208452 215218
rect 208400 215154 208452 215160
rect 208412 214878 208440 215154
rect 208400 214872 208452 214878
rect 208400 214814 208452 214820
rect 209044 214872 209096 214878
rect 209044 214814 209096 214820
rect 209056 184249 209084 214814
rect 211816 199442 211844 234398
rect 213368 229968 213420 229974
rect 213368 229910 213420 229916
rect 213276 225820 213328 225826
rect 213276 225762 213328 225768
rect 211804 199436 211856 199442
rect 211804 199378 211856 199384
rect 213184 198280 213236 198286
rect 213184 198222 213236 198228
rect 209134 191176 209190 191185
rect 209134 191111 209190 191120
rect 209042 184240 209098 184249
rect 209042 184175 209098 184184
rect 209044 181620 209096 181626
rect 209044 181562 209096 181568
rect 208400 153876 208452 153882
rect 208400 153818 208452 153824
rect 208412 150346 208440 153818
rect 208492 150544 208544 150550
rect 208492 150486 208544 150492
rect 208400 150340 208452 150346
rect 208400 150282 208452 150288
rect 208504 144226 208532 150486
rect 208492 144220 208544 144226
rect 208492 144162 208544 144168
rect 207848 116068 207900 116074
rect 207848 116010 207900 116016
rect 207756 100836 207808 100842
rect 207756 100778 207808 100784
rect 207662 93800 207718 93809
rect 207662 93735 207718 93744
rect 206468 85468 206520 85474
rect 206468 85410 206520 85416
rect 207768 74526 207796 100778
rect 207860 94586 207888 116010
rect 207848 94580 207900 94586
rect 207848 94522 207900 94528
rect 207756 74520 207808 74526
rect 207756 74462 207808 74468
rect 206284 35352 206336 35358
rect 206284 35294 206336 35300
rect 209056 22846 209084 181562
rect 209148 86290 209176 191111
rect 210424 185836 210476 185842
rect 210424 185778 210476 185784
rect 209228 142248 209280 142254
rect 209228 142190 209280 142196
rect 209136 86284 209188 86290
rect 209136 86226 209188 86232
rect 209240 79898 209268 142190
rect 209228 79892 209280 79898
rect 209228 79834 209280 79840
rect 210436 39574 210464 185778
rect 211804 176248 211856 176254
rect 211804 176190 211856 176196
rect 210516 132932 210568 132938
rect 210516 132874 210568 132880
rect 210528 82822 210556 132874
rect 210516 82816 210568 82822
rect 210516 82758 210568 82764
rect 210424 39568 210476 39574
rect 210424 39510 210476 39516
rect 211816 36650 211844 176190
rect 211896 139528 211948 139534
rect 211896 139470 211948 139476
rect 211908 92410 211936 139470
rect 211988 102196 212040 102202
rect 211988 102138 212040 102144
rect 211896 92404 211948 92410
rect 211896 92346 211948 92352
rect 212000 91050 212028 102138
rect 211988 91044 212040 91050
rect 211988 90986 212040 90992
rect 211804 36644 211856 36650
rect 211804 36586 211856 36592
rect 209044 22840 209096 22846
rect 209044 22782 209096 22788
rect 202144 11824 202196 11830
rect 202144 11766 202196 11772
rect 213196 4894 213224 198222
rect 213288 198014 213316 225762
rect 213276 198008 213328 198014
rect 213276 197950 213328 197956
rect 213276 195560 213328 195566
rect 213276 195502 213328 195508
rect 213288 28354 213316 195502
rect 213380 185842 213408 229910
rect 213932 224738 213960 239822
rect 216692 228954 216720 239822
rect 218704 237448 218756 237454
rect 218704 237390 218756 237396
rect 216680 228948 216732 228954
rect 216680 228890 216732 228896
rect 216692 227798 216720 228890
rect 216680 227792 216732 227798
rect 216680 227734 216732 227740
rect 217324 227792 217376 227798
rect 217324 227734 217376 227740
rect 215942 227080 215998 227089
rect 215942 227015 215998 227024
rect 213920 224732 213972 224738
rect 213920 224674 213972 224680
rect 213932 224466 213960 224674
rect 213920 224460 213972 224466
rect 213920 224402 213972 224408
rect 214656 224460 214708 224466
rect 214656 224402 214708 224408
rect 214668 207874 214696 224402
rect 214656 207868 214708 207874
rect 214656 207810 214708 207816
rect 214564 207664 214616 207670
rect 214564 207606 214616 207612
rect 213368 185836 213420 185842
rect 213368 185778 213420 185784
rect 214576 178673 214604 207606
rect 214656 182232 214708 182238
rect 214656 182174 214708 182180
rect 214562 178664 214618 178673
rect 214562 178599 214618 178608
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 176225 213960 176598
rect 213918 176216 213974 176225
rect 213918 176151 213974 176160
rect 214104 176180 214156 176186
rect 214104 176122 214156 176128
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175137 213960 175170
rect 214012 175160 214064 175166
rect 213918 175128 213974 175137
rect 214012 175102 214064 175108
rect 213918 175063 213974 175072
rect 214024 174729 214052 175102
rect 214010 174720 214066 174729
rect 214010 174655 214066 174664
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173777 213960 173810
rect 214012 173800 214064 173806
rect 213918 173768 213974 173777
rect 214012 173742 214064 173748
rect 213918 173703 213974 173712
rect 214024 173369 214052 173742
rect 214010 173360 214066 173369
rect 214010 173295 214066 173304
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172417 213960 172450
rect 213918 172408 213974 172417
rect 213918 172343 213974 172352
rect 214116 172009 214144 176122
rect 214102 172000 214158 172009
rect 214102 171935 214158 171944
rect 214012 171080 214064 171086
rect 213918 171048 213974 171057
rect 214012 171022 214064 171028
rect 213918 170983 213920 170992
rect 213972 170983 213974 170992
rect 213920 170954 213972 170960
rect 214024 170785 214052 171022
rect 214010 170776 214066 170785
rect 214010 170711 214066 170720
rect 214668 169425 214696 182174
rect 214748 176928 214800 176934
rect 214748 176870 214800 176876
rect 214654 169416 214710 169425
rect 214654 169351 214710 169360
rect 214012 168360 214064 168366
rect 213918 168328 213974 168337
rect 214012 168302 214064 168308
rect 213918 168263 213920 168272
rect 213972 168263 213974 168272
rect 213920 168234 213972 168240
rect 214024 168065 214052 168302
rect 214010 168056 214066 168065
rect 214010 167991 214066 168000
rect 214104 167000 214156 167006
rect 213918 166968 213974 166977
rect 214104 166942 214156 166948
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 213932 166870 213960 166903
rect 214012 166874 214064 166880
rect 213920 166864 213972 166870
rect 213920 166806 213972 166812
rect 214024 166161 214052 166874
rect 214116 166705 214144 166942
rect 214102 166696 214158 166705
rect 214102 166631 214158 166640
rect 214010 166152 214066 166161
rect 214010 166087 214066 166096
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 165345 213960 165514
rect 214012 165504 214064 165510
rect 214012 165446 214064 165452
rect 213918 165336 213974 165345
rect 213918 165271 213974 165280
rect 214024 164801 214052 165446
rect 214010 164792 214066 164801
rect 214010 164727 214066 164736
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163441 213960 164154
rect 213918 163432 213974 163441
rect 213918 163367 213974 163376
rect 214012 162852 214064 162858
rect 214012 162794 214064 162800
rect 213920 162784 213972 162790
rect 213918 162752 213920 162761
rect 213972 162752 213974 162761
rect 213918 162687 213974 162696
rect 214024 162081 214052 162794
rect 214010 162072 214066 162081
rect 214010 162007 214066 162016
rect 213920 161424 213972 161430
rect 213918 161392 213920 161401
rect 213972 161392 213974 161401
rect 213918 161327 213974 161336
rect 214012 161356 214064 161362
rect 214012 161298 214064 161304
rect 214024 160857 214052 161298
rect 214010 160848 214066 160857
rect 214010 160783 214066 160792
rect 214012 160064 214064 160070
rect 214012 160006 214064 160012
rect 213920 159996 213972 160002
rect 213920 159938 213972 159944
rect 213932 159905 213960 159938
rect 213918 159896 213974 159905
rect 213918 159831 213974 159840
rect 214024 159497 214052 160006
rect 214010 159488 214066 159497
rect 214010 159423 214066 159432
rect 213920 158704 213972 158710
rect 213920 158646 213972 158652
rect 213932 157457 213960 158646
rect 213918 157448 213974 157457
rect 213918 157383 213974 157392
rect 213920 157344 213972 157350
rect 213918 157312 213920 157321
rect 213972 157312 213974 157321
rect 213918 157247 213974 157256
rect 214012 157276 214064 157282
rect 214012 157218 214064 157224
rect 214024 156913 214052 157218
rect 214010 156904 214066 156913
rect 214010 156839 214066 156848
rect 213918 155952 213974 155961
rect 213918 155887 213920 155896
rect 213972 155887 213974 155896
rect 213920 155858 213972 155864
rect 214012 155848 214064 155854
rect 214012 155790 214064 155796
rect 214024 155417 214052 155790
rect 214010 155408 214066 155417
rect 214010 155343 214066 155352
rect 213918 153912 213974 153921
rect 213918 153847 213974 153856
rect 213932 153270 213960 153847
rect 213920 153264 213972 153270
rect 213366 153232 213422 153241
rect 213920 153206 213972 153212
rect 213366 153167 213422 153176
rect 213380 88058 213408 153167
rect 214010 152688 214066 152697
rect 214010 152623 214066 152632
rect 213918 152008 213974 152017
rect 213918 151943 213974 151952
rect 213932 151910 213960 151943
rect 213920 151904 213972 151910
rect 213920 151846 213972 151852
rect 214024 151842 214052 152623
rect 214012 151836 214064 151842
rect 214012 151778 214064 151784
rect 214010 150920 214066 150929
rect 214010 150855 214066 150864
rect 213918 150648 213974 150657
rect 213918 150583 213974 150592
rect 213932 150482 213960 150583
rect 214024 150550 214052 150855
rect 214012 150544 214064 150550
rect 214012 150486 214064 150492
rect 213920 150476 213972 150482
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 213920 150340 213972 150346
rect 213920 150282 213972 150288
rect 213932 149569 213960 150282
rect 214024 150113 214052 150350
rect 214010 150104 214066 150113
rect 214010 150039 214066 150048
rect 213918 149560 213974 149569
rect 213918 149495 213974 149504
rect 214760 148889 214788 176870
rect 214932 174548 214984 174554
rect 214932 174490 214984 174496
rect 214944 169697 214972 174490
rect 214930 169688 214986 169697
rect 214930 169623 214986 169632
rect 215022 151872 215078 151881
rect 215022 151807 215078 151816
rect 214746 148880 214802 148889
rect 214746 148815 214802 148824
rect 214562 148064 214618 148073
rect 214562 147999 214618 148008
rect 214010 146704 214066 146713
rect 214010 146639 214066 146648
rect 213918 146432 213974 146441
rect 213918 146367 213920 146376
rect 213972 146367 213974 146376
rect 213920 146338 213972 146344
rect 214024 146334 214052 146639
rect 214012 146328 214064 146334
rect 214012 146270 214064 146276
rect 213918 145344 213974 145353
rect 213918 145279 213974 145288
rect 213932 144974 213960 145279
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 214010 143984 214066 143993
rect 214010 143919 214066 143928
rect 213920 143676 213972 143682
rect 213920 143618 213972 143624
rect 213932 143585 213960 143618
rect 214024 143614 214052 143919
rect 214012 143608 214064 143614
rect 213918 143576 213974 143585
rect 214012 143550 214064 143556
rect 213918 143511 213974 143520
rect 214010 142760 214066 142769
rect 214010 142695 214066 142704
rect 213918 142352 213974 142361
rect 213918 142287 213974 142296
rect 213932 142254 213960 142287
rect 213920 142248 213972 142254
rect 213920 142190 213972 142196
rect 214024 142186 214052 142695
rect 214012 142180 214064 142186
rect 214012 142122 214064 142128
rect 214010 141400 214066 141409
rect 214010 141335 214066 141344
rect 214024 140894 214052 141335
rect 214012 140888 214064 140894
rect 213918 140856 213974 140865
rect 214012 140830 214064 140836
rect 213918 140791 213920 140800
rect 213972 140791 213974 140800
rect 213920 140762 213972 140768
rect 213918 140040 213974 140049
rect 213918 139975 213974 139984
rect 213932 139466 213960 139975
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 213918 138816 213974 138825
rect 213918 138751 213974 138760
rect 213932 138038 213960 138751
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 214010 137456 214066 137465
rect 214010 137391 214066 137400
rect 213918 136776 213974 136785
rect 213918 136711 213920 136720
rect 213972 136711 213974 136720
rect 213920 136682 213972 136688
rect 214024 136678 214052 137391
rect 214012 136672 214064 136678
rect 214012 136614 214064 136620
rect 213918 136096 213974 136105
rect 213918 136031 213974 136040
rect 213932 135318 213960 136031
rect 213920 135312 213972 135318
rect 213920 135254 213972 135260
rect 214010 134328 214066 134337
rect 214010 134263 214066 134272
rect 213918 134056 213974 134065
rect 214024 134026 214052 134263
rect 213918 133991 213974 134000
rect 214012 134020 214064 134026
rect 213932 133958 213960 133991
rect 214012 133962 214064 133968
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 213918 132968 213974 132977
rect 213918 132903 213920 132912
rect 213972 132903 213974 132912
rect 213920 132874 213972 132880
rect 213918 132832 213974 132841
rect 213918 132767 213974 132776
rect 213932 132530 213960 132767
rect 213920 132524 213972 132530
rect 213920 132466 213972 132472
rect 213918 131472 213974 131481
rect 213918 131407 213974 131416
rect 213932 131170 213960 131407
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 214010 130112 214066 130121
rect 214010 130047 214066 130056
rect 213920 129872 213972 129878
rect 213918 129840 213920 129849
rect 213972 129840 213974 129849
rect 214024 129810 214052 130047
rect 213918 129775 213974 129784
rect 214012 129804 214064 129810
rect 214012 129746 214064 129752
rect 213918 128888 213974 128897
rect 213918 128823 213974 128832
rect 213932 128382 213960 128823
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 214010 127528 214066 127537
rect 214010 127463 214066 127472
rect 213918 127120 213974 127129
rect 214024 127090 214052 127463
rect 213918 127055 213974 127064
rect 214012 127084 214064 127090
rect 213932 127022 213960 127055
rect 214012 127026 214064 127032
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 214010 126168 214066 126177
rect 214010 126103 214066 126112
rect 213918 125760 213974 125769
rect 214024 125730 214052 126103
rect 213918 125695 213974 125704
rect 214012 125724 214064 125730
rect 213932 125662 213960 125695
rect 214012 125666 214064 125672
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214010 124808 214066 124817
rect 214010 124743 214066 124752
rect 213918 124400 213974 124409
rect 213918 124335 213974 124344
rect 213932 124302 213960 124335
rect 213920 124296 213972 124302
rect 213920 124238 213972 124244
rect 214024 124234 214052 124743
rect 214012 124228 214064 124234
rect 214012 124170 214064 124176
rect 214010 123584 214066 123593
rect 214010 123519 214066 123528
rect 213918 123176 213974 123185
rect 213918 123111 213974 123120
rect 213932 122942 213960 123111
rect 213920 122936 213972 122942
rect 213920 122878 213972 122884
rect 214024 122874 214052 123519
rect 214012 122868 214064 122874
rect 214012 122810 214064 122816
rect 214010 122224 214066 122233
rect 214010 122159 214066 122168
rect 214024 121582 214052 122159
rect 214012 121576 214064 121582
rect 213918 121544 213974 121553
rect 214012 121518 214064 121524
rect 213918 121479 213920 121488
rect 213972 121479 213974 121488
rect 213920 121450 213972 121456
rect 214010 120864 214066 120873
rect 214010 120799 214066 120808
rect 214024 120222 214052 120799
rect 214012 120216 214064 120222
rect 213918 120184 213974 120193
rect 214012 120158 214064 120164
rect 213918 120119 213920 120128
rect 213972 120119 213974 120128
rect 213920 120090 213972 120096
rect 214010 119640 214066 119649
rect 214010 119575 214066 119584
rect 213458 119096 213514 119105
rect 213458 119031 213514 119040
rect 213368 88052 213420 88058
rect 213368 87994 213420 88000
rect 213472 78674 213500 119031
rect 213918 118960 213974 118969
rect 213918 118895 213974 118904
rect 213932 118794 213960 118895
rect 214024 118862 214052 119575
rect 214012 118856 214064 118862
rect 214012 118798 214064 118804
rect 213920 118788 213972 118794
rect 213920 118730 213972 118736
rect 214010 117600 214066 117609
rect 214010 117535 214066 117544
rect 213920 117428 213972 117434
rect 213920 117370 213972 117376
rect 213932 117337 213960 117370
rect 214024 117366 214052 117535
rect 214012 117360 214064 117366
rect 213918 117328 213974 117337
rect 214012 117302 214064 117308
rect 213918 117263 213974 117272
rect 214010 116240 214066 116249
rect 214010 116175 214066 116184
rect 213920 116068 213972 116074
rect 213920 116010 213972 116016
rect 213932 115977 213960 116010
rect 214024 116006 214052 116175
rect 214012 116000 214064 116006
rect 213918 115968 213974 115977
rect 214012 115942 214064 115948
rect 213918 115903 213974 115912
rect 213918 115016 213974 115025
rect 213918 114951 213974 114960
rect 213932 114578 213960 114951
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 214010 113656 214066 113665
rect 214010 113591 214066 113600
rect 214024 113286 214052 113591
rect 214012 113280 214064 113286
rect 213918 113248 213974 113257
rect 214012 113222 214064 113228
rect 213918 113183 213920 113192
rect 213972 113183 213974 113192
rect 213920 113154 213972 113160
rect 214010 112296 214066 112305
rect 214010 112231 214066 112240
rect 213920 111920 213972 111926
rect 213918 111888 213920 111897
rect 213972 111888 213974 111897
rect 214024 111858 214052 112231
rect 213918 111823 213974 111832
rect 214012 111852 214064 111858
rect 214012 111794 214064 111800
rect 214010 110936 214066 110945
rect 214010 110871 214066 110880
rect 213920 110560 213972 110566
rect 213918 110528 213920 110537
rect 213972 110528 213974 110537
rect 214024 110498 214052 110871
rect 213918 110463 213974 110472
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 214010 109712 214066 109721
rect 214010 109647 214066 109656
rect 213918 109168 213974 109177
rect 213918 109103 213920 109112
rect 213972 109103 213974 109112
rect 213920 109074 213972 109080
rect 214024 109070 214052 109647
rect 214012 109064 214064 109070
rect 214012 109006 214064 109012
rect 214010 108352 214066 108361
rect 214010 108287 214066 108296
rect 213918 107944 213974 107953
rect 213918 107879 213974 107888
rect 213932 107710 213960 107879
rect 214024 107778 214052 108287
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 106992 214066 107001
rect 214010 106927 214066 106936
rect 213918 106584 213974 106593
rect 213918 106519 213974 106528
rect 213932 106350 213960 106519
rect 214024 106418 214052 106927
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 214010 105768 214066 105777
rect 214010 105703 214066 105712
rect 213918 105088 213974 105097
rect 213918 105023 213974 105032
rect 213932 104990 213960 105023
rect 213920 104984 213972 104990
rect 213920 104926 213972 104932
rect 214024 104922 214052 105703
rect 214012 104916 214064 104922
rect 214012 104858 214064 104864
rect 213918 103728 213974 103737
rect 213918 103663 213974 103672
rect 213932 103562 213960 103663
rect 213920 103556 213972 103562
rect 213920 103498 213972 103504
rect 213918 102504 213974 102513
rect 213918 102439 213974 102448
rect 213932 102202 213960 102439
rect 213920 102196 213972 102202
rect 213920 102138 213972 102144
rect 214010 101280 214066 101289
rect 214010 101215 214066 101224
rect 213918 101144 213974 101153
rect 213918 101079 213974 101088
rect 213932 100774 213960 101079
rect 214024 100842 214052 101215
rect 214012 100836 214064 100842
rect 214012 100778 214064 100784
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214010 99784 214066 99793
rect 214010 99719 214066 99728
rect 213918 99512 213974 99521
rect 213918 99447 213974 99456
rect 213932 99414 213960 99447
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214024 98666 214052 99719
rect 214012 98660 214064 98666
rect 214012 98602 214064 98608
rect 214010 98424 214066 98433
rect 214010 98359 214066 98368
rect 213920 98048 213972 98054
rect 213918 98016 213920 98025
rect 213972 98016 213974 98025
rect 213918 97951 213974 97960
rect 214024 94518 214052 98359
rect 214576 95946 214604 147999
rect 215036 145586 215064 151807
rect 215024 145580 215076 145586
rect 215024 145522 215076 145528
rect 214746 144936 214802 144945
rect 214746 144871 214802 144880
rect 214760 140078 214788 144871
rect 214748 140072 214800 140078
rect 214748 140014 214800 140020
rect 214654 139632 214710 139641
rect 214654 139567 214710 139576
rect 214668 139534 214696 139567
rect 214656 139528 214708 139534
rect 214656 139470 214708 139476
rect 214654 138136 214710 138145
rect 214654 138071 214710 138080
rect 214668 100065 214696 138071
rect 214838 102368 214894 102377
rect 214838 102303 214894 102312
rect 214654 100056 214710 100065
rect 214654 99991 214710 100000
rect 214654 97064 214710 97073
rect 214654 96999 214710 97008
rect 214564 95940 214616 95946
rect 214564 95882 214616 95888
rect 214012 94512 214064 94518
rect 214012 94454 214064 94460
rect 214668 84182 214696 96999
rect 214746 95840 214802 95849
rect 214746 95775 214802 95784
rect 214760 86970 214788 95775
rect 214852 93838 214880 102303
rect 214840 93832 214892 93838
rect 214840 93774 214892 93780
rect 214748 86964 214800 86970
rect 214748 86906 214800 86912
rect 214656 84176 214708 84182
rect 214656 84118 214708 84124
rect 213460 78668 213512 78674
rect 213460 78610 213512 78616
rect 213276 28348 213328 28354
rect 213276 28290 213328 28296
rect 215956 7682 215984 227015
rect 216036 214600 216088 214606
rect 216036 214542 216088 214548
rect 216048 25634 216076 214542
rect 217336 202434 217364 227734
rect 218716 222086 218744 237390
rect 218808 233034 218836 239822
rect 220648 237454 220676 240040
rect 223178 239850 223206 240040
rect 225110 239850 225138 240040
rect 222212 239822 223206 239850
rect 224972 239822 225138 239850
rect 220636 237448 220688 237454
rect 220636 237390 220688 237396
rect 218796 233028 218848 233034
rect 218796 232970 218848 232976
rect 218704 222080 218756 222086
rect 218704 222022 218756 222028
rect 217324 202428 217376 202434
rect 217324 202370 217376 202376
rect 218716 188494 218744 222022
rect 218808 209098 218836 232970
rect 222212 226302 222240 239822
rect 224224 234048 224276 234054
rect 224224 233990 224276 233996
rect 222200 226296 222252 226302
rect 222200 226238 222252 226244
rect 222212 225010 222240 226238
rect 222200 225004 222252 225010
rect 222200 224946 222252 224952
rect 222936 225004 222988 225010
rect 222936 224946 222988 224952
rect 218796 209092 218848 209098
rect 218796 209034 218848 209040
rect 222844 207936 222896 207942
rect 222844 207878 222896 207884
rect 218704 188488 218756 188494
rect 218704 188430 218756 188436
rect 216128 181756 216180 181762
rect 216128 181698 216180 181704
rect 216140 92478 216168 181698
rect 222856 180130 222884 207878
rect 222948 205018 222976 224946
rect 222936 205012 222988 205018
rect 222936 204954 222988 204960
rect 222844 180124 222896 180130
rect 222844 180066 222896 180072
rect 224236 175953 224264 233990
rect 224972 210526 225000 239822
rect 227088 235929 227116 240040
rect 229664 237454 229692 240040
rect 231550 239816 231578 240040
rect 233482 239816 233510 240040
rect 230492 239788 231578 239816
rect 233252 239788 233510 239816
rect 228548 237448 228600 237454
rect 228548 237390 228600 237396
rect 229652 237448 229704 237454
rect 229652 237390 229704 237396
rect 227074 235920 227130 235929
rect 227074 235855 227130 235864
rect 228364 233980 228416 233986
rect 228364 233922 228416 233928
rect 226984 231124 227036 231130
rect 226984 231066 227036 231072
rect 224960 210520 225012 210526
rect 224960 210462 225012 210468
rect 224972 209774 225000 210462
rect 224880 209746 225000 209774
rect 224880 192710 224908 209746
rect 224868 192704 224920 192710
rect 224868 192646 224920 192652
rect 226996 177614 227024 231066
rect 227076 218952 227128 218958
rect 227076 218894 227128 218900
rect 227088 184210 227116 218894
rect 227076 184204 227128 184210
rect 227076 184146 227128 184152
rect 228376 183122 228404 233922
rect 228456 221604 228508 221610
rect 228456 221546 228508 221552
rect 228364 183116 228416 183122
rect 228364 183058 228416 183064
rect 228468 181762 228496 221546
rect 228560 219366 228588 237390
rect 230492 220658 230520 239788
rect 231124 224324 231176 224330
rect 231124 224266 231176 224272
rect 230480 220652 230532 220658
rect 230480 220594 230532 220600
rect 228548 219360 228600 219366
rect 228548 219302 228600 219308
rect 228560 190126 228588 219302
rect 228548 190120 228600 190126
rect 228548 190062 228600 190068
rect 228456 181756 228508 181762
rect 228456 181698 228508 181704
rect 226984 177608 227036 177614
rect 226984 177550 227036 177556
rect 231136 177546 231164 224266
rect 232504 223032 232556 223038
rect 232504 222974 232556 222980
rect 231216 220652 231268 220658
rect 231216 220594 231268 220600
rect 231228 187202 231256 220594
rect 231216 187196 231268 187202
rect 231216 187138 231268 187144
rect 232516 180169 232544 222974
rect 233252 216578 233280 239788
rect 236104 237454 236132 240040
rect 237990 239816 238018 240040
rect 239922 239834 239950 240040
rect 237392 239788 238018 239816
rect 238760 239828 238812 239834
rect 235264 237448 235316 237454
rect 235264 237390 235316 237396
rect 236092 237448 236144 237454
rect 236092 237390 236144 237396
rect 233884 229900 233936 229906
rect 233884 229842 233936 229848
rect 233240 216572 233292 216578
rect 233240 216514 233292 216520
rect 233252 214606 233280 216514
rect 233240 214600 233292 214606
rect 233240 214542 233292 214548
rect 232596 202292 232648 202298
rect 232596 202234 232648 202240
rect 232608 184482 232636 202234
rect 232596 184476 232648 184482
rect 232596 184418 232648 184424
rect 233896 181626 233924 229842
rect 235276 227594 235304 237390
rect 235264 227588 235316 227594
rect 235264 227530 235316 227536
rect 235276 187338 235304 227530
rect 237392 221950 237420 239788
rect 238760 239770 238812 239776
rect 239910 239828 239962 239834
rect 239910 239770 239962 239776
rect 238772 223446 238800 239770
rect 241900 238754 241928 240040
rect 241900 238726 242204 238754
rect 241900 238678 241928 238726
rect 241888 238672 241940 238678
rect 241888 238614 241940 238620
rect 238760 223440 238812 223446
rect 238760 223382 238812 223388
rect 239404 223440 239456 223446
rect 239404 223382 239456 223388
rect 237380 221944 237432 221950
rect 237380 221886 237432 221892
rect 236644 218884 236696 218890
rect 236644 218826 236696 218832
rect 235264 187332 235316 187338
rect 235264 187274 235316 187280
rect 236656 183190 236684 218826
rect 237392 217394 237420 221886
rect 238208 217592 238260 217598
rect 238208 217534 238260 217540
rect 237380 217388 237432 217394
rect 237380 217330 237432 217336
rect 238024 208004 238076 208010
rect 238024 207946 238076 207952
rect 236644 183184 236696 183190
rect 236644 183126 236696 183132
rect 233884 181620 233936 181626
rect 233884 181562 233936 181568
rect 232502 180160 232558 180169
rect 232502 180095 232558 180104
rect 231124 177540 231176 177546
rect 231124 177482 231176 177488
rect 238036 175982 238064 207946
rect 238116 199504 238168 199510
rect 238116 199446 238168 199452
rect 238128 176118 238156 199446
rect 238220 196858 238248 217534
rect 239416 207670 239444 223382
rect 240784 214804 240836 214810
rect 240784 214746 240836 214752
rect 239404 207664 239456 207670
rect 239404 207606 239456 207612
rect 238208 196852 238260 196858
rect 238208 196794 238260 196800
rect 238116 176112 238168 176118
rect 238116 176054 238168 176060
rect 238024 175976 238076 175982
rect 224222 175944 224278 175953
rect 238024 175918 238076 175924
rect 224222 175879 224278 175888
rect 240796 175846 240824 214746
rect 240876 209296 240928 209302
rect 240876 209238 240928 209244
rect 240888 178809 240916 209238
rect 240968 204944 241020 204950
rect 240968 204886 241020 204892
rect 240980 185609 241008 204886
rect 242176 196790 242204 238726
rect 244476 238513 244504 240040
rect 244462 238504 244518 238513
rect 244462 238439 244518 238448
rect 246408 237454 246436 240040
rect 248294 239834 248322 240040
rect 247040 239828 247092 239834
rect 247040 239770 247092 239776
rect 248282 239828 248334 239834
rect 250870 239816 250898 240040
rect 248282 239770 248334 239776
rect 249812 239788 250898 239816
rect 244924 237448 244976 237454
rect 244924 237390 244976 237396
rect 246396 237448 246448 237454
rect 246396 237390 246448 237396
rect 244936 231538 244964 237390
rect 244924 231532 244976 231538
rect 244924 231474 244976 231480
rect 242256 200932 242308 200938
rect 242256 200874 242308 200880
rect 242164 196784 242216 196790
rect 242164 196726 242216 196732
rect 240966 185600 241022 185609
rect 240966 185535 241022 185544
rect 240874 178800 240930 178809
rect 240874 178735 240930 178744
rect 242268 177682 242296 200874
rect 243544 196716 243596 196722
rect 243544 196658 243596 196664
rect 243556 178945 243584 196658
rect 243542 178936 243598 178945
rect 244936 178906 244964 231474
rect 247052 220862 247080 239770
rect 247040 220856 247092 220862
rect 247040 220798 247092 220804
rect 247052 220726 247080 220798
rect 247040 220720 247092 220726
rect 247040 220662 247092 220668
rect 249064 217456 249116 217462
rect 249064 217398 249116 217404
rect 246304 213376 246356 213382
rect 246304 213318 246356 213324
rect 245016 210588 245068 210594
rect 245016 210530 245068 210536
rect 245028 181830 245056 210530
rect 245108 192772 245160 192778
rect 245108 192714 245160 192720
rect 245016 181824 245068 181830
rect 245016 181766 245068 181772
rect 243542 178871 243598 178880
rect 244924 178900 244976 178906
rect 244924 178842 244976 178848
rect 242256 177676 242308 177682
rect 242256 177618 242308 177624
rect 245120 176089 245148 192714
rect 246316 180470 246344 213318
rect 246304 180464 246356 180470
rect 246304 180406 246356 180412
rect 245106 176080 245162 176089
rect 245106 176015 245162 176024
rect 240784 175840 240836 175846
rect 248052 175840 248104 175846
rect 240784 175782 240836 175788
rect 248050 175808 248052 175817
rect 248104 175808 248106 175817
rect 248050 175743 248106 175752
rect 249076 171134 249104 217398
rect 249812 206990 249840 239788
rect 252848 238814 252876 240040
rect 252836 238808 252888 238814
rect 252834 238776 252836 238785
rect 252888 238776 252890 238785
rect 252834 238711 252890 238720
rect 254780 237454 254808 240040
rect 251640 237448 251692 237454
rect 251640 237390 251692 237396
rect 254768 237448 254820 237454
rect 254768 237390 254820 237396
rect 251652 235822 251680 237390
rect 251640 235816 251692 235822
rect 251640 235758 251692 235764
rect 251652 229094 251680 235758
rect 256712 234598 256740 240040
rect 259242 239834 259270 240040
rect 261174 239850 261202 240040
rect 263106 239850 263134 240040
rect 265682 239850 265710 240040
rect 258080 239828 258132 239834
rect 258080 239770 258132 239776
rect 259230 239828 259282 239834
rect 259230 239770 259282 239776
rect 260852 239822 261202 239850
rect 262232 239822 263134 239850
rect 265636 239822 265710 239850
rect 267614 239834 267642 240040
rect 266360 239828 266412 239834
rect 256700 234592 256752 234598
rect 256700 234534 256752 234540
rect 256712 234190 256740 234534
rect 256700 234184 256752 234190
rect 256700 234126 256752 234132
rect 257344 234184 257396 234190
rect 257344 234126 257396 234132
rect 255596 229764 255648 229770
rect 255596 229706 255648 229712
rect 251652 229066 251864 229094
rect 249892 217524 249944 217530
rect 249892 217466 249944 217472
rect 249800 206984 249852 206990
rect 249800 206926 249852 206932
rect 249800 187128 249852 187134
rect 249800 187070 249852 187076
rect 249156 181552 249208 181558
rect 249156 181494 249208 181500
rect 249168 175273 249196 181494
rect 249340 178764 249392 178770
rect 249340 178706 249392 178712
rect 249248 177608 249300 177614
rect 249248 177550 249300 177556
rect 249154 175264 249210 175273
rect 249154 175199 249210 175208
rect 249260 172825 249288 177550
rect 249246 172816 249302 172825
rect 249246 172751 249302 172760
rect 249352 171465 249380 178706
rect 249338 171456 249394 171465
rect 249338 171391 249394 171400
rect 249076 171106 249196 171134
rect 249168 161537 249196 171106
rect 249154 161528 249210 161537
rect 249154 161463 249210 161472
rect 249812 139505 249840 187070
rect 249904 149841 249932 217466
rect 250076 198144 250128 198150
rect 250076 198086 250128 198092
rect 250088 190454 250116 198086
rect 251180 198076 251232 198082
rect 251180 198018 251232 198024
rect 250088 190426 250300 190454
rect 249984 188420 250036 188426
rect 249984 188362 250036 188368
rect 249996 171134 250024 188362
rect 249996 171106 250116 171134
rect 250088 155417 250116 171106
rect 250272 169561 250300 190426
rect 250258 169552 250314 169561
rect 250258 169487 250314 169496
rect 251192 156369 251220 198018
rect 251836 181694 251864 229066
rect 251914 228304 251970 228313
rect 251914 228239 251970 228248
rect 251928 183054 251956 228239
rect 252836 227044 252888 227050
rect 252836 226986 252888 226992
rect 252006 225584 252062 225593
rect 252006 225519 252062 225528
rect 252020 188329 252048 225519
rect 252744 207800 252796 207806
rect 252744 207742 252796 207748
rect 252652 193928 252704 193934
rect 252652 193870 252704 193876
rect 252006 188320 252062 188329
rect 252006 188255 252062 188264
rect 251916 183048 251968 183054
rect 251916 182990 251968 182996
rect 251272 181688 251324 181694
rect 251272 181630 251324 181636
rect 251824 181688 251876 181694
rect 251824 181630 251876 181636
rect 251284 167278 251312 181630
rect 251364 180396 251416 180402
rect 251364 180338 251416 180344
rect 251272 167272 251324 167278
rect 251272 167214 251324 167220
rect 251376 159225 251404 180338
rect 251456 178968 251508 178974
rect 251456 178910 251508 178916
rect 251468 160177 251496 178910
rect 252468 175160 252520 175166
rect 252468 175102 252520 175108
rect 252480 174729 252508 175102
rect 252466 174720 252522 174729
rect 252466 174655 252522 174664
rect 252468 173868 252520 173874
rect 252468 173810 252520 173816
rect 252480 173777 252508 173810
rect 252466 173768 252522 173777
rect 252466 173703 252522 173712
rect 252376 172508 252428 172514
rect 252376 172450 252428 172456
rect 252388 171873 252416 172450
rect 252466 172408 252522 172417
rect 252466 172343 252522 172352
rect 252480 172174 252508 172343
rect 252468 172168 252520 172174
rect 252468 172110 252520 172116
rect 252374 171864 252430 171873
rect 252374 171799 252430 171808
rect 252468 171080 252520 171086
rect 252468 171022 252520 171028
rect 252376 171012 252428 171018
rect 252376 170954 252428 170960
rect 252388 170513 252416 170954
rect 252480 170921 252508 171022
rect 252466 170912 252522 170921
rect 252466 170847 252522 170856
rect 252468 170604 252520 170610
rect 252468 170546 252520 170552
rect 252374 170504 252430 170513
rect 252374 170439 252430 170448
rect 252480 170105 252508 170546
rect 252466 170096 252522 170105
rect 252466 170031 252522 170040
rect 252376 168360 252428 168366
rect 252376 168302 252428 168308
rect 251548 167272 251600 167278
rect 252388 167249 252416 168302
rect 252466 168192 252522 168201
rect 252466 168127 252522 168136
rect 252480 168094 252508 168127
rect 252468 168088 252520 168094
rect 252468 168030 252520 168036
rect 251548 167214 251600 167220
rect 252374 167240 252430 167249
rect 251454 160168 251510 160177
rect 251454 160103 251510 160112
rect 251362 159216 251418 159225
rect 251362 159151 251418 159160
rect 251560 156913 251588 167214
rect 252374 167175 252430 167184
rect 252376 166728 252428 166734
rect 252376 166670 252428 166676
rect 252466 166696 252522 166705
rect 252388 166297 252416 166670
rect 252466 166631 252468 166640
rect 252520 166631 252522 166640
rect 252468 166602 252520 166608
rect 252374 166288 252430 166297
rect 252374 166223 252430 166232
rect 252468 166116 252520 166122
rect 252468 166058 252520 166064
rect 252480 165753 252508 166058
rect 252466 165744 252522 165753
rect 252466 165679 252522 165688
rect 252468 165572 252520 165578
rect 252468 165514 252520 165520
rect 252376 165504 252428 165510
rect 252376 165446 252428 165452
rect 252388 164801 252416 165446
rect 252480 165345 252508 165514
rect 252466 165336 252522 165345
rect 252466 165271 252522 165280
rect 252374 164792 252430 164801
rect 252374 164727 252430 164736
rect 252468 164212 252520 164218
rect 252468 164154 252520 164160
rect 252376 164144 252428 164150
rect 252376 164086 252428 164092
rect 252388 163033 252416 164086
rect 252480 163985 252508 164154
rect 252466 163976 252522 163985
rect 252466 163911 252522 163920
rect 252374 163024 252430 163033
rect 252374 162959 252430 162968
rect 252376 162852 252428 162858
rect 252376 162794 252428 162800
rect 252388 162081 252416 162794
rect 252468 162784 252520 162790
rect 252468 162726 252520 162732
rect 252480 162489 252508 162726
rect 252466 162480 252522 162489
rect 252466 162415 252522 162424
rect 252374 162072 252430 162081
rect 252374 162007 252430 162016
rect 252468 161424 252520 161430
rect 252468 161366 252520 161372
rect 252480 160585 252508 161366
rect 252466 160576 252522 160585
rect 252376 160540 252428 160546
rect 252466 160511 252522 160520
rect 252376 160482 252428 160488
rect 252388 158273 252416 160482
rect 252468 160064 252520 160070
rect 252468 160006 252520 160012
rect 252480 159633 252508 160006
rect 252466 159624 252522 159633
rect 252466 159559 252522 159568
rect 252468 158704 252520 158710
rect 252468 158646 252520 158652
rect 252374 158264 252430 158273
rect 252374 158199 252430 158208
rect 252480 157865 252508 158646
rect 252466 157856 252522 157865
rect 252466 157791 252522 157800
rect 252468 157344 252520 157350
rect 252466 157312 252468 157321
rect 252520 157312 252522 157321
rect 252466 157247 252522 157256
rect 251546 156904 251602 156913
rect 251546 156839 251602 156848
rect 251178 156360 251234 156369
rect 251178 156295 251234 156304
rect 252374 155952 252430 155961
rect 252374 155887 252430 155896
rect 252468 155916 252520 155922
rect 252388 155854 252416 155887
rect 252468 155858 252520 155864
rect 252376 155848 252428 155854
rect 252376 155790 252428 155796
rect 250074 155408 250130 155417
rect 250074 155343 250130 155352
rect 252480 155009 252508 155858
rect 252466 155000 252522 155009
rect 252466 154935 252522 154944
rect 252468 154556 252520 154562
rect 252468 154498 252520 154504
rect 251456 154488 251508 154494
rect 252480 154465 252508 154498
rect 251456 154430 251508 154436
rect 252466 154456 252522 154465
rect 251468 153377 251496 154430
rect 252466 154391 252522 154400
rect 251454 153368 251510 153377
rect 251454 153303 251510 153312
rect 252284 153196 252336 153202
rect 252284 153138 252336 153144
rect 252296 152153 252324 153138
rect 252468 153128 252520 153134
rect 252466 153096 252468 153105
rect 252520 153096 252522 153105
rect 252376 153060 252428 153066
rect 252466 153031 252522 153040
rect 252376 153002 252428 153008
rect 252388 152697 252416 153002
rect 252374 152688 252430 152697
rect 252374 152623 252430 152632
rect 252282 152144 252338 152153
rect 252282 152079 252338 152088
rect 252664 151745 252692 193870
rect 252756 164393 252784 207742
rect 252848 169153 252876 226986
rect 255412 224256 255464 224262
rect 255412 224198 255464 224204
rect 254032 222964 254084 222970
rect 254032 222906 254084 222912
rect 253940 220108 253992 220114
rect 253940 220050 253992 220056
rect 252834 169144 252890 169153
rect 252834 169079 252890 169088
rect 252742 164384 252798 164393
rect 252742 164319 252798 164328
rect 253388 158024 253440 158030
rect 253388 157966 253440 157972
rect 253204 156664 253256 156670
rect 253204 156606 253256 156612
rect 252650 151736 252706 151745
rect 252650 151671 252706 151680
rect 252468 151496 252520 151502
rect 252468 151438 252520 151444
rect 251456 151360 251508 151366
rect 251456 151302 251508 151308
rect 251468 150793 251496 151302
rect 252480 151201 252508 151438
rect 252466 151192 252522 151201
rect 251824 151156 251876 151162
rect 252466 151127 252522 151136
rect 251824 151098 251876 151104
rect 251454 150784 251510 150793
rect 251454 150719 251510 150728
rect 251364 150340 251416 150346
rect 251364 150282 251416 150288
rect 249890 149832 249946 149841
rect 249890 149767 249946 149776
rect 251376 149297 251404 150282
rect 251362 149288 251418 149297
rect 251362 149223 251418 149232
rect 251364 147552 251416 147558
rect 251364 147494 251416 147500
rect 251376 146577 251404 147494
rect 251362 146568 251418 146577
rect 251362 146503 251418 146512
rect 249798 139496 249854 139505
rect 249798 139431 249854 139440
rect 250628 139460 250680 139466
rect 250628 139402 250680 139408
rect 250536 138032 250588 138038
rect 250536 137974 250588 137980
rect 250444 136672 250496 136678
rect 250444 136614 250496 136620
rect 216678 114608 216734 114617
rect 216678 114543 216734 114552
rect 216128 92472 216180 92478
rect 216128 92414 216180 92420
rect 216692 86902 216720 114543
rect 249064 113212 249116 113218
rect 249064 113154 249116 113160
rect 222844 96008 222896 96014
rect 222844 95950 222896 95956
rect 216680 86896 216732 86902
rect 216680 86838 216732 86844
rect 222856 37262 222884 95950
rect 242164 87644 242216 87650
rect 242164 87586 242216 87592
rect 238024 82136 238076 82142
rect 238024 82078 238076 82084
rect 232504 79416 232556 79422
rect 232504 79358 232556 79364
rect 226984 69760 227036 69766
rect 226984 69702 227036 69708
rect 222844 37256 222896 37262
rect 222844 37198 222896 37204
rect 216036 25628 216088 25634
rect 216036 25570 216088 25576
rect 226996 10334 227024 69702
rect 232516 38078 232544 79358
rect 232596 53100 232648 53106
rect 232596 53042 232648 53048
rect 232504 38072 232556 38078
rect 232504 38014 232556 38020
rect 232608 20058 232636 53042
rect 232596 20052 232648 20058
rect 232596 19994 232648 20000
rect 226984 10328 227036 10334
rect 226984 10270 227036 10276
rect 215944 7676 215996 7682
rect 215944 7618 215996 7624
rect 213184 4888 213236 4894
rect 213184 4830 213236 4836
rect 195428 3596 195480 3602
rect 195428 3538 195480 3544
rect 171966 3431 172022 3440
rect 188528 3460 188580 3466
rect 171980 480 172008 3431
rect 188528 3402 188580 3408
rect 238036 3126 238064 82078
rect 240784 50448 240836 50454
rect 240784 50390 240836 50396
rect 240796 6914 240824 50390
rect 240520 6886 240824 6914
rect 239220 4956 239272 4962
rect 239220 4898 239272 4904
rect 239232 4078 239260 4898
rect 239220 4072 239272 4078
rect 240520 4049 240548 6886
rect 242176 6866 242204 87586
rect 244280 86284 244332 86290
rect 244280 86226 244332 86232
rect 243544 51876 243596 51882
rect 243544 51818 243596 51824
rect 243556 10985 243584 51818
rect 244292 16574 244320 86226
rect 246304 79348 246356 79354
rect 246304 79290 246356 79296
rect 246316 31278 246344 79290
rect 246396 68332 246448 68338
rect 246396 68274 246448 68280
rect 246408 58886 246436 68274
rect 246396 58880 246448 58886
rect 246396 58822 246448 58828
rect 247960 53100 248012 53106
rect 247960 53042 248012 53048
rect 247972 51066 248000 53042
rect 247040 51060 247092 51066
rect 247040 51002 247092 51008
rect 247960 51060 248012 51066
rect 247960 51002 248012 51008
rect 246304 31272 246356 31278
rect 246304 31214 246356 31220
rect 246304 18624 246356 18630
rect 246304 18566 246356 18572
rect 244924 17400 244976 17406
rect 244924 17342 244976 17348
rect 244292 16546 244872 16574
rect 242898 10976 242954 10985
rect 242898 10911 242954 10920
rect 243542 10976 243598 10985
rect 243542 10911 243598 10920
rect 242164 6860 242216 6866
rect 242164 6802 242216 6808
rect 239220 4014 239272 4020
rect 240506 4040 240562 4049
rect 235816 3120 235868 3126
rect 235816 3062 235868 3068
rect 238024 3120 238076 3126
rect 238024 3062 238076 3068
rect 239232 3074 239260 4014
rect 240506 3975 240562 3984
rect 235828 480 235856 3062
rect 239232 3046 239352 3074
rect 239324 480 239352 3046
rect 240520 480 240548 3975
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 354 241786 480
rect 242176 354 242204 6802
rect 242912 3534 242940 10911
rect 242992 3596 243044 3602
rect 242992 3538 243044 3544
rect 242900 3528 242952 3534
rect 242900 3470 242952 3476
rect 243004 3369 243032 3538
rect 244096 3528 244148 3534
rect 244096 3470 244148 3476
rect 244844 3482 244872 16546
rect 244936 3602 244964 17342
rect 246316 16574 246344 18566
rect 247052 16574 247080 51002
rect 246316 16546 246436 16574
rect 247052 16546 247632 16574
rect 246408 4146 246436 16546
rect 246396 4140 246448 4146
rect 246396 4082 246448 4088
rect 244924 3596 244976 3602
rect 244924 3538 244976 3544
rect 242990 3360 243046 3369
rect 242912 3318 242990 3346
rect 242912 480 242940 3318
rect 242990 3295 243046 3304
rect 244108 480 244136 3470
rect 244844 3454 245240 3482
rect 245212 480 245240 3454
rect 246408 480 246436 4082
rect 247604 480 247632 16546
rect 248420 12504 248472 12510
rect 248420 12446 248472 12452
rect 241674 326 242204 354
rect 241674 -960 241786 326
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 354 248460 12446
rect 249076 8974 249104 113154
rect 249248 95260 249300 95266
rect 249248 95202 249300 95208
rect 249156 89684 249208 89690
rect 249156 89626 249208 89632
rect 249168 19310 249196 89626
rect 249260 51746 249288 95202
rect 249248 51740 249300 51746
rect 249248 51682 249300 51688
rect 250456 29714 250484 136614
rect 250548 43518 250576 137974
rect 250640 54534 250668 139402
rect 251180 126880 251232 126886
rect 251180 126822 251232 126828
rect 251192 125769 251220 126822
rect 251178 125760 251234 125769
rect 251178 125695 251234 125704
rect 251732 123480 251784 123486
rect 251732 123422 251784 123428
rect 251744 118833 251772 123422
rect 251730 118824 251786 118833
rect 251730 118759 251786 118768
rect 251836 117337 251864 151098
rect 252468 150408 252520 150414
rect 252468 150350 252520 150356
rect 252480 150249 252508 150350
rect 252466 150240 252522 150249
rect 252466 150175 252522 150184
rect 252468 149048 252520 149054
rect 252468 148990 252520 148996
rect 252376 148980 252428 148986
rect 252376 148922 252428 148928
rect 252388 148345 252416 148922
rect 252480 148889 252508 148990
rect 252466 148880 252522 148889
rect 252466 148815 252522 148824
rect 252374 148336 252430 148345
rect 252374 148271 252430 148280
rect 252468 147620 252520 147626
rect 252468 147562 252520 147568
rect 252480 147529 252508 147562
rect 252466 147520 252522 147529
rect 252100 147484 252152 147490
rect 252466 147455 252522 147464
rect 252100 147426 252152 147432
rect 252112 146985 252140 147426
rect 252098 146976 252154 146985
rect 252098 146911 252154 146920
rect 252376 146260 252428 146266
rect 252376 146202 252428 146208
rect 252388 145081 252416 146202
rect 252468 146192 252520 146198
rect 252468 146134 252520 146140
rect 252480 145625 252508 146134
rect 252466 145616 252522 145625
rect 252466 145551 252522 145560
rect 252374 145072 252430 145081
rect 252374 145007 252430 145016
rect 252376 144900 252428 144906
rect 252376 144842 252428 144848
rect 252388 143721 252416 144842
rect 252468 144832 252520 144838
rect 252468 144774 252520 144780
rect 252480 144129 252508 144774
rect 252466 144120 252522 144129
rect 252466 144055 252522 144064
rect 252374 143712 252430 143721
rect 251916 143676 251968 143682
rect 252374 143647 252430 143656
rect 251916 143618 251968 143624
rect 251928 121145 251956 143618
rect 252468 143540 252520 143546
rect 252468 143482 252520 143488
rect 252376 143472 252428 143478
rect 252376 143414 252428 143420
rect 252388 142769 252416 143414
rect 252480 143177 252508 143482
rect 252466 143168 252522 143177
rect 252466 143103 252522 143112
rect 252374 142760 252430 142769
rect 252374 142695 252430 142704
rect 252192 141500 252244 141506
rect 252192 141442 252244 141448
rect 252204 135289 252232 141442
rect 253216 140865 253244 156606
rect 253296 142860 253348 142866
rect 253296 142802 253348 142808
rect 253202 140856 253258 140865
rect 253202 140791 253258 140800
rect 252468 140752 252520 140758
rect 252468 140694 252520 140700
rect 252480 139913 252508 140694
rect 252466 139904 252522 139913
rect 252466 139839 252522 139848
rect 252468 139392 252520 139398
rect 252468 139334 252520 139340
rect 252480 138553 252508 139334
rect 252466 138544 252522 138553
rect 252466 138479 252522 138488
rect 253204 138100 253256 138106
rect 253204 138042 253256 138048
rect 252468 137964 252520 137970
rect 252468 137906 252520 137912
rect 252480 136785 252508 137906
rect 252466 136776 252522 136785
rect 252466 136711 252522 136720
rect 252466 136640 252522 136649
rect 252284 136604 252336 136610
rect 252466 136575 252522 136584
rect 252284 136546 252336 136552
rect 252296 136241 252324 136546
rect 252480 136542 252508 136575
rect 252468 136536 252520 136542
rect 252468 136478 252520 136484
rect 252376 136468 252428 136474
rect 252376 136410 252428 136416
rect 252282 136232 252338 136241
rect 252282 136167 252338 136176
rect 252388 135697 252416 136410
rect 252374 135688 252430 135697
rect 252374 135623 252430 135632
rect 252190 135280 252246 135289
rect 252190 135215 252246 135224
rect 252376 135244 252428 135250
rect 252376 135186 252428 135192
rect 252388 134337 252416 135186
rect 252468 135176 252520 135182
rect 252468 135118 252520 135124
rect 252480 134745 252508 135118
rect 252466 134736 252522 134745
rect 252466 134671 252522 134680
rect 252374 134328 252430 134337
rect 252374 134263 252430 134272
rect 252468 133884 252520 133890
rect 252468 133826 252520 133832
rect 252284 133816 252336 133822
rect 252480 133793 252508 133826
rect 252284 133758 252336 133764
rect 252466 133784 252522 133793
rect 252296 133385 252324 133758
rect 252376 133748 252428 133754
rect 252466 133719 252522 133728
rect 252376 133690 252428 133696
rect 252282 133376 252338 133385
rect 252282 133311 252338 133320
rect 252388 132841 252416 133690
rect 252374 132832 252430 132841
rect 252374 132767 252430 132776
rect 252284 132456 252336 132462
rect 252284 132398 252336 132404
rect 252466 132424 252522 132433
rect 252296 131889 252324 132398
rect 252466 132359 252468 132368
rect 252520 132359 252522 132368
rect 252468 132330 252520 132336
rect 252376 132320 252428 132326
rect 252376 132262 252428 132268
rect 252282 131880 252338 131889
rect 252282 131815 252338 131824
rect 252388 131481 252416 132262
rect 252374 131472 252430 131481
rect 252374 131407 252430 131416
rect 252468 131096 252520 131102
rect 252468 131038 252520 131044
rect 252376 131028 252428 131034
rect 252376 130970 252428 130976
rect 252388 130529 252416 130970
rect 252480 130937 252508 131038
rect 252466 130928 252522 130937
rect 252466 130863 252522 130872
rect 252374 130520 252430 130529
rect 252374 130455 252430 130464
rect 252468 130212 252520 130218
rect 252468 130154 252520 130160
rect 252480 130121 252508 130154
rect 252466 130112 252522 130121
rect 252466 130047 252522 130056
rect 252284 129736 252336 129742
rect 252284 129678 252336 129684
rect 252296 129169 252324 129678
rect 252468 129668 252520 129674
rect 252468 129610 252520 129616
rect 252376 129600 252428 129606
rect 252480 129577 252508 129610
rect 252376 129542 252428 129548
rect 252466 129568 252522 129577
rect 252282 129160 252338 129169
rect 252282 129095 252338 129104
rect 252388 128625 252416 129542
rect 252466 129503 252522 129512
rect 252374 128616 252430 128625
rect 252374 128551 252430 128560
rect 252376 128308 252428 128314
rect 252376 128250 252428 128256
rect 252282 128208 252338 128217
rect 252282 128143 252284 128152
rect 252336 128143 252338 128152
rect 252284 128114 252336 128120
rect 252192 127628 252244 127634
rect 252192 127570 252244 127576
rect 252100 125588 252152 125594
rect 252100 125530 252152 125536
rect 252112 125361 252140 125530
rect 252098 125352 252154 125361
rect 252098 125287 252154 125296
rect 252204 124001 252232 127570
rect 252388 127265 252416 128250
rect 252468 128240 252520 128246
rect 252468 128182 252520 128188
rect 252480 127673 252508 128182
rect 252466 127664 252522 127673
rect 252466 127599 252522 127608
rect 252374 127256 252430 127265
rect 252374 127191 252430 127200
rect 252468 126948 252520 126954
rect 252468 126890 252520 126896
rect 252480 126721 252508 126890
rect 252466 126712 252522 126721
rect 252466 126647 252522 126656
rect 252468 126472 252520 126478
rect 252468 126414 252520 126420
rect 252480 126313 252508 126414
rect 252466 126304 252522 126313
rect 252284 126268 252336 126274
rect 252466 126239 252522 126248
rect 252284 126210 252336 126216
rect 252190 123992 252246 124001
rect 252190 123927 252246 123936
rect 252296 123049 252324 126210
rect 252468 125520 252520 125526
rect 252468 125462 252520 125468
rect 252376 125452 252428 125458
rect 252376 125394 252428 125400
rect 252388 124409 252416 125394
rect 252480 124817 252508 125462
rect 252466 124808 252522 124817
rect 252466 124743 252522 124752
rect 252374 124400 252430 124409
rect 252374 124335 252430 124344
rect 252468 124160 252520 124166
rect 252468 124102 252520 124108
rect 252480 123457 252508 124102
rect 252466 123448 252522 123457
rect 252466 123383 252522 123392
rect 252282 123040 252338 123049
rect 252282 122975 252338 122984
rect 252468 122800 252520 122806
rect 252468 122742 252520 122748
rect 252376 122732 252428 122738
rect 252376 122674 252428 122680
rect 252284 122664 252336 122670
rect 252284 122606 252336 122612
rect 252296 121553 252324 122606
rect 252388 122097 252416 122674
rect 252480 122505 252508 122742
rect 252466 122496 252522 122505
rect 252466 122431 252522 122440
rect 252374 122088 252430 122097
rect 252374 122023 252430 122032
rect 252282 121544 252338 121553
rect 252282 121479 252338 121488
rect 252468 121440 252520 121446
rect 252468 121382 252520 121388
rect 251914 121136 251970 121145
rect 251914 121071 251970 121080
rect 252480 120601 252508 121382
rect 252466 120592 252522 120601
rect 252466 120527 252522 120536
rect 252468 120352 252520 120358
rect 252468 120294 252520 120300
rect 252480 120193 252508 120294
rect 252466 120184 252522 120193
rect 252466 120119 252522 120128
rect 252468 120080 252520 120086
rect 252468 120022 252520 120028
rect 252480 119649 252508 120022
rect 252466 119640 252522 119649
rect 252466 119575 252522 119584
rect 251916 119400 251968 119406
rect 251916 119342 251968 119348
rect 251822 117328 251878 117337
rect 251822 117263 251878 117272
rect 251732 108928 251784 108934
rect 251732 108870 251784 108876
rect 251744 107953 251772 108870
rect 251824 108384 251876 108390
rect 251824 108326 251876 108332
rect 251730 107944 251786 107953
rect 251730 107879 251786 107888
rect 251732 107568 251784 107574
rect 251732 107510 251784 107516
rect 251744 106593 251772 107510
rect 251730 106584 251786 106593
rect 251730 106519 251786 106528
rect 250720 106344 250772 106350
rect 250720 106286 250772 106292
rect 250628 54528 250680 54534
rect 250628 54470 250680 54476
rect 250732 50522 250760 106286
rect 251364 102060 251416 102066
rect 251364 102002 251416 102008
rect 251376 101833 251404 102002
rect 251362 101824 251418 101833
rect 251362 101759 251418 101768
rect 251836 100881 251864 108326
rect 251822 100872 251878 100881
rect 251822 100807 251878 100816
rect 251928 98569 251956 119342
rect 252466 119232 252522 119241
rect 252466 119167 252522 119176
rect 252480 118998 252508 119167
rect 252468 118992 252520 118998
rect 252468 118934 252520 118940
rect 252468 118652 252520 118658
rect 252468 118594 252520 118600
rect 252376 118584 252428 118590
rect 252376 118526 252428 118532
rect 252100 117972 252152 117978
rect 252100 117914 252152 117920
rect 252112 113121 252140 117914
rect 252388 117881 252416 118526
rect 252480 118289 252508 118594
rect 252466 118280 252522 118289
rect 252466 118215 252522 118224
rect 252374 117872 252430 117881
rect 252374 117807 252430 117816
rect 252376 117292 252428 117298
rect 252376 117234 252428 117240
rect 252284 117224 252336 117230
rect 252284 117166 252336 117172
rect 252296 115977 252324 117166
rect 252388 116929 252416 117234
rect 252374 116920 252430 116929
rect 252374 116855 252430 116864
rect 252468 116884 252520 116890
rect 252468 116826 252520 116832
rect 252480 116385 252508 116826
rect 252466 116376 252522 116385
rect 252466 116311 252522 116320
rect 252282 115968 252338 115977
rect 252282 115903 252338 115912
rect 252468 115932 252520 115938
rect 252468 115874 252520 115880
rect 252376 115864 252428 115870
rect 252376 115806 252428 115812
rect 252388 115025 252416 115806
rect 252480 115433 252508 115874
rect 252466 115424 252522 115433
rect 252466 115359 252522 115368
rect 252374 115016 252430 115025
rect 252374 114951 252430 114960
rect 252376 114572 252428 114578
rect 252376 114514 252428 114520
rect 252388 113529 252416 114514
rect 252468 114504 252520 114510
rect 252468 114446 252520 114452
rect 252480 114073 252508 114446
rect 252466 114064 252522 114073
rect 252466 113999 252522 114008
rect 252468 113824 252520 113830
rect 252468 113766 252520 113772
rect 252374 113520 252430 113529
rect 252374 113455 252430 113464
rect 252480 113174 252508 113766
rect 252388 113146 252508 113174
rect 252098 113112 252154 113121
rect 252098 113047 252154 113056
rect 252100 112532 252152 112538
rect 252100 112474 252152 112480
rect 252112 107001 252140 112474
rect 252192 112464 252244 112470
rect 252192 112406 252244 112412
rect 252204 108361 252232 112406
rect 252282 111752 252338 111761
rect 252282 111687 252284 111696
rect 252336 111687 252338 111696
rect 252284 111658 252336 111664
rect 252388 111217 252416 113146
rect 252468 112940 252520 112946
rect 252468 112882 252520 112888
rect 252480 112713 252508 112882
rect 252466 112704 252522 112713
rect 252466 112639 252522 112648
rect 252466 112160 252522 112169
rect 252466 112095 252522 112104
rect 252480 111926 252508 112095
rect 252468 111920 252520 111926
rect 252468 111862 252520 111868
rect 252468 111784 252520 111790
rect 252468 111726 252520 111732
rect 252374 111208 252430 111217
rect 252374 111143 252430 111152
rect 252480 110809 252508 111726
rect 252466 110800 252522 110809
rect 252466 110735 252522 110744
rect 252284 110424 252336 110430
rect 252284 110366 252336 110372
rect 252296 109313 252324 110366
rect 252376 110356 252428 110362
rect 252376 110298 252428 110304
rect 252388 109857 252416 110298
rect 252468 110288 252520 110294
rect 252466 110256 252468 110265
rect 252520 110256 252522 110265
rect 252466 110191 252522 110200
rect 252374 109848 252430 109857
rect 252374 109783 252430 109792
rect 252282 109304 252338 109313
rect 252282 109239 252338 109248
rect 252468 108996 252520 109002
rect 252468 108938 252520 108944
rect 252480 108905 252508 108938
rect 252466 108896 252522 108905
rect 252466 108831 252522 108840
rect 252190 108352 252246 108361
rect 252190 108287 252246 108296
rect 252468 107636 252520 107642
rect 252468 107578 252520 107584
rect 252480 107545 252508 107578
rect 252466 107536 252522 107545
rect 252466 107471 252522 107480
rect 252098 106992 252154 107001
rect 252098 106927 252154 106936
rect 252376 106276 252428 106282
rect 252376 106218 252428 106224
rect 252284 106140 252336 106146
rect 252284 106082 252336 106088
rect 252296 105097 252324 106082
rect 252388 105641 252416 106218
rect 252468 106208 252520 106214
rect 252468 106150 252520 106156
rect 252480 106049 252508 106150
rect 252466 106040 252522 106049
rect 252466 105975 252522 105984
rect 252374 105632 252430 105641
rect 252374 105567 252430 105576
rect 252282 105088 252338 105097
rect 252282 105023 252338 105032
rect 252376 104848 252428 104854
rect 252376 104790 252428 104796
rect 252284 104712 252336 104718
rect 252284 104654 252336 104660
rect 252296 104145 252324 104654
rect 252282 104136 252338 104145
rect 252282 104071 252338 104080
rect 252388 103737 252416 104790
rect 252468 104780 252520 104786
rect 252468 104722 252520 104728
rect 252480 104689 252508 104722
rect 252466 104680 252522 104689
rect 252466 104615 252522 104624
rect 252374 103728 252430 103737
rect 252374 103663 252430 103672
rect 252468 103488 252520 103494
rect 252468 103430 252520 103436
rect 252480 103193 252508 103430
rect 252466 103184 252522 103193
rect 252466 103119 252522 103128
rect 252376 103080 252428 103086
rect 252376 103022 252428 103028
rect 252388 102241 252416 103022
rect 252468 102944 252520 102950
rect 252468 102886 252520 102892
rect 252480 102785 252508 102886
rect 252466 102776 252522 102785
rect 252466 102711 252522 102720
rect 252374 102232 252430 102241
rect 252374 102167 252430 102176
rect 252468 102128 252520 102134
rect 252468 102070 252520 102076
rect 252192 101448 252244 101454
rect 252480 101425 252508 102070
rect 252192 101390 252244 101396
rect 252466 101416 252522 101425
rect 251914 98560 251970 98569
rect 251914 98495 251970 98504
rect 252204 98025 252232 101390
rect 252466 101351 252522 101360
rect 252376 100700 252428 100706
rect 252376 100642 252428 100648
rect 252284 100632 252336 100638
rect 252284 100574 252336 100580
rect 252296 99521 252324 100574
rect 252388 99929 252416 100642
rect 252468 100564 252520 100570
rect 252468 100506 252520 100512
rect 252480 100473 252508 100506
rect 252466 100464 252522 100473
rect 252466 100399 252522 100408
rect 252374 99920 252430 99929
rect 252374 99855 252430 99864
rect 252282 99512 252338 99521
rect 252282 99447 252338 99456
rect 252468 99340 252520 99346
rect 252468 99282 252520 99288
rect 252480 98977 252508 99282
rect 252466 98968 252522 98977
rect 252466 98903 252522 98912
rect 252468 98660 252520 98666
rect 252468 98602 252520 98608
rect 252190 98016 252246 98025
rect 252190 97951 252246 97960
rect 252480 97617 252508 98602
rect 252466 97608 252522 97617
rect 252466 97543 252522 97552
rect 252468 96756 252520 96762
rect 252468 96698 252520 96704
rect 251824 96688 251876 96694
rect 252480 96665 252508 96698
rect 251824 96630 251876 96636
rect 252466 96656 252522 96665
rect 251178 96248 251234 96257
rect 251178 96183 251234 96192
rect 251192 82142 251220 96183
rect 251362 82240 251418 82249
rect 251362 82175 251418 82184
rect 251180 82136 251232 82142
rect 251180 82078 251232 82084
rect 250720 50516 250772 50522
rect 250720 50458 250772 50464
rect 250536 43512 250588 43518
rect 250536 43454 250588 43460
rect 250444 29708 250496 29714
rect 250444 29650 250496 29656
rect 249800 20052 249852 20058
rect 249800 19994 249852 20000
rect 249246 19952 249302 19961
rect 249246 19887 249302 19896
rect 249156 19304 249208 19310
rect 249156 19246 249208 19252
rect 249260 13734 249288 19887
rect 249812 16574 249840 19994
rect 251376 16574 251404 82175
rect 251836 46306 251864 96630
rect 252466 96591 252522 96600
rect 251916 54528 251968 54534
rect 251916 54470 251968 54476
rect 251824 46300 251876 46306
rect 251824 46242 251876 46248
rect 249812 16546 250024 16574
rect 251376 16546 251864 16574
rect 249248 13728 249300 13734
rect 249248 13670 249300 13676
rect 249260 12510 249288 13670
rect 249248 12504 249300 12510
rect 249248 12446 249300 12452
rect 249064 8968 249116 8974
rect 249064 8910 249116 8916
rect 249996 480 250024 16546
rect 251180 5500 251232 5506
rect 251180 5442 251232 5448
rect 251192 5030 251220 5442
rect 251180 5024 251232 5030
rect 251180 4966 251232 4972
rect 251192 480 251220 4966
rect 251836 3482 251864 16546
rect 251928 5030 251956 54470
rect 253216 40798 253244 138042
rect 253308 102066 253336 142802
rect 253400 126886 253428 157966
rect 253952 147558 253980 220050
rect 254044 150346 254072 222906
rect 254124 203652 254176 203658
rect 254124 203594 254176 203600
rect 254136 151366 254164 203594
rect 254216 195424 254268 195430
rect 254216 195366 254268 195372
rect 254228 154494 254256 195366
rect 255424 155854 255452 224198
rect 255504 206440 255556 206446
rect 255504 206382 255556 206388
rect 255412 155848 255464 155854
rect 255412 155790 255464 155796
rect 254216 154488 254268 154494
rect 254216 154430 254268 154436
rect 254584 151836 254636 151842
rect 254584 151778 254636 151784
rect 254124 151360 254176 151366
rect 254124 151302 254176 151308
rect 254032 150340 254084 150346
rect 254032 150282 254084 150288
rect 253940 147552 253992 147558
rect 253940 147494 253992 147500
rect 253478 141808 253534 141817
rect 253478 141743 253534 141752
rect 253492 141001 253520 141743
rect 253572 141432 253624 141438
rect 253572 141374 253624 141380
rect 253478 140992 253534 141001
rect 253478 140927 253534 140936
rect 253388 126880 253440 126886
rect 253388 126822 253440 126828
rect 253584 125594 253612 141374
rect 253572 125588 253624 125594
rect 253572 125530 253624 125536
rect 254596 111722 254624 151778
rect 254860 149116 254912 149122
rect 254860 149058 254912 149064
rect 254768 147688 254820 147694
rect 254768 147630 254820 147636
rect 254676 135312 254728 135318
rect 254676 135254 254728 135260
rect 254584 111716 254636 111722
rect 254584 111658 254636 111664
rect 253388 110492 253440 110498
rect 253388 110434 253440 110440
rect 253296 102060 253348 102066
rect 253296 102002 253348 102008
rect 253296 86352 253348 86358
rect 253296 86294 253348 86300
rect 253204 40792 253256 40798
rect 253204 40734 253256 40740
rect 253308 22098 253336 86294
rect 253400 72554 253428 110434
rect 254584 106412 254636 106418
rect 254584 106354 254636 106360
rect 253388 72548 253440 72554
rect 253388 72490 253440 72496
rect 253296 22092 253348 22098
rect 253296 22034 253348 22040
rect 253308 21622 253336 22034
rect 252560 21616 252612 21622
rect 252560 21558 252612 21564
rect 253296 21616 253348 21622
rect 253296 21558 253348 21564
rect 252572 16574 252600 21558
rect 254596 17474 254624 106354
rect 254688 47666 254716 135254
rect 254780 107574 254808 147630
rect 254872 108934 254900 149058
rect 255516 147490 255544 206382
rect 255608 151502 255636 229706
rect 256976 211948 257028 211954
rect 256976 211890 257028 211896
rect 256792 188352 256844 188358
rect 256792 188294 256844 188300
rect 256700 176112 256752 176118
rect 256700 176054 256752 176060
rect 256712 170610 256740 176054
rect 256700 170604 256752 170610
rect 256700 170546 256752 170552
rect 256804 165510 256832 188294
rect 256884 177676 256936 177682
rect 256884 177618 256936 177624
rect 256896 168366 256924 177618
rect 256884 168360 256936 168366
rect 256884 168302 256936 168308
rect 256792 165504 256844 165510
rect 256792 165446 256844 165452
rect 255596 151496 255648 151502
rect 255596 151438 255648 151444
rect 255964 151088 256016 151094
rect 255964 151030 256016 151036
rect 255504 147484 255556 147490
rect 255504 147426 255556 147432
rect 255976 112946 256004 151030
rect 256988 148986 257016 211890
rect 257356 178770 257384 234126
rect 258092 224874 258120 239770
rect 258080 224868 258132 224874
rect 258080 224810 258132 224816
rect 258724 224868 258776 224874
rect 258724 224810 258776 224816
rect 258264 213308 258316 213314
rect 258264 213250 258316 213256
rect 258172 190052 258224 190058
rect 258172 189994 258224 190000
rect 257344 178764 257396 178770
rect 257344 178706 257396 178712
rect 258080 176044 258132 176050
rect 258080 175986 258132 175992
rect 258092 172174 258120 175986
rect 258184 175166 258212 189994
rect 258172 175160 258224 175166
rect 258172 175102 258224 175108
rect 258080 172168 258132 172174
rect 258080 172110 258132 172116
rect 258276 166734 258304 213250
rect 258736 211954 258764 224810
rect 259460 220244 259512 220250
rect 259460 220186 259512 220192
rect 258724 211948 258776 211954
rect 258724 211890 258776 211896
rect 258356 177540 258408 177546
rect 258356 177482 258408 177488
rect 258264 166728 258316 166734
rect 258264 166670 258316 166676
rect 258368 166666 258396 177482
rect 259000 168428 259052 168434
rect 259000 168370 259052 168376
rect 258356 166660 258408 166666
rect 258356 166602 258408 166608
rect 258724 164892 258776 164898
rect 258724 164834 258776 164840
rect 257620 163532 257672 163538
rect 257620 163474 257672 163480
rect 257344 157412 257396 157418
rect 257344 157354 257396 157360
rect 256976 148980 257028 148986
rect 256976 148922 257028 148928
rect 256148 144968 256200 144974
rect 256148 144910 256200 144916
rect 256056 143608 256108 143614
rect 256056 143550 256108 143556
rect 255964 112940 256016 112946
rect 255964 112882 256016 112888
rect 254860 108928 254912 108934
rect 254860 108870 254912 108876
rect 255964 107908 256016 107914
rect 255964 107850 256016 107856
rect 254768 107568 254820 107574
rect 254768 107510 254820 107516
rect 254768 83496 254820 83502
rect 254768 83438 254820 83444
rect 254780 55826 254808 83438
rect 254768 55820 254820 55826
rect 254768 55762 254820 55768
rect 254676 47660 254728 47666
rect 254676 47602 254728 47608
rect 254584 17468 254636 17474
rect 254584 17410 254636 17416
rect 252572 16546 253520 16574
rect 251916 5024 251968 5030
rect 251916 4966 251968 4972
rect 251836 3454 252416 3482
rect 252388 480 252416 3454
rect 253492 480 253520 16546
rect 254780 6914 254808 55762
rect 255976 31210 256004 107850
rect 256068 103086 256096 143550
rect 256160 104718 256188 144910
rect 256240 142180 256292 142186
rect 256240 142122 256292 142128
rect 256252 108390 256280 142122
rect 257356 118590 257384 157354
rect 257528 146328 257580 146334
rect 257528 146270 257580 146276
rect 257434 145616 257490 145625
rect 257434 145551 257490 145560
rect 257344 118584 257396 118590
rect 257344 118526 257396 118532
rect 256240 108384 256292 108390
rect 256240 108326 256292 108332
rect 257344 104916 257396 104922
rect 257344 104858 257396 104864
rect 256148 104712 256200 104718
rect 256148 104654 256200 104660
rect 256056 103080 256108 103086
rect 256056 103022 256108 103028
rect 256056 98048 256108 98054
rect 256056 97990 256108 97996
rect 256068 55894 256096 97990
rect 256700 97980 256752 97986
rect 256700 97922 256752 97928
rect 256712 96762 256740 97922
rect 256700 96756 256752 96762
rect 256700 96698 256752 96704
rect 256712 89690 256740 96698
rect 256700 89684 256752 89690
rect 256700 89626 256752 89632
rect 256056 55888 256108 55894
rect 256056 55830 256108 55836
rect 255964 31204 256016 31210
rect 255964 31146 256016 31152
rect 257356 21554 257384 104858
rect 257448 97986 257476 145551
rect 257540 106146 257568 146270
rect 257632 128178 257660 163474
rect 257620 128172 257672 128178
rect 257620 128114 257672 128120
rect 258736 126478 258764 164834
rect 258816 153332 258868 153338
rect 258816 153274 258868 153280
rect 258724 126472 258776 126478
rect 258724 126414 258776 126420
rect 258724 116000 258776 116006
rect 258724 115942 258776 115948
rect 257528 106140 257580 106146
rect 257528 106082 257580 106088
rect 257436 97980 257488 97986
rect 257436 97922 257488 97928
rect 257436 87712 257488 87718
rect 257436 87654 257488 87660
rect 257344 21548 257396 21554
rect 257344 21490 257396 21496
rect 255872 11824 255924 11830
rect 255872 11766 255924 11772
rect 254688 6886 254808 6914
rect 254688 480 254716 6886
rect 255884 480 255912 11766
rect 257448 5506 257476 87654
rect 258736 44878 258764 115942
rect 258828 111926 258856 153274
rect 258908 153264 258960 153270
rect 258908 153206 258960 153212
rect 258920 114578 258948 153206
rect 259012 130218 259040 168370
rect 259472 168094 259500 220186
rect 260852 208350 260880 239822
rect 262232 228818 262260 239822
rect 265636 233073 265664 239822
rect 266360 239770 266412 239776
rect 267602 239828 267654 239834
rect 269546 239816 269574 240040
rect 272122 239816 272150 240040
rect 274054 239816 274082 240040
rect 267602 239770 267654 239776
rect 269132 239788 269574 239816
rect 271892 239788 272150 239816
rect 273272 239788 274082 239816
rect 265622 233064 265678 233073
rect 265622 232999 265678 233008
rect 262864 229832 262916 229838
rect 262864 229774 262916 229780
rect 262220 228812 262272 228818
rect 262220 228754 262272 228760
rect 262232 227798 262260 228754
rect 262220 227792 262272 227798
rect 262220 227734 262272 227740
rect 260840 208344 260892 208350
rect 260840 208286 260892 208292
rect 260852 207126 260880 208286
rect 260840 207120 260892 207126
rect 260840 207062 260892 207068
rect 261484 207120 261536 207126
rect 261484 207062 261536 207068
rect 260932 199572 260984 199578
rect 260932 199514 260984 199520
rect 260840 189916 260892 189922
rect 260840 189858 260892 189864
rect 259552 185836 259604 185842
rect 259552 185778 259604 185784
rect 259460 168088 259512 168094
rect 259460 168030 259512 168036
rect 259564 165578 259592 185778
rect 259736 181756 259788 181762
rect 259736 181698 259788 181704
rect 259642 176080 259698 176089
rect 259642 176015 259698 176024
rect 259552 165572 259604 165578
rect 259552 165514 259604 165520
rect 259656 160546 259684 176015
rect 259748 166122 259776 181698
rect 259736 166116 259788 166122
rect 259736 166058 259788 166064
rect 259644 160540 259696 160546
rect 259644 160482 259696 160488
rect 260472 160200 260524 160206
rect 260472 160142 260524 160148
rect 260104 160132 260156 160138
rect 260104 160074 260156 160080
rect 260116 143682 260144 160074
rect 260380 158772 260432 158778
rect 260380 158714 260432 158720
rect 260288 155984 260340 155990
rect 260288 155926 260340 155932
rect 260104 143676 260156 143682
rect 260104 143618 260156 143624
rect 260196 143676 260248 143682
rect 260196 143618 260248 143624
rect 259000 130212 259052 130218
rect 259000 130154 259052 130160
rect 260104 120148 260156 120154
rect 260104 120090 260156 120096
rect 258908 114572 258960 114578
rect 258908 114514 258960 114520
rect 258816 111920 258868 111926
rect 258816 111862 258868 111868
rect 258908 102196 258960 102202
rect 258908 102138 258960 102144
rect 258920 55962 258948 102138
rect 259458 60752 259514 60761
rect 259458 60687 259514 60696
rect 258908 55956 258960 55962
rect 258908 55898 258960 55904
rect 258724 44872 258776 44878
rect 258724 44814 258776 44820
rect 258264 10328 258316 10334
rect 258264 10270 258316 10276
rect 257068 5500 257120 5506
rect 257068 5442 257120 5448
rect 257436 5500 257488 5506
rect 257436 5442 257488 5448
rect 257080 480 257108 5442
rect 258276 480 258304 10270
rect 259472 480 259500 60687
rect 260116 22914 260144 120090
rect 260208 102950 260236 143618
rect 260300 116890 260328 155926
rect 260392 118998 260420 158714
rect 260484 120358 260512 160142
rect 260852 146198 260880 189858
rect 260944 158710 260972 199514
rect 261496 199510 261524 207062
rect 262220 202360 262272 202366
rect 262220 202302 262272 202308
rect 261484 199504 261536 199510
rect 261484 199446 261536 199452
rect 261024 187264 261076 187270
rect 261024 187206 261076 187212
rect 261036 172514 261064 187206
rect 261024 172508 261076 172514
rect 261024 172450 261076 172456
rect 261484 171828 261536 171834
rect 261484 171770 261536 171776
rect 260932 158704 260984 158710
rect 260932 158646 260984 158652
rect 260840 146192 260892 146198
rect 260840 146134 260892 146140
rect 260472 120352 260524 120358
rect 260472 120294 260524 120300
rect 260380 118992 260432 118998
rect 260380 118934 260432 118940
rect 260288 116884 260340 116890
rect 260288 116826 260340 116832
rect 260196 102944 260248 102950
rect 260196 102886 260248 102892
rect 261496 99346 261524 171770
rect 261668 169788 261720 169794
rect 261668 169730 261720 169736
rect 261680 131034 261708 169730
rect 261760 154624 261812 154630
rect 261760 154566 261812 154572
rect 261668 131028 261720 131034
rect 261668 130970 261720 130976
rect 261576 129804 261628 129810
rect 261576 129746 261628 129752
rect 261484 99340 261536 99346
rect 261484 99282 261536 99288
rect 261482 84824 261538 84833
rect 261482 84759 261538 84768
rect 260194 79384 260250 79393
rect 260194 79319 260250 79328
rect 260208 62121 260236 79319
rect 260194 62112 260250 62121
rect 260194 62047 260250 62056
rect 260208 60761 260236 62047
rect 260194 60752 260250 60761
rect 260194 60687 260250 60696
rect 261496 57934 261524 84759
rect 261588 60110 261616 129746
rect 261668 117360 261720 117366
rect 261668 117302 261720 117308
rect 261576 60104 261628 60110
rect 261576 60046 261628 60052
rect 261484 57928 261536 57934
rect 261484 57870 261536 57876
rect 261496 57458 261524 57870
rect 260840 57452 260892 57458
rect 260840 57394 260892 57400
rect 261484 57452 261536 57458
rect 261484 57394 261536 57400
rect 260104 22908 260156 22914
rect 260104 22850 260156 22856
rect 259552 22840 259604 22846
rect 259552 22782 259604 22788
rect 259564 16574 259592 22782
rect 260852 16574 260880 57394
rect 261680 57254 261708 117302
rect 261772 114510 261800 154566
rect 262232 144838 262260 202302
rect 262312 198212 262364 198218
rect 262312 198154 262364 198160
rect 262324 171018 262352 198154
rect 262404 182844 262456 182850
rect 262404 182786 262456 182792
rect 262416 173874 262444 182786
rect 262876 181558 262904 229774
rect 262956 227792 263008 227798
rect 262956 227734 263008 227740
rect 262968 204950 262996 227734
rect 263600 218816 263652 218822
rect 263600 218758 263652 218764
rect 262956 204944 263008 204950
rect 262956 204886 263008 204892
rect 262864 181552 262916 181558
rect 262864 181494 262916 181500
rect 263048 173936 263100 173942
rect 263048 173878 263100 173884
rect 262404 173868 262456 173874
rect 262404 173810 262456 173816
rect 262312 171012 262364 171018
rect 262312 170954 262364 170960
rect 262864 161492 262916 161498
rect 262864 161434 262916 161440
rect 262220 144832 262272 144838
rect 262220 144774 262272 144780
rect 262876 122670 262904 161434
rect 262956 139528 263008 139534
rect 262956 139470 263008 139476
rect 262864 122664 262916 122670
rect 262864 122606 262916 122612
rect 261760 114504 261812 114510
rect 261760 114446 261812 114452
rect 262864 99408 262916 99414
rect 262864 99350 262916 99356
rect 262220 71800 262272 71806
rect 262220 71742 262272 71748
rect 261668 57248 261720 57254
rect 261668 57190 261720 57196
rect 262232 16574 262260 71742
rect 259564 16546 260696 16574
rect 260852 16546 261800 16574
rect 262232 16546 262536 16574
rect 260668 480 260696 16546
rect 261772 480 261800 16546
rect 248758 354 248870 480
rect 248432 326 248870 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 16546
rect 262876 14550 262904 99350
rect 262968 98666 262996 139470
rect 263060 136474 263088 173878
rect 263612 171086 263640 218758
rect 264980 192636 265032 192642
rect 264980 192578 265032 192584
rect 263784 183184 263836 183190
rect 263784 183126 263836 183132
rect 263692 181824 263744 181830
rect 263692 181766 263744 181772
rect 263600 171080 263652 171086
rect 263600 171022 263652 171028
rect 263704 161430 263732 181766
rect 263796 164150 263824 183126
rect 264428 167068 264480 167074
rect 264428 167010 264480 167016
rect 264336 166320 264388 166326
rect 264336 166262 264388 166268
rect 263784 164144 263836 164150
rect 263784 164086 263836 164092
rect 263692 161424 263744 161430
rect 263692 161366 263744 161372
rect 264244 139596 264296 139602
rect 264244 139538 264296 139544
rect 263048 136468 263100 136474
rect 263048 136410 263100 136416
rect 263048 119468 263100 119474
rect 263048 119410 263100 119416
rect 263060 100570 263088 119410
rect 263048 100564 263100 100570
rect 263048 100506 263100 100512
rect 262956 98660 263008 98666
rect 262956 98602 263008 98608
rect 262956 93152 263008 93158
rect 262956 93094 263008 93100
rect 262968 73098 262996 93094
rect 262956 73092 263008 73098
rect 262956 73034 263008 73040
rect 262968 71806 262996 73034
rect 262956 71800 263008 71806
rect 262956 71742 263008 71748
rect 264256 24138 264284 139538
rect 264348 132326 264376 166262
rect 264336 132320 264388 132326
rect 264336 132262 264388 132268
rect 264440 129606 264468 167010
rect 264992 162790 265020 192578
rect 265636 188358 265664 232999
rect 266372 219434 266400 239770
rect 268384 235272 268436 235278
rect 268384 235214 268436 235220
rect 266360 219428 266412 219434
rect 266360 219370 266412 219376
rect 266372 218074 266400 219370
rect 266360 218068 266412 218074
rect 266360 218010 266412 218016
rect 267004 218068 267056 218074
rect 267004 218010 267056 218016
rect 266360 203788 266412 203794
rect 266360 203730 266412 203736
rect 265624 188352 265676 188358
rect 265624 188294 265676 188300
rect 265072 183116 265124 183122
rect 265072 183058 265124 183064
rect 264980 162784 265032 162790
rect 264980 162726 265032 162732
rect 264520 158840 264572 158846
rect 264520 158782 264572 158788
rect 264428 129600 264480 129606
rect 264428 129542 264480 129548
rect 264336 128376 264388 128382
rect 264336 128318 264388 128324
rect 264348 53174 264376 128318
rect 264532 123486 264560 158782
rect 265084 155922 265112 183058
rect 265808 174004 265860 174010
rect 265808 173946 265860 173952
rect 265716 171148 265768 171154
rect 265716 171090 265768 171096
rect 265072 155916 265124 155922
rect 265072 155858 265124 155864
rect 265624 147756 265676 147762
rect 265624 147698 265676 147704
rect 264520 123480 264572 123486
rect 264520 123422 264572 123428
rect 265636 107642 265664 147698
rect 265728 133754 265756 171090
rect 265820 141506 265848 173946
rect 266372 143546 266400 203730
rect 266544 184476 266596 184482
rect 266544 184418 266596 184424
rect 266452 180328 266504 180334
rect 266452 180270 266504 180276
rect 266360 143540 266412 143546
rect 266360 143482 266412 143488
rect 266464 143478 266492 180270
rect 266556 162858 266584 184418
rect 267016 176050 267044 218010
rect 267740 195288 267792 195294
rect 267740 195230 267792 195236
rect 267004 176044 267056 176050
rect 267004 175986 267056 175992
rect 267188 169856 267240 169862
rect 267188 169798 267240 169804
rect 266544 162852 266596 162858
rect 266544 162794 266596 162800
rect 267004 156052 267056 156058
rect 267004 155994 267056 156000
rect 266452 143472 266504 143478
rect 266452 143414 266504 143420
rect 265808 141500 265860 141506
rect 265808 141442 265860 141448
rect 265808 134564 265860 134570
rect 265808 134506 265860 134512
rect 265716 133748 265768 133754
rect 265716 133690 265768 133696
rect 265716 113280 265768 113286
rect 265716 113222 265768 113228
rect 265624 107636 265676 107642
rect 265624 107578 265676 107584
rect 265624 104984 265676 104990
rect 265624 104926 265676 104932
rect 264428 100768 264480 100774
rect 264428 100710 264480 100716
rect 264336 53168 264388 53174
rect 264336 53110 264388 53116
rect 264440 37942 264468 100710
rect 264520 98116 264572 98122
rect 264520 98058 264572 98064
rect 264532 58682 264560 98058
rect 264980 58880 265032 58886
rect 264980 58822 265032 58828
rect 264992 58682 265020 58822
rect 264520 58676 264572 58682
rect 264520 58618 264572 58624
rect 264980 58676 265032 58682
rect 264980 58618 265032 58624
rect 264428 37936 264480 37942
rect 264428 37878 264480 37884
rect 264336 35216 264388 35222
rect 264336 35158 264388 35164
rect 264348 24818 264376 35158
rect 264336 24812 264388 24818
rect 264336 24754 264388 24760
rect 264244 24132 264296 24138
rect 264244 24074 264296 24080
rect 264348 23526 264376 24754
rect 263600 23520 263652 23526
rect 263600 23462 263652 23468
rect 264336 23520 264388 23526
rect 264336 23462 264388 23468
rect 263612 16574 263640 23462
rect 263612 16546 264192 16574
rect 262864 14544 262916 14550
rect 262864 14486 262916 14492
rect 264164 480 264192 16546
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 264992 354 265020 58618
rect 265636 18698 265664 104926
rect 265728 26926 265756 113222
rect 265820 106214 265848 134506
rect 267016 117230 267044 155994
rect 267096 140820 267148 140826
rect 267096 140762 267148 140768
rect 267004 117224 267056 117230
rect 267004 117166 267056 117172
rect 267004 111852 267056 111858
rect 267004 111794 267056 111800
rect 265808 106208 265860 106214
rect 265808 106150 265860 106156
rect 266360 84924 266412 84930
rect 266360 84866 266412 84872
rect 266372 78674 266400 84866
rect 266360 78668 266412 78674
rect 266360 78610 266412 78616
rect 265716 26920 265768 26926
rect 265716 26862 265768 26868
rect 265624 18692 265676 18698
rect 265624 18634 265676 18640
rect 266372 16574 266400 78610
rect 266372 16546 266584 16574
rect 266556 480 266584 16546
rect 267016 7614 267044 111794
rect 267108 101454 267136 140762
rect 267200 131102 267228 169798
rect 267752 146266 267780 195230
rect 267832 189848 267884 189854
rect 267832 189790 267884 189796
rect 267844 156670 267872 189790
rect 268396 189106 268424 235214
rect 269132 231810 269160 239788
rect 269120 231804 269172 231810
rect 269120 231746 269172 231752
rect 269764 231804 269816 231810
rect 269764 231746 269816 231752
rect 269776 200938 269804 231746
rect 271892 215286 271920 239788
rect 271880 215280 271932 215286
rect 271880 215222 271932 215228
rect 271892 214810 271920 215222
rect 271880 214804 271932 214810
rect 271880 214746 271932 214752
rect 272524 214804 272576 214810
rect 272524 214746 272576 214752
rect 270500 214668 270552 214674
rect 270500 214610 270552 214616
rect 269764 200932 269816 200938
rect 269764 200874 269816 200880
rect 269120 191208 269172 191214
rect 269120 191150 269172 191156
rect 268384 189100 268436 189106
rect 268384 189042 268436 189048
rect 267924 178832 267976 178838
rect 267924 178774 267976 178780
rect 267832 156664 267884 156670
rect 267832 156606 267884 156612
rect 267936 153066 267964 178774
rect 268384 167136 268436 167142
rect 268384 167078 268436 167084
rect 267924 153060 267976 153066
rect 267924 153002 267976 153008
rect 267740 146260 267792 146266
rect 267740 146202 267792 146208
rect 267188 131096 267240 131102
rect 267188 131038 267240 131044
rect 268396 128246 268424 167078
rect 268476 151904 268528 151910
rect 268476 151846 268528 151852
rect 268384 128240 268436 128246
rect 268384 128182 268436 128188
rect 268384 120216 268436 120222
rect 268384 120158 268436 120164
rect 267188 103556 267240 103562
rect 267188 103498 267240 103504
rect 267096 101448 267148 101454
rect 267096 101390 267148 101396
rect 267200 75206 267228 103498
rect 267188 75200 267240 75206
rect 267188 75142 267240 75148
rect 268396 58818 268424 120158
rect 268488 113830 268516 151846
rect 269132 144906 269160 191150
rect 269212 189100 269264 189106
rect 269212 189042 269264 189048
rect 269224 153134 269252 189042
rect 269856 164280 269908 164286
rect 269856 164222 269908 164228
rect 269212 153128 269264 153134
rect 269212 153070 269264 153076
rect 269120 144900 269172 144906
rect 269120 144842 269172 144848
rect 269764 142248 269816 142254
rect 269764 142190 269816 142196
rect 268568 127696 268620 127702
rect 268568 127638 268620 127644
rect 268476 113824 268528 113830
rect 268476 113766 268528 113772
rect 268580 100638 268608 127638
rect 269776 102134 269804 142190
rect 269868 125526 269896 164222
rect 270512 164218 270540 214610
rect 271972 196852 272024 196858
rect 271972 196794 272024 196800
rect 271878 195256 271934 195265
rect 271878 195191 271934 195200
rect 270684 188556 270736 188562
rect 270684 188498 270736 188504
rect 270592 187060 270644 187066
rect 270592 187002 270644 187008
rect 270500 164212 270552 164218
rect 270500 164154 270552 164160
rect 269948 161560 270000 161566
rect 269948 161502 270000 161508
rect 269856 125520 269908 125526
rect 269856 125462 269908 125468
rect 269960 122738 269988 161502
rect 270604 147626 270632 187002
rect 270696 157350 270724 188498
rect 271144 165640 271196 165646
rect 271144 165582 271196 165588
rect 270684 157344 270736 157350
rect 270684 157286 270736 157292
rect 270592 147620 270644 147626
rect 270592 147562 270644 147568
rect 271156 128314 271184 165582
rect 271236 154692 271288 154698
rect 271236 154634 271288 154640
rect 271144 128308 271196 128314
rect 271144 128250 271196 128256
rect 269948 122732 270000 122738
rect 269948 122674 270000 122680
rect 269856 121508 269908 121514
rect 269856 121450 269908 121456
rect 269764 102128 269816 102134
rect 269764 102070 269816 102076
rect 268568 100632 268620 100638
rect 268568 100574 268620 100580
rect 269764 96756 269816 96762
rect 269764 96698 269816 96704
rect 268476 60104 268528 60110
rect 268476 60046 268528 60052
rect 268384 58812 268436 58818
rect 268384 58754 268436 58760
rect 268488 20641 268516 60046
rect 269120 49632 269172 49638
rect 269120 49574 269172 49580
rect 267738 20632 267794 20641
rect 267738 20567 267794 20576
rect 268474 20632 268530 20641
rect 268474 20567 268530 20576
rect 267752 16574 267780 20567
rect 269132 16574 269160 49574
rect 269776 36582 269804 96698
rect 269868 73914 269896 121450
rect 271248 115870 271276 154634
rect 271892 136542 271920 195191
rect 271984 153202 272012 196794
rect 272536 192642 272564 214746
rect 273272 213926 273300 239788
rect 276032 237114 276060 240040
rect 277918 239850 277946 240040
rect 280494 239850 280522 240040
rect 282426 239850 282454 240040
rect 277412 239822 277946 239850
rect 280172 239822 280522 239850
rect 281552 239822 282454 239850
rect 276020 237108 276072 237114
rect 276020 237050 276072 237056
rect 276032 236026 276060 237050
rect 276020 236020 276072 236026
rect 276020 235962 276072 235968
rect 276664 236020 276716 236026
rect 276664 235962 276716 235968
rect 276676 224262 276704 235962
rect 277412 231606 277440 239822
rect 277400 231600 277452 231606
rect 277400 231542 277452 231548
rect 278044 231600 278096 231606
rect 278044 231542 278096 231548
rect 276664 224256 276716 224262
rect 276664 224198 276716 224204
rect 273260 213920 273312 213926
rect 273260 213862 273312 213868
rect 273904 213920 273956 213926
rect 273904 213862 273956 213868
rect 272524 192636 272576 192642
rect 272524 192578 272576 192584
rect 273444 191140 273496 191146
rect 273444 191082 273496 191088
rect 273352 185632 273404 185638
rect 273352 185574 273404 185580
rect 273260 184408 273312 184414
rect 273260 184350 273312 184356
rect 272064 180464 272116 180470
rect 272064 180406 272116 180412
rect 271972 153196 272024 153202
rect 271972 153138 272024 153144
rect 272076 149054 272104 180406
rect 272524 163600 272576 163606
rect 272524 163542 272576 163548
rect 272064 149048 272116 149054
rect 272064 148990 272116 148996
rect 271880 136536 271932 136542
rect 271880 136478 271932 136484
rect 272536 126954 272564 163542
rect 272616 146396 272668 146402
rect 272616 146338 272668 146344
rect 272524 126948 272576 126954
rect 272524 126890 272576 126896
rect 272524 124228 272576 124234
rect 272524 124170 272576 124176
rect 271236 115864 271288 115870
rect 271236 115806 271288 115812
rect 271144 114572 271196 114578
rect 271144 114514 271196 114520
rect 269948 100836 270000 100842
rect 269948 100778 270000 100784
rect 269856 73908 269908 73914
rect 269856 73850 269908 73856
rect 269856 65612 269908 65618
rect 269856 65554 269908 65560
rect 269868 49638 269896 65554
rect 269960 62830 269988 100778
rect 269948 62824 270000 62830
rect 269948 62766 270000 62772
rect 269856 49632 269908 49638
rect 269856 49574 269908 49580
rect 271156 49026 271184 114514
rect 271878 61568 271934 61577
rect 271878 61503 271934 61512
rect 271144 49020 271196 49026
rect 271144 48962 271196 48968
rect 269764 36576 269816 36582
rect 269764 36518 269816 36524
rect 270500 26920 270552 26926
rect 270500 26862 270552 26868
rect 270512 16574 270540 26862
rect 267752 16546 268424 16574
rect 269132 16546 270080 16574
rect 270512 16546 270816 16574
rect 267004 7608 267056 7614
rect 267004 7550 267056 7556
rect 267740 3596 267792 3602
rect 267740 3538 267792 3544
rect 267752 480 267780 3538
rect 265318 354 265430 480
rect 264992 326 265430 354
rect 265318 -960 265430 326
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 354 268424 16546
rect 270052 480 270080 16546
rect 268814 354 268926 480
rect 268396 326 268926 354
rect 268814 -960 268926 326
rect 270010 -960 270122 480
rect 270788 354 270816 16546
rect 271892 3482 271920 61503
rect 272536 61470 272564 124170
rect 272628 104786 272656 146338
rect 273272 140758 273300 184350
rect 273364 148345 273392 185574
rect 273456 160070 273484 191082
rect 273916 180334 273944 213862
rect 274640 211880 274692 211886
rect 274640 211822 274692 211828
rect 273904 180328 273956 180334
rect 273904 180270 273956 180276
rect 273444 160064 273496 160070
rect 273444 160006 273496 160012
rect 273904 158908 273956 158914
rect 273904 158850 273956 158856
rect 273350 148336 273406 148345
rect 273350 148271 273406 148280
rect 273260 140752 273312 140758
rect 273260 140694 273312 140700
rect 273916 120086 273944 158850
rect 274652 137970 274680 211822
rect 274732 200864 274784 200870
rect 274732 200806 274784 200812
rect 274744 154562 274772 200806
rect 276664 199640 276716 199646
rect 276664 199582 276716 199588
rect 274732 154556 274784 154562
rect 274732 154498 274784 154504
rect 275376 153400 275428 153406
rect 275376 153342 275428 153348
rect 274640 137964 274692 137970
rect 274640 137906 274692 137912
rect 275284 125656 275336 125662
rect 275284 125598 275336 125604
rect 273904 120080 273956 120086
rect 273904 120022 273956 120028
rect 273904 116068 273956 116074
rect 273904 116010 273956 116016
rect 272616 104780 272668 104786
rect 272616 104722 272668 104728
rect 272616 99476 272668 99482
rect 272616 99418 272668 99424
rect 272524 61464 272576 61470
rect 272524 61406 272576 61412
rect 272628 39370 272656 99418
rect 273166 61568 273222 61577
rect 273166 61503 273222 61512
rect 273180 61402 273208 61503
rect 273168 61396 273220 61402
rect 273168 61338 273220 61344
rect 273260 47388 273312 47394
rect 273260 47330 273312 47336
rect 272616 39364 272668 39370
rect 272616 39306 272668 39312
rect 271972 25628 272024 25634
rect 271972 25570 272024 25576
rect 271984 3602 272012 25570
rect 271972 3596 272024 3602
rect 271972 3538 272024 3544
rect 271892 3454 272472 3482
rect 272444 480 272472 3454
rect 271206 354 271318 480
rect 270788 326 271318 354
rect 271206 -960 271318 326
rect 272402 -960 272514 480
rect 273272 354 273300 47330
rect 273916 33862 273944 116010
rect 273996 110560 274048 110566
rect 273996 110502 274048 110508
rect 274008 47598 274036 110502
rect 274088 64252 274140 64258
rect 274088 64194 274140 64200
rect 274100 48278 274128 64194
rect 274088 48272 274140 48278
rect 274088 48214 274140 48220
rect 273996 47592 274048 47598
rect 273996 47534 274048 47540
rect 274100 47394 274128 48214
rect 274088 47388 274140 47394
rect 274088 47330 274140 47336
rect 273904 33856 273956 33862
rect 273904 33798 273956 33804
rect 274640 28348 274692 28354
rect 274640 28290 274692 28296
rect 274652 16574 274680 28290
rect 275296 22778 275324 125598
rect 275388 117978 275416 153342
rect 275376 117972 275428 117978
rect 275376 117914 275428 117920
rect 275376 103624 275428 103630
rect 275376 103566 275428 103572
rect 275388 54670 275416 103566
rect 276018 76664 276074 76673
rect 276018 76599 276074 76608
rect 275376 54664 275428 54670
rect 275376 54606 275428 54612
rect 275284 22772 275336 22778
rect 275284 22714 275336 22720
rect 274652 16546 274864 16574
rect 274836 480 274864 16546
rect 276032 6914 276060 76599
rect 276676 64258 276704 199582
rect 278056 185638 278084 231542
rect 280172 230450 280200 239822
rect 280160 230444 280212 230450
rect 280160 230386 280212 230392
rect 281448 230444 281500 230450
rect 281448 230386 281500 230392
rect 281460 229770 281488 230386
rect 281448 229764 281500 229770
rect 281448 229706 281500 229712
rect 278780 218748 278832 218754
rect 278780 218690 278832 218696
rect 278044 185632 278096 185638
rect 278044 185574 278096 185580
rect 278044 184340 278096 184346
rect 278044 184282 278096 184288
rect 276756 172576 276808 172582
rect 276756 172518 276808 172524
rect 276768 135182 276796 172518
rect 277032 145580 277084 145586
rect 277032 145522 277084 145528
rect 276940 144220 276992 144226
rect 276940 144162 276992 144168
rect 276756 135176 276808 135182
rect 276756 135118 276808 135124
rect 276848 116136 276900 116142
rect 276848 116078 276900 116084
rect 276756 103692 276808 103698
rect 276756 103634 276808 103640
rect 276664 64252 276716 64258
rect 276664 64194 276716 64200
rect 276662 29608 276718 29617
rect 276662 29543 276718 29552
rect 276676 11778 276704 29543
rect 276768 13122 276796 103634
rect 276860 28286 276888 116078
rect 276952 104854 276980 144162
rect 277044 117298 277072 145522
rect 277032 117292 277084 117298
rect 277032 117234 277084 117240
rect 276940 104848 276992 104854
rect 276940 104790 276992 104796
rect 278056 93838 278084 184282
rect 278228 171216 278280 171222
rect 278228 171158 278280 171164
rect 278240 132394 278268 171158
rect 278792 150414 278820 218690
rect 281552 209778 281580 239822
rect 284404 237454 284432 240040
rect 286934 239834 286962 240040
rect 285680 239828 285732 239834
rect 285680 239770 285732 239776
rect 286922 239828 286974 239834
rect 286922 239770 286974 239776
rect 283564 237448 283616 237454
rect 283564 237390 283616 237396
rect 284392 237448 284444 237454
rect 284392 237390 284444 237396
rect 283576 218006 283604 237390
rect 283564 218000 283616 218006
rect 283564 217942 283616 217948
rect 281540 209772 281592 209778
rect 281540 209714 281592 209720
rect 281552 208418 281580 209714
rect 281540 208412 281592 208418
rect 281540 208354 281592 208360
rect 282276 208412 282328 208418
rect 282276 208354 282328 208360
rect 282184 206372 282236 206378
rect 282184 206314 282236 206320
rect 280804 203720 280856 203726
rect 280804 203662 280856 203668
rect 280160 202224 280212 202230
rect 280160 202166 280212 202172
rect 279422 181520 279478 181529
rect 279422 181455 279478 181464
rect 278780 150408 278832 150414
rect 278780 150350 278832 150356
rect 278228 132388 278280 132394
rect 278228 132330 278280 132336
rect 278136 131164 278188 131170
rect 278136 131106 278188 131112
rect 278044 93832 278096 93838
rect 278044 93774 278096 93780
rect 278044 62824 278096 62830
rect 278044 62766 278096 62772
rect 277400 30320 277452 30326
rect 277400 30262 277452 30268
rect 276848 28280 276900 28286
rect 276848 28222 276900 28228
rect 277412 16574 277440 30262
rect 278056 29617 278084 62766
rect 278148 60042 278176 131106
rect 279436 122126 279464 181455
rect 279516 150612 279568 150618
rect 279516 150554 279568 150560
rect 279424 122120 279476 122126
rect 279424 122062 279476 122068
rect 278320 118856 278372 118862
rect 278320 118798 278372 118804
rect 278228 77988 278280 77994
rect 278228 77930 278280 77936
rect 278136 60036 278188 60042
rect 278136 59978 278188 59984
rect 278240 30326 278268 77930
rect 278332 71058 278360 118798
rect 279528 110294 279556 150554
rect 280172 139398 280200 202166
rect 280160 139392 280212 139398
rect 280160 139334 280212 139340
rect 279516 110288 279568 110294
rect 279516 110230 279568 110236
rect 279424 107772 279476 107778
rect 279424 107714 279476 107720
rect 278320 71052 278372 71058
rect 278320 70994 278372 71000
rect 278780 64252 278832 64258
rect 278780 64194 278832 64200
rect 278228 30320 278280 30326
rect 278228 30262 278280 30268
rect 278042 29608 278098 29617
rect 278042 29543 278098 29552
rect 278792 16574 278820 64194
rect 279436 29646 279464 107714
rect 280816 89078 280844 203662
rect 281080 156120 281132 156126
rect 281080 156062 281132 156068
rect 280988 135380 281040 135386
rect 280988 135322 281040 135328
rect 280896 114640 280948 114646
rect 280896 114582 280948 114588
rect 280804 89072 280856 89078
rect 280804 89014 280856 89020
rect 280802 62792 280858 62801
rect 280802 62727 280858 62736
rect 279424 29640 279476 29646
rect 279424 29582 279476 29588
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 276756 13116 276808 13122
rect 276756 13058 276808 13064
rect 276676 11750 276796 11778
rect 276032 6886 276704 6914
rect 276020 3460 276072 3466
rect 276020 3402 276072 3408
rect 276032 480 276060 3402
rect 273598 354 273710 480
rect 273272 326 273710 354
rect 273598 -960 273710 326
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 354 276704 6886
rect 276768 3466 276796 11750
rect 276756 3460 276808 3466
rect 276756 3402 276808 3408
rect 278332 480 278360 16546
rect 277094 354 277206 480
rect 276676 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279068 354 279096 16546
rect 280816 8226 280844 62727
rect 280908 11762 280936 114582
rect 281000 32434 281028 135322
rect 281092 115938 281120 156062
rect 281080 115932 281132 115938
rect 281080 115874 281132 115880
rect 280988 32428 281040 32434
rect 280988 32370 281040 32376
rect 282196 16574 282224 206314
rect 282288 96626 282316 208354
rect 283576 177546 283604 217942
rect 285692 205630 285720 239770
rect 288912 234666 288940 240040
rect 290798 239816 290826 240040
rect 289832 239788 290826 239816
rect 292796 239816 292824 240040
rect 292796 239788 293264 239816
rect 288900 234660 288952 234666
rect 288900 234602 288952 234608
rect 289452 234660 289504 234666
rect 289452 234602 289504 234608
rect 289464 233209 289492 234602
rect 289450 233200 289506 233209
rect 289450 233135 289506 233144
rect 289832 226234 289860 239788
rect 293236 234569 293264 239788
rect 293222 234560 293278 234569
rect 293222 234495 293278 234504
rect 289820 226228 289872 226234
rect 289820 226170 289872 226176
rect 289832 225010 289860 226170
rect 289820 225004 289872 225010
rect 289820 224946 289872 224952
rect 290464 225004 290516 225010
rect 290464 224946 290516 224952
rect 289084 220176 289136 220182
rect 289084 220118 289136 220124
rect 287702 211984 287758 211993
rect 287702 211919 287758 211928
rect 285680 205624 285732 205630
rect 285680 205566 285732 205572
rect 285692 205154 285720 205566
rect 285680 205148 285732 205154
rect 285680 205090 285732 205096
rect 286416 205148 286468 205154
rect 286416 205090 286468 205096
rect 286324 193996 286376 194002
rect 286324 193938 286376 193944
rect 283564 177540 283616 177546
rect 283564 177482 283616 177488
rect 284944 174072 284996 174078
rect 284944 174014 284996 174020
rect 283564 157480 283616 157486
rect 283564 157422 283616 157428
rect 283576 151162 283604 157422
rect 283564 151156 283616 151162
rect 283564 151098 283616 151104
rect 283656 149184 283708 149190
rect 283656 149126 283708 149132
rect 283564 125724 283616 125730
rect 283564 125666 283616 125672
rect 282368 117428 282420 117434
rect 282368 117370 282420 117376
rect 282276 96620 282328 96626
rect 282276 96562 282328 96568
rect 281920 16546 282224 16574
rect 280896 11756 280948 11762
rect 280896 11698 280948 11704
rect 280804 8220 280856 8226
rect 280804 8162 280856 8168
rect 280816 6914 280844 8162
rect 280724 6886 280844 6914
rect 280724 480 280752 6886
rect 281920 6866 281948 16546
rect 282276 16040 282328 16046
rect 282276 15982 282328 15988
rect 281908 6860 281960 6866
rect 281908 6802 281960 6808
rect 281920 480 281948 6802
rect 282288 4078 282316 15982
rect 282380 10402 282408 117370
rect 283576 17270 283604 125666
rect 283668 109002 283696 149126
rect 284956 136610 284984 174014
rect 285128 146464 285180 146470
rect 285128 146406 285180 146412
rect 284944 136604 284996 136610
rect 284944 136546 284996 136552
rect 284944 128444 284996 128450
rect 284944 128386 284996 128392
rect 283656 108996 283708 109002
rect 283656 108938 283708 108944
rect 283656 105052 283708 105058
rect 283656 104994 283708 105000
rect 283564 17264 283616 17270
rect 283564 17206 283616 17212
rect 283564 11756 283616 11762
rect 283564 11698 283616 11704
rect 282368 10396 282420 10402
rect 282368 10338 282420 10344
rect 283576 8294 283604 11698
rect 283668 9042 283696 104994
rect 284298 46880 284354 46889
rect 284298 46815 284354 46824
rect 283656 9036 283708 9042
rect 283656 8978 283708 8984
rect 283564 8288 283616 8294
rect 283564 8230 283616 8236
rect 282276 4072 282328 4078
rect 282276 4014 282328 4020
rect 279486 354 279598 480
rect 279068 326 279598 354
rect 279486 -960 279598 326
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 354 283186 480
rect 283576 354 283604 8230
rect 284312 480 284340 46815
rect 284392 31272 284444 31278
rect 284392 31214 284444 31220
rect 284404 6914 284432 31214
rect 284956 14618 284984 128386
rect 285036 124296 285088 124302
rect 285036 124238 285088 124244
rect 285048 46374 285076 124238
rect 285140 106282 285168 146406
rect 285128 106276 285180 106282
rect 285128 106218 285180 106224
rect 285128 100904 285180 100910
rect 285128 100846 285180 100852
rect 285036 46368 285088 46374
rect 285036 46310 285088 46316
rect 285140 42090 285168 100846
rect 286336 68338 286364 193938
rect 286428 193934 286456 205090
rect 286416 193928 286468 193934
rect 286416 193870 286468 193876
rect 286508 140888 286560 140894
rect 286508 140830 286560 140836
rect 286416 133952 286468 133958
rect 286416 133894 286468 133900
rect 286324 68332 286376 68338
rect 286324 68274 286376 68280
rect 285680 66224 285732 66230
rect 285680 66166 285732 66172
rect 285218 61432 285274 61441
rect 285218 61367 285274 61376
rect 285232 46889 285260 61367
rect 285218 46880 285274 46889
rect 285218 46815 285274 46824
rect 285128 42084 285180 42090
rect 285128 42026 285180 42032
rect 284944 14612 284996 14618
rect 284944 14554 284996 14560
rect 285692 6914 285720 66166
rect 286428 15978 286456 133894
rect 286520 100706 286548 140830
rect 286508 100700 286560 100706
rect 286508 100642 286560 100648
rect 286508 78056 286560 78062
rect 286508 77998 286560 78004
rect 286520 66230 286548 77998
rect 287716 67590 287744 211919
rect 287980 160268 288032 160274
rect 287980 160210 288032 160216
rect 287796 138168 287848 138174
rect 287796 138110 287848 138116
rect 287704 67584 287756 67590
rect 287704 67526 287756 67532
rect 286508 66224 286560 66230
rect 286508 66166 286560 66172
rect 287808 39438 287836 138110
rect 287992 121446 288020 160210
rect 287980 121440 288032 121446
rect 287980 121382 288032 121388
rect 287888 120284 287940 120290
rect 287888 120226 287940 120232
rect 287900 71126 287928 120226
rect 289096 94518 289124 220118
rect 290476 195294 290504 224946
rect 293236 220114 293264 234495
rect 293224 220108 293276 220114
rect 293224 220050 293276 220056
rect 295352 216646 295380 240040
rect 297238 239850 297266 240040
rect 296732 239822 297266 239850
rect 296732 224874 296760 239822
rect 299216 238678 299244 240040
rect 301746 239850 301774 240040
rect 301516 239822 301774 239850
rect 299204 238672 299256 238678
rect 299204 238614 299256 238620
rect 299216 231849 299244 238614
rect 301516 235754 301544 239822
rect 303724 237182 303752 240040
rect 304264 238876 304316 238882
rect 304264 238818 304316 238824
rect 304276 238610 304304 238818
rect 305656 238649 305684 240040
rect 308186 239850 308214 240040
rect 310118 239850 310146 240040
rect 307772 239822 308214 239850
rect 309152 239822 310146 239850
rect 305642 238640 305698 238649
rect 304264 238604 304316 238610
rect 305642 238575 305698 238584
rect 304264 238546 304316 238552
rect 303712 237176 303764 237182
rect 303712 237118 303764 237124
rect 303724 236026 303752 237118
rect 303712 236020 303764 236026
rect 303712 235962 303764 235968
rect 304264 236020 304316 236026
rect 304264 235962 304316 235968
rect 301504 235748 301556 235754
rect 301504 235690 301556 235696
rect 299202 231840 299258 231849
rect 299202 231775 299258 231784
rect 296720 224868 296772 224874
rect 296720 224810 296772 224816
rect 297364 224868 297416 224874
rect 297364 224810 297416 224816
rect 295340 216640 295392 216646
rect 295340 216582 295392 216588
rect 295352 215354 295380 216582
rect 295340 215348 295392 215354
rect 295340 215290 295392 215296
rect 295984 215348 296036 215354
rect 295984 215290 296036 215296
rect 291844 213444 291896 213450
rect 291844 213386 291896 213392
rect 290464 195288 290516 195294
rect 290464 195230 290516 195236
rect 289268 147824 289320 147830
rect 289268 147766 289320 147772
rect 289176 135448 289228 135454
rect 289176 135390 289228 135396
rect 289084 94512 289136 94518
rect 289084 94454 289136 94460
rect 289082 75168 289138 75177
rect 289082 75103 289138 75112
rect 287888 71120 287940 71126
rect 287888 71062 287940 71068
rect 288348 39636 288400 39642
rect 288348 39578 288400 39584
rect 287796 39432 287848 39438
rect 287796 39374 287848 39380
rect 288360 37262 288388 39578
rect 287060 37256 287112 37262
rect 287060 37198 287112 37204
rect 288348 37256 288400 37262
rect 288348 37198 288400 37204
rect 287072 16574 287100 37198
rect 289096 34474 289124 75103
rect 289188 49094 289216 135390
rect 289280 112538 289308 147766
rect 290464 137284 290516 137290
rect 290464 137226 290516 137232
rect 290476 118658 290504 137226
rect 290556 131232 290608 131238
rect 290556 131174 290608 131180
rect 290464 118652 290516 118658
rect 290464 118594 290516 118600
rect 290464 114708 290516 114714
rect 290464 114650 290516 114656
rect 289268 112532 289320 112538
rect 289268 112474 289320 112480
rect 289268 109064 289320 109070
rect 289268 109006 289320 109012
rect 289176 49088 289228 49094
rect 289176 49030 289228 49036
rect 289084 34468 289136 34474
rect 289084 34410 289136 34416
rect 289096 33182 289124 34410
rect 288440 33176 288492 33182
rect 288440 33118 288492 33124
rect 289084 33176 289136 33182
rect 289084 33118 289136 33124
rect 288452 16574 288480 33118
rect 289280 31142 289308 109006
rect 289820 67584 289872 67590
rect 289820 67526 289872 67532
rect 289832 66978 289860 67526
rect 289820 66972 289872 66978
rect 289820 66914 289872 66920
rect 289268 31136 289320 31142
rect 289268 31078 289320 31084
rect 287072 16546 287376 16574
rect 288452 16546 289032 16574
rect 286416 15972 286468 15978
rect 286416 15914 286468 15920
rect 284404 6886 284984 6914
rect 285692 6886 286640 6914
rect 283074 326 283604 354
rect 283074 -960 283186 326
rect 284270 -960 284382 480
rect 284956 354 284984 6886
rect 286612 480 286640 6886
rect 285374 354 285486 480
rect 284956 326 285486 354
rect 285374 -960 285486 326
rect 286570 -960 286682 480
rect 287348 354 287376 16546
rect 289004 480 289032 16546
rect 287766 354 287878 480
rect 287348 326 287878 354
rect 287766 -960 287878 326
rect 288962 -960 289074 480
rect 289832 354 289860 66914
rect 290476 33794 290504 114650
rect 290568 72486 290596 131174
rect 291856 84182 291884 213386
rect 295996 178838 296024 215290
rect 297376 189854 297404 224810
rect 301516 222970 301544 235690
rect 301504 222964 301556 222970
rect 301504 222906 301556 222912
rect 304276 210526 304304 235962
rect 305656 227050 305684 238575
rect 307024 233300 307076 233306
rect 307024 233242 307076 233248
rect 305644 227044 305696 227050
rect 305644 226986 305696 226992
rect 304264 210520 304316 210526
rect 304264 210462 304316 210468
rect 297364 189848 297416 189854
rect 297364 189790 297416 189796
rect 307036 181762 307064 233242
rect 307772 211818 307800 239822
rect 309152 222154 309180 239822
rect 312096 238610 312124 240040
rect 313982 239850 314010 240040
rect 313292 239822 314010 239850
rect 312084 238604 312136 238610
rect 312084 238546 312136 238552
rect 312096 237454 312124 238546
rect 312084 237448 312136 237454
rect 312084 237390 312136 237396
rect 312544 237448 312596 237454
rect 312544 237390 312596 237396
rect 309140 222148 309192 222154
rect 309140 222090 309192 222096
rect 309876 222148 309928 222154
rect 309876 222090 309928 222096
rect 307760 211812 307812 211818
rect 307760 211754 307812 211760
rect 307772 211698 307800 211754
rect 307680 211670 307800 211698
rect 307024 181756 307076 181762
rect 307024 181698 307076 181704
rect 295984 178832 296036 178838
rect 295984 178774 296036 178780
rect 294696 177472 294748 177478
rect 294696 177414 294748 177420
rect 291936 167680 291988 167686
rect 291936 167622 291988 167628
rect 291948 129674 291976 167622
rect 293316 162920 293368 162926
rect 293316 162862 293368 162868
rect 292028 132524 292080 132530
rect 292028 132466 292080 132472
rect 291936 129668 291988 129674
rect 291936 129610 291988 129616
rect 291936 113348 291988 113354
rect 291936 113290 291988 113296
rect 291844 84176 291896 84182
rect 291844 84118 291896 84124
rect 291856 82890 291884 84118
rect 291200 82884 291252 82890
rect 291200 82826 291252 82832
rect 291844 82884 291896 82890
rect 291844 82826 291896 82832
rect 290556 72480 290608 72486
rect 290556 72422 290608 72428
rect 290464 33788 290516 33794
rect 290464 33730 290516 33736
rect 291212 16574 291240 82826
rect 291212 16546 291424 16574
rect 291396 480 291424 16546
rect 291948 4826 291976 113290
rect 292040 53242 292068 132466
rect 293224 127016 293276 127022
rect 293224 126958 293276 126964
rect 292580 68332 292632 68338
rect 292580 68274 292632 68280
rect 292028 53236 292080 53242
rect 292028 53178 292080 53184
rect 292592 16574 292620 68274
rect 293236 31074 293264 126958
rect 293328 126274 293356 162862
rect 294604 131300 294656 131306
rect 294604 131242 294656 131248
rect 293316 126268 293368 126274
rect 293316 126210 293368 126216
rect 293316 123004 293368 123010
rect 293316 122946 293368 122952
rect 293328 68406 293356 122946
rect 293316 68400 293368 68406
rect 293316 68342 293368 68348
rect 293960 35352 294012 35358
rect 293960 35294 294012 35300
rect 293972 35222 294000 35294
rect 293960 35216 294012 35222
rect 293960 35158 294012 35164
rect 293224 31068 293276 31074
rect 293224 31010 293276 31016
rect 292592 16546 293264 16574
rect 291936 4820 291988 4826
rect 291936 4762 291988 4768
rect 292580 3052 292632 3058
rect 292580 2994 292632 3000
rect 292592 480 292620 2994
rect 290158 354 290270 480
rect 289832 326 290270 354
rect 290158 -960 290270 326
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293236 354 293264 16546
rect 293972 3058 294000 35158
rect 294616 24206 294644 131242
rect 294708 94994 294736 177414
rect 307680 176118 307708 211670
rect 309784 190120 309836 190126
rect 309784 190062 309836 190068
rect 308404 187332 308456 187338
rect 308404 187274 308456 187280
rect 307668 176112 307720 176118
rect 307668 176054 307720 176060
rect 307390 175264 307446 175273
rect 307390 175199 307446 175208
rect 307298 173632 307354 173641
rect 307298 173567 307354 173576
rect 302884 172712 302936 172718
rect 302884 172654 302936 172660
rect 298744 172644 298796 172650
rect 298744 172586 298796 172592
rect 297456 169924 297508 169930
rect 297456 169866 297508 169872
rect 295984 166388 296036 166394
rect 295984 166330 296036 166336
rect 295996 133822 296024 166330
rect 296076 151972 296128 151978
rect 296076 151914 296128 151920
rect 295984 133816 296036 133822
rect 295984 133758 296036 133764
rect 295984 127084 296036 127090
rect 295984 127026 296036 127032
rect 294788 110628 294840 110634
rect 294788 110570 294840 110576
rect 294696 94988 294748 94994
rect 294696 94930 294748 94936
rect 294800 67046 294828 110570
rect 294788 67040 294840 67046
rect 294788 66982 294840 66988
rect 295340 36644 295392 36650
rect 295340 36586 295392 36592
rect 294604 24200 294656 24206
rect 294604 24142 294656 24148
rect 295352 16574 295380 36586
rect 295352 16546 295656 16574
rect 294880 4888 294932 4894
rect 294880 4830 294932 4836
rect 293960 3052 294012 3058
rect 293960 2994 294012 3000
rect 294892 480 294920 4830
rect 293654 354 293766 480
rect 293236 326 293766 354
rect 293654 -960 293766 326
rect 294850 -960 294962 480
rect 295628 354 295656 16546
rect 295996 6186 296024 127026
rect 296088 111790 296116 151914
rect 297364 132592 297416 132598
rect 297364 132534 297416 132540
rect 296168 125792 296220 125798
rect 296168 125734 296220 125740
rect 296076 111784 296128 111790
rect 296076 111726 296128 111732
rect 296076 99544 296128 99550
rect 296076 99486 296128 99492
rect 296088 25566 296116 99486
rect 296180 56030 296208 125734
rect 296168 56024 296220 56030
rect 296168 55966 296220 55972
rect 297376 54602 297404 132534
rect 297468 132462 297496 169866
rect 298756 133890 298784 172586
rect 300308 168496 300360 168502
rect 300308 168438 300360 168444
rect 299020 161628 299072 161634
rect 299020 161570 299072 161576
rect 298928 150544 298980 150550
rect 298928 150486 298980 150492
rect 298744 133884 298796 133890
rect 298744 133826 298796 133832
rect 297456 132456 297508 132462
rect 297456 132398 297508 132404
rect 298836 128512 298888 128518
rect 298836 128454 298888 128460
rect 298744 121644 298796 121650
rect 298744 121586 298796 121592
rect 297456 121576 297508 121582
rect 297456 121518 297508 121524
rect 297468 75274 297496 121518
rect 297548 102264 297600 102270
rect 297548 102206 297600 102212
rect 297456 75268 297508 75274
rect 297456 75210 297508 75216
rect 297560 65550 297588 102206
rect 297640 75200 297692 75206
rect 297640 75142 297692 75148
rect 297548 65544 297600 65550
rect 297548 65486 297600 65492
rect 297364 54596 297416 54602
rect 297364 54538 297416 54544
rect 297652 45558 297680 75142
rect 296720 45552 296772 45558
rect 296720 45494 296772 45500
rect 297640 45552 297692 45558
rect 297640 45494 297692 45500
rect 296076 25560 296128 25566
rect 296076 25502 296128 25508
rect 296732 16574 296760 45494
rect 298100 28960 298152 28966
rect 298100 28902 298152 28908
rect 296732 16546 297312 16574
rect 295984 6180 296036 6186
rect 295984 6122 296036 6128
rect 297284 480 297312 16546
rect 296046 354 296158 480
rect 295628 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 28902
rect 298756 21486 298784 121586
rect 298848 66910 298876 128454
rect 298940 110362 298968 150486
rect 299032 122806 299060 161570
rect 300124 135516 300176 135522
rect 300124 135458 300176 135464
rect 299020 122800 299072 122806
rect 299020 122742 299072 122748
rect 298928 110356 298980 110362
rect 298928 110298 298980 110304
rect 298928 98184 298980 98190
rect 298928 98126 298980 98132
rect 298836 66904 298888 66910
rect 298836 66846 298888 66852
rect 298940 50386 298968 98126
rect 298928 50380 298980 50386
rect 298928 50322 298980 50328
rect 298836 44872 298888 44878
rect 298836 44814 298888 44820
rect 298848 28966 298876 44814
rect 299480 38072 299532 38078
rect 299480 38014 299532 38020
rect 299492 37942 299520 38014
rect 300136 38010 300164 135458
rect 300216 132660 300268 132666
rect 300216 132602 300268 132608
rect 300228 51814 300256 132602
rect 300320 129742 300348 168438
rect 301596 164348 301648 164354
rect 301596 164290 301648 164296
rect 301504 129940 301556 129946
rect 301504 129882 301556 129888
rect 300308 129736 300360 129742
rect 300308 129678 300360 129684
rect 300308 118720 300360 118726
rect 300308 118662 300360 118668
rect 300320 64190 300348 118662
rect 300308 64184 300360 64190
rect 300308 64126 300360 64132
rect 300216 51808 300268 51814
rect 300216 51750 300268 51756
rect 300768 39500 300820 39506
rect 300768 39442 300820 39448
rect 300780 38690 300808 39442
rect 300768 38684 300820 38690
rect 300768 38626 300820 38632
rect 300124 38004 300176 38010
rect 300124 37946 300176 37952
rect 299480 37936 299532 37942
rect 299480 37878 299532 37884
rect 298836 28960 298888 28966
rect 298836 28902 298888 28908
rect 298744 21480 298796 21486
rect 298744 21422 298796 21428
rect 299492 16574 299520 37878
rect 299492 16546 299704 16574
rect 299676 480 299704 16546
rect 300768 4140 300820 4146
rect 300768 4082 300820 4088
rect 300780 480 300808 4082
rect 301516 2174 301544 129882
rect 301608 125458 301636 164290
rect 302896 135250 302924 172654
rect 307312 172582 307340 173567
rect 307300 172576 307352 172582
rect 307300 172518 307352 172524
rect 306746 172272 306802 172281
rect 306746 172207 306802 172216
rect 306760 171134 306788 172207
rect 307114 171864 307170 171873
rect 307404 171834 307432 175199
rect 307574 174856 307630 174865
rect 307574 174791 307630 174800
rect 307482 174448 307538 174457
rect 307482 174383 307538 174392
rect 307496 173942 307524 174383
rect 307588 174078 307616 174791
rect 307576 174072 307628 174078
rect 307576 174014 307628 174020
rect 307666 174040 307722 174049
rect 307666 173975 307668 173984
rect 307720 173975 307722 173984
rect 307668 173946 307720 173952
rect 307484 173936 307536 173942
rect 307484 173878 307536 173884
rect 307482 173224 307538 173233
rect 307482 173159 307538 173168
rect 307496 172718 307524 173159
rect 307484 172712 307536 172718
rect 307484 172654 307536 172660
rect 307666 172680 307722 172689
rect 307666 172615 307668 172624
rect 307720 172615 307722 172624
rect 307668 172586 307720 172592
rect 307114 171799 307170 171808
rect 307392 171828 307444 171834
rect 307128 171154 307156 171799
rect 307392 171770 307444 171776
rect 307666 171456 307722 171465
rect 307666 171391 307722 171400
rect 307680 171222 307708 171391
rect 307668 171216 307720 171222
rect 307668 171158 307720 171164
rect 306668 171106 306788 171134
rect 307116 171148 307168 171154
rect 306562 168872 306618 168881
rect 306562 168807 306618 168816
rect 306576 167686 306604 168807
rect 306564 167680 306616 167686
rect 306564 167622 306616 167628
rect 306562 166424 306618 166433
rect 306668 166394 306696 171106
rect 307116 171090 307168 171096
rect 306746 171048 306802 171057
rect 306746 170983 306802 170992
rect 306760 169930 306788 170983
rect 306930 170640 306986 170649
rect 306930 170575 306986 170584
rect 306748 169924 306800 169930
rect 306748 169866 306800 169872
rect 306746 166832 306802 166841
rect 306746 166767 306802 166776
rect 306562 166359 306618 166368
rect 306656 166388 306708 166394
rect 306576 163606 306604 166359
rect 306656 166330 306708 166336
rect 306760 165646 306788 166767
rect 306944 166326 306972 170575
rect 307666 170232 307722 170241
rect 307666 170167 307722 170176
rect 307680 169862 307708 170167
rect 307668 169856 307720 169862
rect 307482 169824 307538 169833
rect 307668 169798 307720 169804
rect 307482 169759 307484 169768
rect 307536 169759 307538 169768
rect 307484 169730 307536 169736
rect 307574 169280 307630 169289
rect 307574 169215 307630 169224
rect 307588 168434 307616 169215
rect 307668 168496 307720 168502
rect 307666 168464 307668 168473
rect 307720 168464 307722 168473
rect 307576 168428 307628 168434
rect 307666 168399 307722 168408
rect 307576 168370 307628 168376
rect 307298 168056 307354 168065
rect 307298 167991 307354 168000
rect 307312 167074 307340 167991
rect 307574 167648 307630 167657
rect 307574 167583 307630 167592
rect 307300 167068 307352 167074
rect 307300 167010 307352 167016
rect 306932 166320 306984 166326
rect 306932 166262 306984 166268
rect 307482 165880 307538 165889
rect 307482 165815 307538 165824
rect 306748 165640 306800 165646
rect 306748 165582 306800 165588
rect 307206 165472 307262 165481
rect 307206 165407 307262 165416
rect 307022 165064 307078 165073
rect 307022 164999 307078 165008
rect 306930 163840 306986 163849
rect 306930 163775 306986 163784
rect 306564 163600 306616 163606
rect 306564 163542 306616 163548
rect 306944 163033 306972 163775
rect 305642 163024 305698 163033
rect 305642 162959 305698 162968
rect 306930 163024 306986 163033
rect 306930 162959 306986 162968
rect 302976 161696 303028 161702
rect 302976 161638 303028 161644
rect 302884 135244 302936 135250
rect 302884 135186 302936 135192
rect 301596 125452 301648 125458
rect 301596 125394 301648 125400
rect 301688 124364 301740 124370
rect 301688 124306 301740 124312
rect 301596 100972 301648 100978
rect 301596 100914 301648 100920
rect 301504 2168 301556 2174
rect 301504 2110 301556 2116
rect 301608 2106 301636 100914
rect 301700 35290 301728 124306
rect 302988 124166 303016 161638
rect 304356 154760 304408 154766
rect 304356 154702 304408 154708
rect 304368 149705 304396 154702
rect 304354 149696 304410 149705
rect 304354 149631 304410 149640
rect 304264 149252 304316 149258
rect 304264 149194 304316 149200
rect 303158 143984 303214 143993
rect 303158 143919 303214 143928
rect 302976 124160 303028 124166
rect 302976 124102 303028 124108
rect 303068 122868 303120 122874
rect 303068 122810 303120 122816
rect 302884 109132 302936 109138
rect 302884 109074 302936 109080
rect 302240 39568 302292 39574
rect 302240 39510 302292 39516
rect 302252 39370 302280 39510
rect 302240 39364 302292 39370
rect 302240 39306 302292 39312
rect 301688 35284 301740 35290
rect 301688 35226 301740 35232
rect 302252 16574 302280 39306
rect 302896 24274 302924 109074
rect 302976 107704 303028 107710
rect 302976 107646 303028 107652
rect 302988 40730 303016 107646
rect 303080 62898 303108 122810
rect 303172 103494 303200 143919
rect 304276 112470 304304 149194
rect 304356 140956 304408 140962
rect 304356 140898 304408 140904
rect 304368 119406 304396 140898
rect 304448 129872 304500 129878
rect 304448 129814 304500 129820
rect 304356 119400 304408 119406
rect 304356 119342 304408 119348
rect 304264 112464 304316 112470
rect 304264 112406 304316 112412
rect 304356 111920 304408 111926
rect 304356 111862 304408 111868
rect 304264 106480 304316 106486
rect 304264 106422 304316 106428
rect 303160 103488 303212 103494
rect 303160 103430 303212 103436
rect 303068 62892 303120 62898
rect 303068 62834 303120 62840
rect 302976 40724 303028 40730
rect 302976 40666 303028 40672
rect 302884 24268 302936 24274
rect 302884 24210 302936 24216
rect 302252 16546 303200 16574
rect 301780 7676 301832 7682
rect 301780 7618 301832 7624
rect 301792 6798 301820 7618
rect 301780 6792 301832 6798
rect 301780 6734 301832 6740
rect 301596 2100 301648 2106
rect 301596 2042 301648 2048
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301792 354 301820 6734
rect 303172 480 303200 16546
rect 304276 15910 304304 106422
rect 304368 32502 304396 111862
rect 304460 58750 304488 129814
rect 305656 127634 305684 162959
rect 306562 161256 306618 161265
rect 306562 161191 306618 161200
rect 306576 160138 306604 161191
rect 306564 160132 306616 160138
rect 306564 160074 306616 160080
rect 306930 160032 306986 160041
rect 306930 159967 306986 159976
rect 306944 158914 306972 159967
rect 306932 158908 306984 158914
rect 306932 158850 306984 158856
rect 306746 158264 306802 158273
rect 306746 158199 306802 158208
rect 306760 157418 306788 158199
rect 306748 157412 306800 157418
rect 306748 157354 306800 157360
rect 306562 157040 306618 157049
rect 306562 156975 306618 156984
rect 306576 155990 306604 156975
rect 306564 155984 306616 155990
rect 306564 155926 306616 155932
rect 306562 155680 306618 155689
rect 306562 155615 306618 155624
rect 306576 154698 306604 155615
rect 306564 154692 306616 154698
rect 306564 154634 306616 154640
rect 306654 153640 306710 153649
rect 306654 153575 306710 153584
rect 306668 151094 306696 153575
rect 306656 151088 306708 151094
rect 306656 151030 306708 151036
rect 305826 150648 305882 150657
rect 305826 150583 305882 150592
rect 305644 127628 305696 127634
rect 305644 127570 305696 127576
rect 305734 118824 305790 118833
rect 305734 118759 305790 118768
rect 304540 117496 304592 117502
rect 304540 117438 304592 117444
rect 304552 69698 304580 117438
rect 305642 109304 305698 109313
rect 305642 109239 305698 109248
rect 304540 69692 304592 69698
rect 304540 69634 304592 69640
rect 304448 58744 304500 58750
rect 304448 58686 304500 58692
rect 304356 32496 304408 32502
rect 304356 32438 304408 32444
rect 304264 15904 304316 15910
rect 304264 15846 304316 15852
rect 305552 10396 305604 10402
rect 305552 10338 305604 10344
rect 304354 3496 304410 3505
rect 304354 3431 304410 3440
rect 304368 480 304396 3431
rect 305564 480 305592 10338
rect 305656 6254 305684 109239
rect 305748 17338 305776 118759
rect 305840 110430 305868 150583
rect 306746 150240 306802 150249
rect 306746 150175 306802 150184
rect 306760 149190 306788 150175
rect 306748 149184 306800 149190
rect 306748 149126 306800 149132
rect 306930 148472 306986 148481
rect 306930 148407 306986 148416
rect 306944 147830 306972 148407
rect 306932 147824 306984 147830
rect 306932 147766 306984 147772
rect 306746 146840 306802 146849
rect 306746 146775 306802 146784
rect 306760 146334 306788 146775
rect 306748 146328 306800 146334
rect 306748 146270 306800 146276
rect 306930 144256 306986 144265
rect 306930 144191 306986 144200
rect 306944 143614 306972 144191
rect 306932 143608 306984 143614
rect 306932 143550 306984 143556
rect 306562 143032 306618 143041
rect 306562 142967 306618 142976
rect 306576 142186 306604 142967
rect 306564 142180 306616 142186
rect 306564 142122 306616 142128
rect 306562 142080 306618 142089
rect 306562 142015 306618 142024
rect 306576 140894 306604 142015
rect 307036 141438 307064 164999
rect 307116 164348 307168 164354
rect 307116 164290 307168 164296
rect 307128 164257 307156 164290
rect 307114 164248 307170 164257
rect 307114 164183 307170 164192
rect 307220 158030 307248 165407
rect 307496 164898 307524 165815
rect 307484 164892 307536 164898
rect 307484 164834 307536 164840
rect 307588 163538 307616 167583
rect 307666 167240 307722 167249
rect 307666 167175 307722 167184
rect 307680 167142 307708 167175
rect 307668 167136 307720 167142
rect 307668 167078 307720 167084
rect 307666 164656 307722 164665
rect 307666 164591 307722 164600
rect 307680 164286 307708 164591
rect 307668 164280 307720 164286
rect 307668 164222 307720 164228
rect 307576 163532 307628 163538
rect 307576 163474 307628 163480
rect 307390 163432 307446 163441
rect 307390 163367 307446 163376
rect 307404 161702 307432 163367
rect 307666 163024 307722 163033
rect 307666 162959 307722 162968
rect 307680 162926 307708 162959
rect 307668 162920 307720 162926
rect 307668 162862 307720 162868
rect 307482 162480 307538 162489
rect 307482 162415 307538 162424
rect 307392 161696 307444 161702
rect 307392 161638 307444 161644
rect 307496 161634 307524 162415
rect 307574 162072 307630 162081
rect 307574 162007 307630 162016
rect 307484 161628 307536 161634
rect 307484 161570 307536 161576
rect 307588 161566 307616 162007
rect 307666 161664 307722 161673
rect 307666 161599 307722 161608
rect 307576 161560 307628 161566
rect 307576 161502 307628 161508
rect 307680 161498 307708 161599
rect 307668 161492 307720 161498
rect 307668 161434 307720 161440
rect 307574 160848 307630 160857
rect 307574 160783 307630 160792
rect 307588 160274 307616 160783
rect 307666 160440 307722 160449
rect 307666 160375 307722 160384
rect 307576 160268 307628 160274
rect 307576 160210 307628 160216
rect 307680 160206 307708 160375
rect 307668 160200 307720 160206
rect 307668 160142 307720 160148
rect 307574 159624 307630 159633
rect 307574 159559 307630 159568
rect 307588 158778 307616 159559
rect 307666 159080 307722 159089
rect 307666 159015 307722 159024
rect 307680 158846 307708 159015
rect 307668 158840 307720 158846
rect 307668 158782 307720 158788
rect 307576 158772 307628 158778
rect 307576 158714 307628 158720
rect 307390 158672 307446 158681
rect 307390 158607 307446 158616
rect 307208 158024 307260 158030
rect 307208 157966 307260 157972
rect 307114 157448 307170 157457
rect 307114 157383 307170 157392
rect 307128 145586 307156 157383
rect 307298 154864 307354 154873
rect 307298 154799 307354 154808
rect 307312 154630 307340 154799
rect 307300 154624 307352 154630
rect 307300 154566 307352 154572
rect 307298 154456 307354 154465
rect 307298 154391 307354 154400
rect 307312 153270 307340 154391
rect 307300 153264 307352 153270
rect 307300 153206 307352 153212
rect 307404 151814 307432 158607
rect 307482 157856 307538 157865
rect 307482 157791 307538 157800
rect 307496 157486 307524 157791
rect 307484 157480 307536 157486
rect 307484 157422 307536 157428
rect 307574 156632 307630 156641
rect 307574 156567 307630 156576
rect 307588 156058 307616 156567
rect 307666 156224 307722 156233
rect 307666 156159 307722 156168
rect 307680 156126 307708 156159
rect 307668 156120 307720 156126
rect 307668 156062 307720 156068
rect 307576 156052 307628 156058
rect 307576 155994 307628 156000
rect 307666 155272 307722 155281
rect 307666 155207 307722 155216
rect 307680 154766 307708 155207
rect 307668 154760 307720 154766
rect 307668 154702 307720 154708
rect 307574 154048 307630 154057
rect 307574 153983 307630 153992
rect 307588 153406 307616 153983
rect 307576 153400 307628 153406
rect 307576 153342 307628 153348
rect 307668 153332 307720 153338
rect 307668 153274 307720 153280
rect 307680 153241 307708 153274
rect 307666 153232 307722 153241
rect 307666 153167 307722 153176
rect 307482 152688 307538 152697
rect 307482 152623 307538 152632
rect 307496 151842 307524 152623
rect 307574 152280 307630 152289
rect 307574 152215 307630 152224
rect 307588 151910 307616 152215
rect 307668 151972 307720 151978
rect 307668 151914 307720 151920
rect 307576 151904 307628 151910
rect 307680 151881 307708 151914
rect 307576 151846 307628 151852
rect 307666 151872 307722 151881
rect 307220 151786 307432 151814
rect 307484 151836 307536 151842
rect 307116 145580 307168 145586
rect 307116 145522 307168 145528
rect 307114 142488 307170 142497
rect 307114 142423 307170 142432
rect 307024 141432 307076 141438
rect 307024 141374 307076 141380
rect 306564 140888 306616 140894
rect 306564 140830 306616 140836
rect 306562 139088 306618 139097
rect 306562 139023 306618 139032
rect 306576 138106 306604 139023
rect 306564 138100 306616 138106
rect 306564 138042 306616 138048
rect 306562 136640 306618 136649
rect 306562 136575 306618 136584
rect 306576 135318 306604 136575
rect 306564 135312 306616 135318
rect 306564 135254 306616 135260
rect 306562 134872 306618 134881
rect 306562 134807 306618 134816
rect 306576 133958 306604 134807
rect 307022 134056 307078 134065
rect 307022 133991 307078 134000
rect 306564 133952 306616 133958
rect 306564 133894 306616 133900
rect 306562 133648 306618 133657
rect 306562 133583 306618 133592
rect 306576 132530 306604 133583
rect 306930 133240 306986 133249
rect 306930 133175 306986 133184
rect 306944 132666 306972 133175
rect 306932 132660 306984 132666
rect 306932 132602 306984 132608
rect 306564 132524 306616 132530
rect 306564 132466 306616 132472
rect 306562 131064 306618 131073
rect 306562 130999 306618 131008
rect 306576 129810 306604 130999
rect 306930 130656 306986 130665
rect 306930 130591 306986 130600
rect 306944 129878 306972 130591
rect 306932 129872 306984 129878
rect 306932 129814 306984 129820
rect 306564 129804 306616 129810
rect 306564 129746 306616 129752
rect 306930 129296 306986 129305
rect 306930 129231 306986 129240
rect 306944 128450 306972 129231
rect 306932 128444 306984 128450
rect 306932 128386 306984 128392
rect 305918 123312 305974 123321
rect 305918 123247 305974 123256
rect 305828 110424 305880 110430
rect 305828 110366 305880 110372
rect 305826 108352 305882 108361
rect 305826 108287 305882 108296
rect 305840 43450 305868 108287
rect 305932 76566 305960 123247
rect 306562 118688 306618 118697
rect 306562 118623 306618 118632
rect 306576 117434 306604 118623
rect 306564 117428 306616 117434
rect 306564 117370 306616 117376
rect 306746 116648 306802 116657
rect 306746 116583 306802 116592
rect 306760 116142 306788 116583
rect 306748 116136 306800 116142
rect 306748 116078 306800 116084
rect 306930 112704 306986 112713
rect 306930 112639 306986 112648
rect 306944 111858 306972 112639
rect 306932 111852 306984 111858
rect 306932 111794 306984 111800
rect 306746 110256 306802 110265
rect 306746 110191 306802 110200
rect 306760 109313 306788 110191
rect 306746 109304 306802 109313
rect 306746 109239 306802 109248
rect 306930 109304 306986 109313
rect 306930 109239 306986 109248
rect 306944 109138 306972 109239
rect 306932 109132 306984 109138
rect 306932 109074 306984 109080
rect 306930 105904 306986 105913
rect 306930 105839 306986 105848
rect 306944 104922 306972 105839
rect 306932 104916 306984 104922
rect 306932 104858 306984 104864
rect 306930 104680 306986 104689
rect 306930 104615 306986 104624
rect 306944 103698 306972 104615
rect 306932 103692 306984 103698
rect 306932 103634 306984 103640
rect 306562 101280 306618 101289
rect 306562 101215 306618 101224
rect 306576 100978 306604 101215
rect 306564 100972 306616 100978
rect 306564 100914 306616 100920
rect 306930 100872 306986 100881
rect 306930 100807 306986 100816
rect 306944 100774 306972 100807
rect 306932 100768 306984 100774
rect 306932 100710 306984 100716
rect 306562 100464 306618 100473
rect 306562 100399 306618 100408
rect 306576 99550 306604 100399
rect 306564 99544 306616 99550
rect 306564 99486 306616 99492
rect 306930 98696 306986 98705
rect 306930 98631 306986 98640
rect 306944 98190 306972 98631
rect 306932 98184 306984 98190
rect 306932 98126 306984 98132
rect 305920 76560 305972 76566
rect 305920 76502 305972 76508
rect 305828 43444 305880 43450
rect 305828 43386 305880 43392
rect 307036 18766 307064 133991
rect 307128 119474 307156 142423
rect 307220 137290 307248 151786
rect 307666 151807 307722 151816
rect 307484 151778 307536 151784
rect 307574 151464 307630 151473
rect 307574 151399 307630 151408
rect 307588 150618 307616 151399
rect 307666 151056 307722 151065
rect 307666 150991 307722 151000
rect 307576 150612 307628 150618
rect 307576 150554 307628 150560
rect 307680 150550 307708 150991
rect 307668 150544 307720 150550
rect 307668 150486 307720 150492
rect 307666 149832 307722 149841
rect 307666 149767 307722 149776
rect 307574 149288 307630 149297
rect 307680 149258 307708 149767
rect 307574 149223 307630 149232
rect 307668 149252 307720 149258
rect 307588 149122 307616 149223
rect 307668 149194 307720 149200
rect 307576 149116 307628 149122
rect 307576 149058 307628 149064
rect 307574 148880 307630 148889
rect 307574 148815 307630 148824
rect 307588 147762 307616 148815
rect 307666 148064 307722 148073
rect 307666 147999 307722 148008
rect 307576 147756 307628 147762
rect 307576 147698 307628 147704
rect 307680 147694 307708 147999
rect 307668 147688 307720 147694
rect 307390 147656 307446 147665
rect 307668 147630 307720 147636
rect 307390 147591 307446 147600
rect 307298 139632 307354 139641
rect 307298 139567 307354 139576
rect 307312 139466 307340 139567
rect 307300 139460 307352 139466
rect 307300 139402 307352 139408
rect 307298 138680 307354 138689
rect 307298 138615 307354 138624
rect 307312 138174 307340 138615
rect 307300 138168 307352 138174
rect 307300 138110 307352 138116
rect 307208 137284 307260 137290
rect 307208 137226 307260 137232
rect 307206 137048 307262 137057
rect 307206 136983 307262 136992
rect 307116 119468 307168 119474
rect 307116 119410 307168 119416
rect 307114 114064 307170 114073
rect 307114 113999 307170 114008
rect 307128 19990 307156 113999
rect 307220 84862 307248 136983
rect 307300 135448 307352 135454
rect 307300 135390 307352 135396
rect 307312 135289 307340 135390
rect 307298 135280 307354 135289
rect 307298 135215 307354 135224
rect 307404 134570 307432 147591
rect 307574 147248 307630 147257
rect 307574 147183 307630 147192
rect 307588 146470 307616 147183
rect 307576 146464 307628 146470
rect 307576 146406 307628 146412
rect 307666 146432 307722 146441
rect 307666 146367 307668 146376
rect 307720 146367 307722 146376
rect 307668 146338 307720 146344
rect 307666 145888 307722 145897
rect 307666 145823 307722 145832
rect 307574 145480 307630 145489
rect 307574 145415 307630 145424
rect 307588 144226 307616 145415
rect 307680 144974 307708 145823
rect 307668 144968 307720 144974
rect 307668 144910 307720 144916
rect 307666 144664 307722 144673
rect 307666 144599 307722 144608
rect 307576 144220 307628 144226
rect 307576 144162 307628 144168
rect 307574 143848 307630 143857
rect 307574 143783 307630 143792
rect 307588 142866 307616 143783
rect 307680 143682 307708 144599
rect 307668 143676 307720 143682
rect 307668 143618 307720 143624
rect 307666 143440 307722 143449
rect 307666 143375 307722 143384
rect 307576 142860 307628 142866
rect 307576 142802 307628 142808
rect 307680 142254 307708 143375
rect 307668 142248 307720 142254
rect 307668 142190 307720 142196
rect 307574 141672 307630 141681
rect 307574 141607 307630 141616
rect 307482 141264 307538 141273
rect 307482 141199 307538 141208
rect 307496 140962 307524 141199
rect 307484 140956 307536 140962
rect 307484 140898 307536 140904
rect 307588 140570 307616 141607
rect 307666 140856 307722 140865
rect 307666 140791 307668 140800
rect 307720 140791 307722 140800
rect 307668 140762 307720 140768
rect 307496 140542 307616 140570
rect 307392 134564 307444 134570
rect 307392 134506 307444 134512
rect 307298 132696 307354 132705
rect 307298 132631 307354 132640
rect 307312 132598 307340 132631
rect 307300 132592 307352 132598
rect 307300 132534 307352 132540
rect 307496 132494 307524 140542
rect 307574 140448 307630 140457
rect 307574 140383 307630 140392
rect 307588 139534 307616 140383
rect 307666 140040 307722 140049
rect 307666 139975 307722 139984
rect 307680 139602 307708 139975
rect 307668 139596 307720 139602
rect 307668 139538 307720 139544
rect 307576 139528 307628 139534
rect 307576 139470 307628 139476
rect 307666 138272 307722 138281
rect 307666 138207 307722 138216
rect 307680 138038 307708 138207
rect 307668 138032 307720 138038
rect 307668 137974 307720 137980
rect 307666 137864 307722 137873
rect 307666 137799 307722 137808
rect 307680 136678 307708 137799
rect 307668 136672 307720 136678
rect 307668 136614 307720 136620
rect 307574 136232 307630 136241
rect 307574 136167 307630 136176
rect 307588 135386 307616 136167
rect 307666 135688 307722 135697
rect 307666 135623 307722 135632
rect 307680 135522 307708 135623
rect 307668 135516 307720 135522
rect 307668 135458 307720 135464
rect 307576 135380 307628 135386
rect 307576 135322 307628 135328
rect 307404 132466 307524 132494
rect 307404 127702 307432 132466
rect 307482 132288 307538 132297
rect 307482 132223 307538 132232
rect 307496 131306 307524 132223
rect 307574 131880 307630 131889
rect 307574 131815 307630 131824
rect 307484 131300 307536 131306
rect 307484 131242 307536 131248
rect 307588 131238 307616 131815
rect 307666 131472 307722 131481
rect 307666 131407 307722 131416
rect 307576 131232 307628 131238
rect 307576 131174 307628 131180
rect 307680 131170 307708 131407
rect 307668 131164 307720 131170
rect 307668 131106 307720 131112
rect 307484 129940 307536 129946
rect 307484 129882 307536 129888
rect 307496 129849 307524 129882
rect 307482 129840 307538 129849
rect 307482 129775 307538 129784
rect 307666 128888 307722 128897
rect 307666 128823 307722 128832
rect 307680 128518 307708 128823
rect 307668 128512 307720 128518
rect 307574 128480 307630 128489
rect 307668 128454 307720 128460
rect 307574 128415 307630 128424
rect 307588 128382 307616 128415
rect 307576 128376 307628 128382
rect 307576 128318 307628 128324
rect 307574 128072 307630 128081
rect 307574 128007 307630 128016
rect 307392 127696 307444 127702
rect 307392 127638 307444 127644
rect 307588 127090 307616 128007
rect 307666 127256 307722 127265
rect 307666 127191 307722 127200
rect 307576 127084 307628 127090
rect 307576 127026 307628 127032
rect 307680 127022 307708 127191
rect 307668 127016 307720 127022
rect 307668 126958 307720 126964
rect 307482 126848 307538 126857
rect 307482 126783 307538 126792
rect 307496 125730 307524 126783
rect 307574 126440 307630 126449
rect 307574 126375 307630 126384
rect 307484 125724 307536 125730
rect 307484 125666 307536 125672
rect 307588 125662 307616 126375
rect 307666 125896 307722 125905
rect 307666 125831 307722 125840
rect 307680 125798 307708 125831
rect 307668 125792 307720 125798
rect 307668 125734 307720 125740
rect 307576 125656 307628 125662
rect 307576 125598 307628 125604
rect 307482 125488 307538 125497
rect 307482 125423 307538 125432
rect 307298 124264 307354 124273
rect 307496 124234 307524 125423
rect 307574 125080 307630 125089
rect 307574 125015 307630 125024
rect 307588 124302 307616 125015
rect 307666 124672 307722 124681
rect 307666 124607 307722 124616
rect 307680 124370 307708 124607
rect 307668 124364 307720 124370
rect 307668 124306 307720 124312
rect 307576 124296 307628 124302
rect 307576 124238 307628 124244
rect 307298 124199 307354 124208
rect 307484 124228 307536 124234
rect 307312 89010 307340 124199
rect 307484 124170 307536 124176
rect 307574 123856 307630 123865
rect 307574 123791 307630 123800
rect 307588 123010 307616 123791
rect 307666 123040 307722 123049
rect 307576 123004 307628 123010
rect 307666 122975 307722 122984
rect 307576 122946 307628 122952
rect 307680 122874 307708 122975
rect 307668 122868 307720 122874
rect 307668 122810 307720 122816
rect 307482 122496 307538 122505
rect 307482 122431 307538 122440
rect 307496 121582 307524 122431
rect 307666 122088 307722 122097
rect 307666 122023 307722 122032
rect 307574 121680 307630 121689
rect 307680 121650 307708 122023
rect 307574 121615 307630 121624
rect 307668 121644 307720 121650
rect 307484 121576 307536 121582
rect 307484 121518 307536 121524
rect 307588 121514 307616 121615
rect 307668 121586 307720 121592
rect 307576 121508 307628 121514
rect 307576 121450 307628 121456
rect 307482 121272 307538 121281
rect 307482 121207 307538 121216
rect 307496 120222 307524 121207
rect 307666 120864 307722 120873
rect 307666 120799 307722 120808
rect 307574 120456 307630 120465
rect 307574 120391 307630 120400
rect 307484 120216 307536 120222
rect 307484 120158 307536 120164
rect 307588 120154 307616 120391
rect 307680 120290 307708 120799
rect 307668 120284 307720 120290
rect 307668 120226 307720 120232
rect 307576 120148 307628 120154
rect 307576 120090 307628 120096
rect 307482 120048 307538 120057
rect 307482 119983 307538 119992
rect 307496 118726 307524 119983
rect 307574 119640 307630 119649
rect 307574 119575 307630 119584
rect 307588 118833 307616 119575
rect 307666 119096 307722 119105
rect 307666 119031 307722 119040
rect 307680 118862 307708 119031
rect 307668 118856 307720 118862
rect 307574 118824 307630 118833
rect 307668 118798 307720 118804
rect 307574 118759 307630 118768
rect 307484 118720 307536 118726
rect 307484 118662 307536 118668
rect 307574 117872 307630 117881
rect 307574 117807 307630 117816
rect 307588 117502 307616 117807
rect 307576 117496 307628 117502
rect 307576 117438 307628 117444
rect 307666 117464 307722 117473
rect 307666 117399 307722 117408
rect 307680 117366 307708 117399
rect 307668 117360 307720 117366
rect 307668 117302 307720 117308
rect 307574 117056 307630 117065
rect 307574 116991 307630 117000
rect 307588 116006 307616 116991
rect 307666 116240 307722 116249
rect 307666 116175 307722 116184
rect 307680 116074 307708 116175
rect 307668 116068 307720 116074
rect 307668 116010 307720 116016
rect 307576 116000 307628 116006
rect 307576 115942 307628 115948
rect 307482 115696 307538 115705
rect 307482 115631 307538 115640
rect 307496 114578 307524 115631
rect 307574 115288 307630 115297
rect 307574 115223 307630 115232
rect 307588 114646 307616 115223
rect 307666 114880 307722 114889
rect 307666 114815 307722 114824
rect 307680 114714 307708 114815
rect 307668 114708 307720 114714
rect 307668 114650 307720 114656
rect 307576 114640 307628 114646
rect 307576 114582 307628 114588
rect 307484 114572 307536 114578
rect 307484 114514 307536 114520
rect 307666 114472 307722 114481
rect 307666 114407 307722 114416
rect 307574 113656 307630 113665
rect 307574 113591 307630 113600
rect 307588 113286 307616 113591
rect 307680 113354 307708 114407
rect 307668 113348 307720 113354
rect 307668 113290 307720 113296
rect 307576 113280 307628 113286
rect 307576 113222 307628 113228
rect 307666 113248 307722 113257
rect 307666 113183 307668 113192
rect 307720 113183 307722 113192
rect 307668 113154 307720 113160
rect 307668 111920 307720 111926
rect 307666 111888 307668 111897
rect 307720 111888 307722 111897
rect 307666 111823 307722 111832
rect 307482 111480 307538 111489
rect 307482 111415 307538 111424
rect 307496 110634 307524 111415
rect 307574 111072 307630 111081
rect 307574 111007 307630 111016
rect 307484 110628 307536 110634
rect 307484 110570 307536 110576
rect 307588 110566 307616 111007
rect 307666 110664 307722 110673
rect 307666 110599 307722 110608
rect 307576 110560 307628 110566
rect 307576 110502 307628 110508
rect 307680 110498 307708 110599
rect 307668 110492 307720 110498
rect 307668 110434 307720 110440
rect 307666 109848 307722 109857
rect 307666 109783 307722 109792
rect 307680 109070 307708 109783
rect 307668 109064 307720 109070
rect 307668 109006 307720 109012
rect 307574 108896 307630 108905
rect 307574 108831 307630 108840
rect 307588 107710 307616 108831
rect 307666 108080 307722 108089
rect 307666 108015 307722 108024
rect 307680 107914 307708 108015
rect 307668 107908 307720 107914
rect 307668 107850 307720 107856
rect 307668 107772 307720 107778
rect 307668 107714 307720 107720
rect 307576 107704 307628 107710
rect 307680 107681 307708 107714
rect 307576 107646 307628 107652
rect 307666 107672 307722 107681
rect 307666 107607 307722 107616
rect 307574 107264 307630 107273
rect 307574 107199 307630 107208
rect 307482 106856 307538 106865
rect 307482 106791 307538 106800
rect 307496 106418 307524 106791
rect 307588 106486 307616 107199
rect 307576 106480 307628 106486
rect 307576 106422 307628 106428
rect 307666 106448 307722 106457
rect 307484 106412 307536 106418
rect 307666 106383 307722 106392
rect 307484 106354 307536 106360
rect 307680 106350 307708 106383
rect 307668 106344 307720 106350
rect 307668 106286 307720 106292
rect 307482 105496 307538 105505
rect 307482 105431 307538 105440
rect 307496 105058 307524 105431
rect 307666 105088 307722 105097
rect 307484 105052 307536 105058
rect 307666 105023 307722 105032
rect 307484 104994 307536 105000
rect 307680 104990 307708 105023
rect 307668 104984 307720 104990
rect 307668 104926 307720 104932
rect 307574 104272 307630 104281
rect 307574 104207 307630 104216
rect 307588 103562 307616 104207
rect 307666 103864 307722 103873
rect 307666 103799 307722 103808
rect 307680 103630 307708 103799
rect 307668 103624 307720 103630
rect 307668 103566 307720 103572
rect 307576 103556 307628 103562
rect 307576 103498 307628 103504
rect 307574 103456 307630 103465
rect 307574 103391 307630 103400
rect 307588 102202 307616 103391
rect 307666 102504 307722 102513
rect 307666 102439 307722 102448
rect 307680 102270 307708 102439
rect 307668 102264 307720 102270
rect 307668 102206 307720 102212
rect 307576 102196 307628 102202
rect 307576 102138 307628 102144
rect 307666 102096 307722 102105
rect 307666 102031 307722 102040
rect 307574 101688 307630 101697
rect 307574 101623 307630 101632
rect 307588 100842 307616 101623
rect 307680 100910 307708 102031
rect 307668 100904 307720 100910
rect 307668 100846 307720 100852
rect 307576 100836 307628 100842
rect 307576 100778 307628 100784
rect 307574 100056 307630 100065
rect 307574 99991 307630 100000
rect 307588 99414 307616 99991
rect 307666 99648 307722 99657
rect 307666 99583 307722 99592
rect 307680 99482 307708 99583
rect 307668 99476 307720 99482
rect 307668 99418 307720 99424
rect 307576 99408 307628 99414
rect 307576 99350 307628 99356
rect 307574 99104 307630 99113
rect 307574 99039 307630 99048
rect 307588 98122 307616 99039
rect 307666 98288 307722 98297
rect 307666 98223 307722 98232
rect 307576 98116 307628 98122
rect 307576 98058 307628 98064
rect 307680 98054 307708 98223
rect 307668 98048 307720 98054
rect 307668 97990 307720 97996
rect 307482 97880 307538 97889
rect 307482 97815 307538 97824
rect 307496 96694 307524 97815
rect 307668 96756 307720 96762
rect 307668 96698 307720 96704
rect 307484 96688 307536 96694
rect 307680 96665 307708 96698
rect 307484 96630 307536 96636
rect 307666 96656 307722 96665
rect 307666 96591 307722 96600
rect 308416 96490 308444 187274
rect 308494 178120 308550 178129
rect 308494 178055 308550 178064
rect 308508 123457 308536 178055
rect 308494 123448 308550 123457
rect 308494 123383 308550 123392
rect 308496 122120 308548 122126
rect 308496 122062 308548 122068
rect 308404 96484 308456 96490
rect 308404 96426 308456 96432
rect 307666 96248 307722 96257
rect 307666 96183 307722 96192
rect 307680 95266 307708 96183
rect 307668 95260 307720 95266
rect 307668 95202 307720 95208
rect 308508 94926 308536 122062
rect 309138 112296 309194 112305
rect 309138 112231 309194 112240
rect 308496 94920 308548 94926
rect 308496 94862 308548 94868
rect 307300 89004 307352 89010
rect 307300 88946 307352 88952
rect 308404 86352 308456 86358
rect 308404 86294 308456 86300
rect 307208 84856 307260 84862
rect 307208 84798 307260 84804
rect 307208 76560 307260 76566
rect 307208 76502 307260 76508
rect 307220 38690 307248 76502
rect 307208 38684 307260 38690
rect 307208 38626 307260 38632
rect 307116 19984 307168 19990
rect 307116 19926 307168 19932
rect 307024 18760 307076 18766
rect 307024 18702 307076 18708
rect 305736 17332 305788 17338
rect 305736 17274 305788 17280
rect 306748 6928 306800 6934
rect 306748 6870 306800 6876
rect 305644 6248 305696 6254
rect 305644 6190 305696 6196
rect 306760 480 306788 6870
rect 307220 4146 307248 38626
rect 308416 27606 308444 86294
rect 309152 73846 309180 112231
rect 309796 96558 309824 190062
rect 309888 179042 309916 222090
rect 309876 179036 309928 179042
rect 309876 178978 309928 178984
rect 312556 177682 312584 237390
rect 313292 223582 313320 239822
rect 316604 238746 316632 240040
rect 316592 238740 316644 238746
rect 316592 238682 316644 238688
rect 314108 238128 314160 238134
rect 314108 238070 314160 238076
rect 314016 225752 314068 225758
rect 314016 225694 314068 225700
rect 313280 223576 313332 223582
rect 313280 223518 313332 223524
rect 313924 223576 313976 223582
rect 313924 223518 313976 223524
rect 313832 182980 313884 182986
rect 313832 182922 313884 182928
rect 312544 177676 312596 177682
rect 312544 177618 312596 177624
rect 313844 176662 313872 182922
rect 313936 178974 313964 223518
rect 314028 182850 314056 225694
rect 314120 220794 314148 238070
rect 316604 238066 316632 238682
rect 316592 238060 316644 238066
rect 316592 238002 316644 238008
rect 318536 237454 318564 240094
rect 318064 237448 318116 237454
rect 318064 237390 318116 237396
rect 318524 237448 318576 237454
rect 318524 237390 318576 237396
rect 316684 233912 316736 233918
rect 316684 233854 316736 233860
rect 314108 220788 314160 220794
rect 314108 220730 314160 220736
rect 314016 182844 314068 182850
rect 314016 182786 314068 182792
rect 316696 180794 316724 233854
rect 318076 224942 318104 237390
rect 318708 233980 318760 233986
rect 318708 233922 318760 233928
rect 318064 224936 318116 224942
rect 318064 224878 318116 224884
rect 318064 192704 318116 192710
rect 318064 192646 318116 192652
rect 316420 180766 316724 180794
rect 313924 178968 313976 178974
rect 313924 178910 313976 178916
rect 316420 178129 316448 180766
rect 316038 178120 316094 178129
rect 316038 178055 316094 178064
rect 316406 178120 316462 178129
rect 316406 178055 316462 178064
rect 313832 176656 313884 176662
rect 313832 176598 313884 176604
rect 316052 175930 316080 178055
rect 318076 177478 318104 192646
rect 318616 185564 318668 185570
rect 318616 185506 318668 185512
rect 318064 177472 318116 177478
rect 318064 177414 318116 177420
rect 318628 176225 318656 185506
rect 318720 177614 318748 233922
rect 319272 233918 319300 335326
rect 319350 242584 319406 242593
rect 319350 242519 319406 242528
rect 319364 237250 319392 242519
rect 320088 240168 320140 240174
rect 320088 240110 320140 240116
rect 320100 238678 320128 240110
rect 320088 238672 320140 238678
rect 320088 238614 320140 238620
rect 319352 237244 319404 237250
rect 319352 237186 319404 237192
rect 319260 233912 319312 233918
rect 319260 233854 319312 233860
rect 320192 185570 320220 366046
rect 320284 345545 320312 400182
rect 321560 386504 321612 386510
rect 321560 386446 321612 386452
rect 320824 363248 320876 363254
rect 320824 363190 320876 363196
rect 320364 359440 320416 359446
rect 320364 359382 320416 359388
rect 320376 358834 320404 359382
rect 320364 358828 320416 358834
rect 320364 358770 320416 358776
rect 320270 345536 320326 345545
rect 320270 345471 320326 345480
rect 320284 345098 320312 345471
rect 320272 345092 320324 345098
rect 320272 345034 320324 345040
rect 320270 248840 320326 248849
rect 320270 248775 320326 248784
rect 320284 248470 320312 248775
rect 320272 248464 320324 248470
rect 320272 248406 320324 248412
rect 320284 239970 320312 248406
rect 320362 246800 320418 246809
rect 320362 246735 320418 246744
rect 320376 245682 320404 246735
rect 320364 245676 320416 245682
rect 320364 245618 320416 245624
rect 320272 239964 320324 239970
rect 320272 239906 320324 239912
rect 320376 238134 320404 245618
rect 320364 238128 320416 238134
rect 320364 238070 320416 238076
rect 320836 188426 320864 363190
rect 321572 352209 321600 386446
rect 323596 386442 323624 418134
rect 353300 409896 353352 409902
rect 353300 409838 353352 409844
rect 324412 390584 324464 390590
rect 324412 390526 324464 390532
rect 323584 386436 323636 386442
rect 323584 386378 323636 386384
rect 323124 368620 323176 368626
rect 323124 368562 323176 368568
rect 321836 367124 321888 367130
rect 321836 367066 321888 367072
rect 321652 363112 321704 363118
rect 321652 363054 321704 363060
rect 321664 359145 321692 363054
rect 321742 359408 321798 359417
rect 321742 359343 321798 359352
rect 321650 359136 321706 359145
rect 321650 359071 321706 359080
rect 321652 358964 321704 358970
rect 321652 358906 321704 358912
rect 321558 352200 321614 352209
rect 321558 352135 321614 352144
rect 321664 331809 321692 358906
rect 321756 334665 321784 359343
rect 321848 347449 321876 367066
rect 323032 365968 323084 365974
rect 323032 365910 323084 365916
rect 322940 360256 322992 360262
rect 322940 360198 322992 360204
rect 322848 354408 322900 354414
rect 322846 354376 322848 354385
rect 322900 354376 322902 354385
rect 322846 354311 322902 354320
rect 322202 352200 322258 352209
rect 322202 352135 322258 352144
rect 322216 348430 322244 352135
rect 322662 350160 322718 350169
rect 322662 350095 322718 350104
rect 322676 349858 322704 350095
rect 322664 349852 322716 349858
rect 322664 349794 322716 349800
rect 322204 348424 322256 348430
rect 322204 348366 322256 348372
rect 321834 347440 321890 347449
rect 321834 347375 321890 347384
rect 322294 347440 322350 347449
rect 322294 347375 322350 347384
rect 322308 347070 322336 347375
rect 322296 347064 322348 347070
rect 322296 347006 322348 347012
rect 322478 343360 322534 343369
rect 322478 343295 322534 343304
rect 322492 342922 322520 343295
rect 322480 342916 322532 342922
rect 322480 342858 322532 342864
rect 322848 342236 322900 342242
rect 322848 342178 322900 342184
rect 322860 341465 322888 342178
rect 322846 341456 322902 341465
rect 322846 341391 322902 341400
rect 322480 336728 322532 336734
rect 322478 336696 322480 336705
rect 322532 336696 322534 336705
rect 322478 336631 322534 336640
rect 321742 334656 321798 334665
rect 321742 334591 321744 334600
rect 321796 334591 321798 334600
rect 321744 334562 321796 334568
rect 321756 334531 321784 334562
rect 321650 331800 321706 331809
rect 321650 331735 321706 331744
rect 322202 331800 322258 331809
rect 322202 331735 322204 331744
rect 322256 331735 322258 331744
rect 322204 331706 322256 331712
rect 322204 330540 322256 330546
rect 322204 330482 322256 330488
rect 322216 329905 322244 330482
rect 322202 329896 322258 329905
rect 322202 329831 322258 329840
rect 322848 327752 322900 327758
rect 322846 327720 322848 327729
rect 322900 327720 322902 327729
rect 322846 327655 322902 327664
rect 322754 325000 322810 325009
rect 322754 324935 322756 324944
rect 322808 324935 322810 324944
rect 322756 324906 322808 324912
rect 322480 322992 322532 322998
rect 322478 322960 322480 322969
rect 322532 322960 322534 322969
rect 322478 322895 322534 322904
rect 322202 320920 322258 320929
rect 322202 320855 322258 320864
rect 322216 301578 322244 320855
rect 322846 318880 322902 318889
rect 322846 318815 322848 318824
rect 322900 318815 322902 318824
rect 322848 318786 322900 318792
rect 322480 317416 322532 317422
rect 322480 317358 322532 317364
rect 322492 316305 322520 317358
rect 322478 316296 322534 316305
rect 322478 316231 322534 316240
rect 322480 314628 322532 314634
rect 322480 314570 322532 314576
rect 322492 314265 322520 314570
rect 322478 314256 322534 314265
rect 322478 314191 322534 314200
rect 322846 312080 322902 312089
rect 322846 312015 322848 312024
rect 322900 312015 322902 312024
rect 322848 311986 322900 311992
rect 322480 309800 322532 309806
rect 322480 309742 322532 309748
rect 322492 309505 322520 309742
rect 322478 309496 322534 309505
rect 322478 309431 322534 309440
rect 322480 307760 322532 307766
rect 322480 307702 322532 307708
rect 322492 307465 322520 307702
rect 322478 307456 322534 307465
rect 322478 307391 322534 307400
rect 322478 305280 322534 305289
rect 322478 305215 322534 305224
rect 322492 305046 322520 305215
rect 322480 305040 322532 305046
rect 322480 304982 322532 304988
rect 322478 303240 322534 303249
rect 322478 303175 322534 303184
rect 322492 302258 322520 303175
rect 322480 302252 322532 302258
rect 322480 302194 322532 302200
rect 322204 301572 322256 301578
rect 322204 301514 322256 301520
rect 322848 301504 322900 301510
rect 322848 301446 322900 301452
rect 322860 300665 322888 301446
rect 322846 300656 322902 300665
rect 322846 300591 322902 300600
rect 322480 298784 322532 298790
rect 322480 298726 322532 298732
rect 322492 298625 322520 298726
rect 322478 298616 322534 298625
rect 322478 298551 322534 298560
rect 322478 296440 322534 296449
rect 322478 296375 322534 296384
rect 322492 295390 322520 296375
rect 322480 295384 322532 295390
rect 322480 295326 322532 295332
rect 322846 293720 322902 293729
rect 322846 293655 322902 293664
rect 322860 293282 322888 293655
rect 322848 293276 322900 293282
rect 322848 293218 322900 293224
rect 322846 291680 322902 291689
rect 322846 291615 322902 291624
rect 322860 291242 322888 291615
rect 322848 291236 322900 291242
rect 322848 291178 322900 291184
rect 322846 289640 322902 289649
rect 322846 289575 322902 289584
rect 322860 288454 322888 289575
rect 322848 288448 322900 288454
rect 322848 288390 322900 288396
rect 321558 286920 321614 286929
rect 321558 286855 321614 286864
rect 321572 235890 321600 286855
rect 322204 286340 322256 286346
rect 322204 286282 322256 286288
rect 322216 285025 322244 286282
rect 322202 285016 322258 285025
rect 322202 284951 322258 284960
rect 322478 282976 322534 282985
rect 322478 282911 322480 282920
rect 322532 282911 322534 282920
rect 322480 282882 322532 282888
rect 322478 280800 322534 280809
rect 322478 280735 322534 280744
rect 322492 280226 322520 280735
rect 322480 280220 322532 280226
rect 322480 280162 322532 280168
rect 322202 278080 322258 278089
rect 322202 278015 322258 278024
rect 322216 276146 322244 278015
rect 322204 276140 322256 276146
rect 322204 276082 322256 276088
rect 321650 255640 321706 255649
rect 321650 255575 321706 255584
rect 321560 235884 321612 235890
rect 321560 235826 321612 235832
rect 321572 234734 321600 235826
rect 321560 234728 321612 234734
rect 321560 234670 321612 234676
rect 321664 233986 321692 255575
rect 321744 242956 321796 242962
rect 321744 242898 321796 242904
rect 321756 242593 321784 242898
rect 321742 242584 321798 242593
rect 321742 242519 321798 242528
rect 321742 240000 321798 240009
rect 321742 239935 321798 239944
rect 321652 233980 321704 233986
rect 321652 233922 321704 233928
rect 321756 229094 321784 239935
rect 322216 237386 322244 276082
rect 322848 276072 322900 276078
rect 322846 276040 322848 276049
rect 322900 276040 322902 276049
rect 322846 275975 322902 275984
rect 322388 274644 322440 274650
rect 322388 274586 322440 274592
rect 322400 274145 322428 274586
rect 322386 274136 322442 274145
rect 322386 274071 322442 274080
rect 322846 271280 322902 271289
rect 322846 271215 322902 271224
rect 322860 270570 322888 271215
rect 322848 270564 322900 270570
rect 322848 270506 322900 270512
rect 322846 269240 322902 269249
rect 322846 269175 322902 269184
rect 322860 269142 322888 269175
rect 322848 269136 322900 269142
rect 322848 269078 322900 269084
rect 322480 267708 322532 267714
rect 322480 267650 322532 267656
rect 322492 267345 322520 267650
rect 322478 267336 322534 267345
rect 322478 267271 322534 267280
rect 322478 265160 322534 265169
rect 322478 265095 322534 265104
rect 322492 264994 322520 265095
rect 322480 264988 322532 264994
rect 322480 264930 322532 264936
rect 322478 262440 322534 262449
rect 322478 262375 322534 262384
rect 322492 262274 322520 262375
rect 322480 262268 322532 262274
rect 322480 262210 322532 262216
rect 322570 260400 322626 260409
rect 322570 260335 322626 260344
rect 322584 259486 322612 260335
rect 322572 259480 322624 259486
rect 322572 259422 322624 259428
rect 322478 251560 322534 251569
rect 322478 251495 322534 251504
rect 322492 251326 322520 251495
rect 322480 251320 322532 251326
rect 322480 251262 322532 251268
rect 322846 244760 322902 244769
rect 322846 244695 322902 244704
rect 322860 244322 322888 244695
rect 322848 244316 322900 244322
rect 322848 244258 322900 244264
rect 322204 237380 322256 237386
rect 322204 237322 322256 237328
rect 322204 234728 322256 234734
rect 322204 234670 322256 234676
rect 321664 229066 321784 229094
rect 321664 228886 321692 229066
rect 321652 228880 321704 228886
rect 321652 228822 321704 228828
rect 320916 205012 320968 205018
rect 320916 204954 320968 204960
rect 320928 190454 320956 204954
rect 321560 202428 321612 202434
rect 321560 202370 321612 202376
rect 320928 190426 321324 190454
rect 320824 188420 320876 188426
rect 320824 188362 320876 188368
rect 320180 185564 320232 185570
rect 320180 185506 320232 185512
rect 318708 177608 318760 177614
rect 318708 177550 318760 177556
rect 318614 176216 318670 176225
rect 318614 176151 318670 176160
rect 316020 175902 316080 175930
rect 321296 169697 321324 190426
rect 321468 176656 321520 176662
rect 321468 176598 321520 176604
rect 321480 176089 321508 176598
rect 321466 176080 321522 176089
rect 321466 176015 321522 176024
rect 321374 175808 321430 175817
rect 321374 175743 321430 175752
rect 321388 173777 321416 175743
rect 321374 173768 321430 173777
rect 321374 173703 321430 173712
rect 321282 169688 321338 169697
rect 321282 169623 321338 169632
rect 321572 129713 321600 202370
rect 321664 162217 321692 228822
rect 322216 202230 322244 234670
rect 322204 202224 322256 202230
rect 322204 202166 322256 202172
rect 321836 199504 321888 199510
rect 321836 199446 321888 199452
rect 321744 177676 321796 177682
rect 321744 177618 321796 177624
rect 321650 162208 321706 162217
rect 321650 162143 321706 162152
rect 321756 133793 321784 177618
rect 321848 172689 321876 199446
rect 321834 172680 321890 172689
rect 321834 172615 321890 172624
rect 322952 160857 322980 360198
rect 323044 338745 323072 365910
rect 323136 349858 323164 368562
rect 323124 349852 323176 349858
rect 323124 349794 323176 349800
rect 323596 342310 323624 386378
rect 324320 360324 324372 360330
rect 324320 360266 324372 360272
rect 323584 342304 323636 342310
rect 323584 342246 323636 342252
rect 323030 338736 323086 338745
rect 323030 338671 323086 338680
rect 323044 338434 323072 338671
rect 323032 338428 323084 338434
rect 323032 338370 323084 338376
rect 323584 338428 323636 338434
rect 323584 338370 323636 338376
rect 323216 324964 323268 324970
rect 323216 324906 323268 324912
rect 323124 177404 323176 177410
rect 323124 177346 323176 177352
rect 323032 176044 323084 176050
rect 323032 175986 323084 175992
rect 322938 160848 322994 160857
rect 322938 160783 322994 160792
rect 323044 154737 323072 175986
rect 323136 159361 323164 177346
rect 323228 174729 323256 324906
rect 323596 194002 323624 338370
rect 323676 318844 323728 318850
rect 323676 318786 323728 318792
rect 323688 237522 323716 318786
rect 324332 293282 324360 360266
rect 324424 327758 324452 390526
rect 335542 389192 335598 389201
rect 335542 389127 335598 389136
rect 331220 376032 331272 376038
rect 331220 375974 331272 375980
rect 327264 374128 327316 374134
rect 327264 374070 327316 374076
rect 327172 372836 327224 372842
rect 327172 372778 327224 372784
rect 324964 370184 325016 370190
rect 324964 370126 325016 370132
rect 324504 367260 324556 367266
rect 324504 367202 324556 367208
rect 324516 354414 324544 367202
rect 324504 354408 324556 354414
rect 324504 354350 324556 354356
rect 324516 353433 324544 354350
rect 324502 353424 324558 353433
rect 324502 353359 324558 353368
rect 324412 327752 324464 327758
rect 324412 327694 324464 327700
rect 324412 312044 324464 312050
rect 324412 311986 324464 311992
rect 324424 311817 324452 311986
rect 324410 311808 324466 311817
rect 324410 311743 324466 311752
rect 324424 311166 324452 311743
rect 324412 311160 324464 311166
rect 324412 311102 324464 311108
rect 324320 293276 324372 293282
rect 324320 293218 324372 293224
rect 324320 291236 324372 291242
rect 324320 291178 324372 291184
rect 323676 237516 323728 237522
rect 323676 237458 323728 237464
rect 323688 237289 323716 237458
rect 323674 237280 323730 237289
rect 323674 237215 323730 237224
rect 324332 229022 324360 291178
rect 324410 258360 324466 258369
rect 324410 258295 324466 258304
rect 324424 258126 324452 258295
rect 324412 258120 324464 258126
rect 324412 258062 324464 258068
rect 324412 244316 324464 244322
rect 324412 244258 324464 244264
rect 324424 233238 324452 244258
rect 324412 233232 324464 233238
rect 324412 233174 324464 233180
rect 324412 232552 324464 232558
rect 324412 232494 324464 232500
rect 324320 229016 324372 229022
rect 324320 228958 324372 228964
rect 323676 220856 323728 220862
rect 323676 220798 323728 220804
rect 323584 193996 323636 194002
rect 323584 193938 323636 193944
rect 323688 178022 323716 220798
rect 323676 178016 323728 178022
rect 323676 177958 323728 177964
rect 323214 174720 323270 174729
rect 323214 174655 323270 174664
rect 324424 174049 324452 232494
rect 324976 181529 325004 370126
rect 327080 365832 327132 365838
rect 327080 365774 327132 365780
rect 325792 364676 325844 364682
rect 325792 364618 325844 364624
rect 325700 331764 325752 331770
rect 325700 331706 325752 331712
rect 325056 301504 325108 301510
rect 325056 301446 325108 301452
rect 325068 290494 325096 301446
rect 325056 290488 325108 290494
rect 325056 290430 325108 290436
rect 325056 276072 325108 276078
rect 325056 276014 325108 276020
rect 325068 240242 325096 276014
rect 325056 240236 325108 240242
rect 325056 240178 325108 240184
rect 325068 237153 325096 240178
rect 325054 237144 325110 237153
rect 325054 237079 325110 237088
rect 324962 181520 325018 181529
rect 324962 181455 325018 181464
rect 324504 180260 324556 180266
rect 324504 180202 324556 180208
rect 324410 174040 324466 174049
rect 324410 173975 324466 173984
rect 324320 169720 324372 169726
rect 324320 169662 324372 169668
rect 324332 168609 324360 169662
rect 324318 168600 324374 168609
rect 324318 168535 324374 168544
rect 324320 168360 324372 168366
rect 324320 168302 324372 168308
rect 324332 167793 324360 168302
rect 324318 167784 324374 167793
rect 324318 167719 324374 167728
rect 324320 165572 324372 165578
rect 324320 165514 324372 165520
rect 324332 165481 324360 165514
rect 324412 165504 324464 165510
rect 324318 165472 324374 165481
rect 324412 165446 324464 165452
rect 324318 165407 324374 165416
rect 324424 164801 324452 165446
rect 324410 164792 324466 164801
rect 324410 164727 324466 164736
rect 324320 164212 324372 164218
rect 324320 164154 324372 164160
rect 324332 163985 324360 164154
rect 324412 164144 324464 164150
rect 324412 164086 324464 164092
rect 324318 163976 324374 163985
rect 324318 163911 324374 163920
rect 324424 163169 324452 164086
rect 324410 163160 324466 163169
rect 324410 163095 324466 163104
rect 324320 162852 324372 162858
rect 324320 162794 324372 162800
rect 324332 162489 324360 162794
rect 324318 162480 324374 162489
rect 324318 162415 324374 162424
rect 323122 159352 323178 159361
rect 323122 159287 323178 159296
rect 324412 158704 324464 158710
rect 324412 158646 324464 158652
rect 324320 158568 324372 158574
rect 324318 158536 324320 158545
rect 324372 158536 324374 158545
rect 324318 158471 324374 158480
rect 324424 157865 324452 158646
rect 324410 157856 324466 157865
rect 324410 157791 324466 157800
rect 324320 156460 324372 156466
rect 324320 156402 324372 156408
rect 324332 156369 324360 156402
rect 324318 156360 324374 156369
rect 324318 156295 324374 156304
rect 323030 154728 323086 154737
rect 323030 154663 323086 154672
rect 324412 154556 324464 154562
rect 324412 154498 324464 154504
rect 324320 154488 324372 154494
rect 324320 154430 324372 154436
rect 324332 154057 324360 154430
rect 324318 154048 324374 154057
rect 324318 153983 324374 153992
rect 324424 153241 324452 154498
rect 324410 153232 324466 153241
rect 324320 153196 324372 153202
rect 324410 153167 324466 153176
rect 324320 153138 324372 153144
rect 324332 152425 324360 153138
rect 324318 152416 324374 152425
rect 324318 152351 324374 152360
rect 324412 151768 324464 151774
rect 324318 151736 324374 151745
rect 324412 151710 324464 151716
rect 324318 151671 324320 151680
rect 324372 151671 324374 151680
rect 324320 151642 324372 151648
rect 324424 150929 324452 151710
rect 324410 150920 324466 150929
rect 324410 150855 324466 150864
rect 324320 150408 324372 150414
rect 324320 150350 324372 150356
rect 324332 150113 324360 150350
rect 324412 150340 324464 150346
rect 324412 150282 324464 150288
rect 324318 150104 324374 150113
rect 324318 150039 324374 150048
rect 324424 149433 324452 150282
rect 324410 149424 324466 149433
rect 324410 149359 324466 149368
rect 324412 149048 324464 149054
rect 324412 148990 324464 148996
rect 324320 148980 324372 148986
rect 324320 148922 324372 148928
rect 324332 148617 324360 148922
rect 324318 148608 324374 148617
rect 324318 148543 324374 148552
rect 324424 147801 324452 148990
rect 324410 147792 324466 147801
rect 324410 147727 324466 147736
rect 324320 147620 324372 147626
rect 324320 147562 324372 147568
rect 324332 147121 324360 147562
rect 324318 147112 324374 147121
rect 324318 147047 324374 147056
rect 324318 146296 324374 146305
rect 324318 146231 324320 146240
rect 324372 146231 324374 146240
rect 324320 146202 324372 146208
rect 324412 145580 324464 145586
rect 324412 145522 324464 145528
rect 324320 144900 324372 144906
rect 324320 144842 324372 144848
rect 324332 144809 324360 144842
rect 324318 144800 324374 144809
rect 324318 144735 324374 144744
rect 324320 143540 324372 143546
rect 324320 143482 324372 143488
rect 324332 142497 324360 143482
rect 324424 143177 324452 145522
rect 324410 143168 324466 143177
rect 324410 143103 324466 143112
rect 324318 142488 324374 142497
rect 324318 142423 324374 142432
rect 324412 142112 324464 142118
rect 324412 142054 324464 142060
rect 324320 142044 324372 142050
rect 324320 141986 324372 141992
rect 324332 141681 324360 141986
rect 324318 141672 324374 141681
rect 324318 141607 324374 141616
rect 324424 140865 324452 142054
rect 324410 140856 324466 140865
rect 324410 140791 324466 140800
rect 324320 139392 324372 139398
rect 324320 139334 324372 139340
rect 324332 138553 324360 139334
rect 324318 138544 324374 138553
rect 324318 138479 324374 138488
rect 324412 137964 324464 137970
rect 324412 137906 324464 137912
rect 324320 137896 324372 137902
rect 324318 137864 324320 137873
rect 324372 137864 324374 137873
rect 324318 137799 324374 137808
rect 324424 137057 324452 137906
rect 324410 137048 324466 137057
rect 324410 136983 324466 136992
rect 324412 136604 324464 136610
rect 324412 136546 324464 136552
rect 324320 136536 324372 136542
rect 324320 136478 324372 136484
rect 324332 136377 324360 136478
rect 324318 136368 324374 136377
rect 324318 136303 324374 136312
rect 324424 135561 324452 136546
rect 324410 135552 324466 135561
rect 324410 135487 324466 135496
rect 323490 134192 323546 134201
rect 323490 134127 323546 134136
rect 323504 133929 323532 134127
rect 323490 133920 323546 133929
rect 323490 133855 323546 133864
rect 321742 133784 321798 133793
rect 321742 133719 321798 133728
rect 324412 131096 324464 131102
rect 324412 131038 324464 131044
rect 324320 131028 324372 131034
rect 324320 130970 324372 130976
rect 324332 130937 324360 130970
rect 324318 130928 324374 130937
rect 324318 130863 324374 130872
rect 324424 130121 324452 131038
rect 324410 130112 324466 130121
rect 324410 130047 324466 130056
rect 324320 129736 324372 129742
rect 321558 129704 321614 129713
rect 324320 129678 324372 129684
rect 321558 129639 321614 129648
rect 324332 128625 324360 129678
rect 324318 128616 324374 128625
rect 324318 128551 324374 128560
rect 324320 128308 324372 128314
rect 324320 128250 324372 128256
rect 324332 127809 324360 128250
rect 324412 128240 324464 128246
rect 324412 128182 324464 128188
rect 324318 127800 324374 127809
rect 324318 127735 324374 127744
rect 324424 127129 324452 128182
rect 324410 127120 324466 127129
rect 324410 127055 324466 127064
rect 324516 126313 324544 180202
rect 324594 176216 324650 176225
rect 324594 176151 324650 176160
rect 324608 170921 324636 176151
rect 324964 171148 325016 171154
rect 324964 171090 325016 171096
rect 324594 170912 324650 170921
rect 324594 170847 324650 170856
rect 324596 149728 324648 149734
rect 324596 149670 324648 149676
rect 324608 145489 324636 149670
rect 324594 145480 324650 145489
rect 324594 145415 324650 145424
rect 324502 126304 324558 126313
rect 324502 126239 324558 126248
rect 324412 125588 324464 125594
rect 324412 125530 324464 125536
rect 324320 125520 324372 125526
rect 324318 125488 324320 125497
rect 324372 125488 324374 125497
rect 324318 125423 324374 125432
rect 324424 124817 324452 125530
rect 324410 124808 324466 124817
rect 324410 124743 324466 124752
rect 324412 124160 324464 124166
rect 324412 124102 324464 124108
rect 324320 124092 324372 124098
rect 324320 124034 324372 124040
rect 324332 124001 324360 124034
rect 324318 123992 324374 124001
rect 324318 123927 324374 123936
rect 324424 123185 324452 124102
rect 324410 123176 324466 123185
rect 324410 123111 324466 123120
rect 324320 122800 324372 122806
rect 324320 122742 324372 122748
rect 324332 122505 324360 122742
rect 324412 122732 324464 122738
rect 324412 122674 324464 122680
rect 324318 122496 324374 122505
rect 324318 122431 324374 122440
rect 324424 121689 324452 122674
rect 324410 121680 324466 121689
rect 324410 121615 324466 121624
rect 324320 121440 324372 121446
rect 324320 121382 324372 121388
rect 324332 120193 324360 121382
rect 324976 120873 325004 171090
rect 325606 160168 325662 160177
rect 325712 160154 325740 331706
rect 325804 330546 325832 364618
rect 325792 330540 325844 330546
rect 325792 330482 325844 330488
rect 327092 309806 327120 365774
rect 327184 336734 327212 372778
rect 327276 342922 327304 374070
rect 329840 358896 329892 358902
rect 329840 358838 329892 358844
rect 327264 342916 327316 342922
rect 327264 342858 327316 342864
rect 327172 336728 327224 336734
rect 327172 336670 327224 336676
rect 328368 336728 328420 336734
rect 328368 336670 328420 336676
rect 328380 336054 328408 336670
rect 328368 336048 328420 336054
rect 328368 335990 328420 335996
rect 328460 334620 328512 334626
rect 328460 334562 328512 334568
rect 327080 309800 327132 309806
rect 327080 309742 327132 309748
rect 327172 305040 327224 305046
rect 327172 304982 327224 304988
rect 327080 302252 327132 302258
rect 327080 302194 327132 302200
rect 326344 269136 326396 269142
rect 326344 269078 326396 269084
rect 325792 251320 325844 251326
rect 325792 251262 325844 251268
rect 325804 248414 325832 251262
rect 325804 248386 325924 248414
rect 325896 233170 325924 248386
rect 326356 235686 326384 269078
rect 327092 240038 327120 302194
rect 327080 240032 327132 240038
rect 327078 240000 327080 240009
rect 327132 240000 327134 240009
rect 327078 239935 327134 239944
rect 326988 236020 327040 236026
rect 326988 235962 327040 235968
rect 327000 235686 327028 235962
rect 326344 235680 326396 235686
rect 326344 235622 326396 235628
rect 326988 235680 327040 235686
rect 326988 235622 327040 235628
rect 325884 233164 325936 233170
rect 325884 233106 325936 233112
rect 327184 230382 327212 304982
rect 327264 288448 327316 288454
rect 327264 288390 327316 288396
rect 327276 234297 327304 288390
rect 327356 259480 327408 259486
rect 327356 259422 327408 259428
rect 327262 234288 327318 234297
rect 327262 234223 327318 234232
rect 327172 230376 327224 230382
rect 327172 230318 327224 230324
rect 327368 229090 327396 259422
rect 327446 234288 327502 234297
rect 327446 234223 327502 234232
rect 327356 229084 327408 229090
rect 327356 229026 327408 229032
rect 327368 228478 327396 229026
rect 327356 228472 327408 228478
rect 327356 228414 327408 228420
rect 325884 216028 325936 216034
rect 325884 215970 325936 215976
rect 325792 192636 325844 192642
rect 325792 192578 325844 192584
rect 325662 160126 325740 160154
rect 325606 160103 325662 160112
rect 324962 120864 325018 120873
rect 324962 120799 325018 120808
rect 324318 120184 324374 120193
rect 324318 120119 324374 120128
rect 324320 120012 324372 120018
rect 324320 119954 324372 119960
rect 324332 119377 324360 119954
rect 324318 119368 324374 119377
rect 324318 119303 324374 119312
rect 324412 118652 324464 118658
rect 324412 118594 324464 118600
rect 324320 118584 324372 118590
rect 324318 118552 324320 118561
rect 324372 118552 324374 118561
rect 324318 118487 324374 118496
rect 324424 117881 324452 118594
rect 324410 117872 324466 117881
rect 324410 117807 324466 117816
rect 324412 117224 324464 117230
rect 324412 117166 324464 117172
rect 324320 117156 324372 117162
rect 324320 117098 324372 117104
rect 324332 117065 324360 117098
rect 324318 117056 324374 117065
rect 324318 116991 324374 117000
rect 324424 116385 324452 117166
rect 324410 116376 324466 116385
rect 324410 116311 324466 116320
rect 324412 115932 324464 115938
rect 324412 115874 324464 115880
rect 324320 115864 324372 115870
rect 324320 115806 324372 115812
rect 324332 115569 324360 115806
rect 324318 115560 324374 115569
rect 324318 115495 324374 115504
rect 324424 114753 324452 115874
rect 324410 114744 324466 114753
rect 324410 114679 324466 114688
rect 324412 114504 324464 114510
rect 324412 114446 324464 114452
rect 324320 114436 324372 114442
rect 324320 114378 324372 114384
rect 324332 114073 324360 114378
rect 324318 114064 324374 114073
rect 324318 113999 324374 114008
rect 324424 113257 324452 114446
rect 324410 113248 324466 113257
rect 324410 113183 324466 113192
rect 324320 113144 324372 113150
rect 324320 113086 324372 113092
rect 324332 112441 324360 113086
rect 324318 112432 324374 112441
rect 324318 112367 324374 112376
rect 324320 111784 324372 111790
rect 324318 111752 324320 111761
rect 324372 111752 324374 111761
rect 324318 111687 324374 111696
rect 324412 111716 324464 111722
rect 324412 111658 324464 111664
rect 324424 110945 324452 111658
rect 324410 110936 324466 110945
rect 324410 110871 324466 110880
rect 324320 110424 324372 110430
rect 324320 110366 324372 110372
rect 324332 109449 324360 110366
rect 324502 110120 324558 110129
rect 324502 110055 324558 110064
rect 324412 109744 324464 109750
rect 324412 109686 324464 109692
rect 324318 109440 324374 109449
rect 324318 109375 324374 109384
rect 324320 108248 324372 108254
rect 324320 108190 324372 108196
rect 324332 107817 324360 108190
rect 324318 107808 324374 107817
rect 324318 107743 324374 107752
rect 324320 107636 324372 107642
rect 324320 107578 324372 107584
rect 324332 107137 324360 107578
rect 324318 107128 324374 107137
rect 324318 107063 324374 107072
rect 322938 106312 322994 106321
rect 322938 106247 322994 106256
rect 321834 105088 321890 105097
rect 321834 105023 321890 105032
rect 321650 102776 321706 102785
rect 321650 102711 321706 102720
rect 321558 99648 321614 99657
rect 321558 99583 321614 99592
rect 321572 96626 321600 99583
rect 321560 96620 321612 96626
rect 321560 96562 321612 96568
rect 309784 96552 309836 96558
rect 309784 96494 309836 96500
rect 321664 96490 321692 102711
rect 321742 102232 321798 102241
rect 321742 102167 321798 102176
rect 321652 96484 321704 96490
rect 321652 96426 321704 96432
rect 321466 95840 321522 95849
rect 321466 95775 321522 95784
rect 321480 95198 321508 95775
rect 321468 95192 321520 95198
rect 321468 95134 321520 95140
rect 321756 95062 321784 102167
rect 321848 95130 321876 105023
rect 322952 96558 322980 106247
rect 324424 104825 324452 109686
rect 324410 104816 324466 104825
rect 324410 104751 324466 104760
rect 324516 103514 324544 110055
rect 324594 108624 324650 108633
rect 324594 108559 324650 108568
rect 324424 103486 324544 103514
rect 323584 102808 323636 102814
rect 323584 102750 323636 102756
rect 322940 96552 322992 96558
rect 322940 96494 322992 96500
rect 321836 95124 321888 95130
rect 321836 95066 321888 95072
rect 321744 95056 321796 95062
rect 321744 94998 321796 95004
rect 323596 93838 323624 102750
rect 324320 102128 324372 102134
rect 324320 102070 324372 102076
rect 324332 101697 324360 102070
rect 324318 101688 324374 101697
rect 324318 101623 324374 101632
rect 324318 99376 324374 99385
rect 324318 99311 324320 99320
rect 324372 99311 324374 99320
rect 324320 99282 324372 99288
rect 324424 98802 324452 103486
rect 324502 100872 324558 100881
rect 324502 100807 324558 100816
rect 324412 98796 324464 98802
rect 324412 98738 324464 98744
rect 324412 98660 324464 98666
rect 324412 98602 324464 98608
rect 324320 97980 324372 97986
rect 324320 97922 324372 97928
rect 324332 97073 324360 97922
rect 324424 97889 324452 98602
rect 324410 97880 324466 97889
rect 324410 97815 324466 97824
rect 324318 97064 324374 97073
rect 324318 96999 324374 97008
rect 324516 94926 324544 100807
rect 324504 94920 324556 94926
rect 324504 94862 324556 94868
rect 324320 94512 324372 94518
rect 324320 94454 324372 94460
rect 323584 93832 323636 93838
rect 323584 93774 323636 93780
rect 320824 93220 320876 93226
rect 320824 93162 320876 93168
rect 311900 89072 311952 89078
rect 311900 89014 311952 89020
rect 309784 79348 309836 79354
rect 309784 79290 309836 79296
rect 309140 73840 309192 73846
rect 309140 73782 309192 73788
rect 308494 40624 308550 40633
rect 308494 40559 308550 40568
rect 307760 27600 307812 27606
rect 307760 27542 307812 27548
rect 308404 27600 308456 27606
rect 308404 27542 308456 27548
rect 307208 4140 307260 4146
rect 307208 4082 307260 4088
rect 307772 3534 307800 27542
rect 308508 6730 308536 40559
rect 309140 40112 309192 40118
rect 309140 40054 309192 40060
rect 309152 6914 309180 40054
rect 309796 16574 309824 79290
rect 311164 73840 311216 73846
rect 311164 73782 311216 73788
rect 311176 49706 311204 73782
rect 310520 49700 310572 49706
rect 310520 49642 310572 49648
rect 311164 49700 311216 49706
rect 311164 49642 311216 49648
rect 310532 16574 310560 49642
rect 311912 16574 311940 89014
rect 316040 84856 316092 84862
rect 316040 84798 316092 84804
rect 316052 81433 316080 84798
rect 316038 81424 316094 81433
rect 316038 81359 316094 81368
rect 313924 80708 313976 80714
rect 313924 80650 313976 80656
rect 313936 42770 313964 80650
rect 315304 47728 315356 47734
rect 315304 47670 315356 47676
rect 313280 42764 313332 42770
rect 313280 42706 313332 42712
rect 313924 42764 313976 42770
rect 313924 42706 313976 42712
rect 313292 16574 313320 42706
rect 309796 16546 309916 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 313292 16546 313872 16574
rect 309152 6886 309824 6914
rect 308496 6724 308548 6730
rect 308496 6666 308548 6672
rect 307760 3528 307812 3534
rect 307760 3470 307812 3476
rect 301934 354 302046 480
rect 301792 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 354 308026 480
rect 308508 354 308536 6666
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309060 480 309088 3470
rect 307914 326 308536 354
rect 307914 -960 308026 326
rect 309018 -960 309130 480
rect 309796 354 309824 6886
rect 309888 6730 309916 16546
rect 309876 6724 309928 6730
rect 309876 6666 309928 6672
rect 311452 480 311480 16546
rect 310214 354 310326 480
rect 309796 326 310326 354
rect 310214 -960 310326 326
rect 311410 -960 311522 480
rect 312188 354 312216 16546
rect 313844 480 313872 16546
rect 315316 13802 315344 47670
rect 314660 13796 314712 13802
rect 314660 13738 314712 13744
rect 315304 13796 315356 13802
rect 315304 13738 315356 13744
rect 312606 354 312718 480
rect 312188 326 312718 354
rect 312606 -960 312718 326
rect 313802 -960 313914 480
rect 314672 354 314700 13738
rect 316052 3482 316080 81359
rect 317420 80096 317472 80102
rect 317420 80038 317472 80044
rect 316130 43480 316186 43489
rect 316130 43415 316186 43424
rect 317326 43480 317382 43489
rect 317326 43415 317328 43424
rect 316144 3602 316172 43415
rect 317380 43415 317382 43424
rect 317328 43386 317380 43392
rect 317432 16574 317460 80038
rect 320836 73166 320864 93162
rect 323596 93090 323624 93774
rect 322940 93084 322992 93090
rect 322940 93026 322992 93032
rect 323584 93084 323636 93090
rect 323584 93026 323636 93032
rect 321560 90364 321612 90370
rect 321560 90306 321612 90312
rect 320824 73160 320876 73166
rect 320824 73102 320876 73108
rect 320836 71806 320864 73102
rect 320180 71800 320232 71806
rect 320180 71742 320232 71748
rect 320824 71800 320876 71806
rect 320824 71742 320876 71748
rect 320192 16574 320220 71742
rect 321572 16574 321600 90306
rect 317432 16546 318104 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 316132 3596 316184 3602
rect 316132 3538 316184 3544
rect 317328 3596 317380 3602
rect 317328 3538 317380 3544
rect 316052 3454 316264 3482
rect 316236 480 316264 3454
rect 317340 480 317368 3538
rect 314998 354 315110 480
rect 314672 326 315110 354
rect 314998 -960 315110 326
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 16546
rect 319720 8968 319772 8974
rect 319720 8910 319772 8916
rect 319732 480 319760 8910
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320468 354 320496 16546
rect 322124 480 322152 16546
rect 320886 354 320998 480
rect 320468 326 320998 354
rect 320886 -960 320998 326
rect 322082 -960 322194 480
rect 322952 354 322980 93026
rect 324332 16574 324360 94454
rect 324608 93770 324636 108559
rect 325606 104272 325662 104281
rect 325804 104258 325832 192578
rect 325896 132433 325924 215970
rect 327264 200932 327316 200938
rect 327264 200874 327316 200880
rect 325976 179036 326028 179042
rect 325976 178978 326028 178984
rect 325882 132424 325938 132433
rect 325882 132359 325938 132368
rect 325988 120018 326016 178978
rect 327172 178832 327224 178838
rect 327172 178774 327224 178780
rect 327080 178016 327132 178022
rect 327080 177958 327132 177964
rect 327092 171154 327120 177958
rect 327080 171148 327132 171154
rect 327080 171090 327132 171096
rect 325976 120012 326028 120018
rect 325976 119954 326028 119960
rect 327184 108254 327212 178774
rect 327276 156466 327304 200874
rect 327460 158574 327488 234223
rect 328368 230376 328420 230382
rect 328368 230318 328420 230324
rect 328380 229838 328408 230318
rect 328368 229832 328420 229838
rect 328368 229774 328420 229780
rect 327448 158568 327500 158574
rect 327448 158510 327500 158516
rect 327264 156460 327316 156466
rect 327264 156402 327316 156408
rect 327724 155236 327776 155242
rect 327724 155178 327776 155184
rect 327736 125526 327764 155178
rect 327724 125520 327776 125526
rect 327724 125462 327776 125468
rect 328472 109750 328500 334562
rect 328552 330540 328604 330546
rect 328552 330482 328604 330488
rect 328564 143546 328592 330482
rect 329852 324970 329880 358838
rect 329840 324964 329892 324970
rect 329840 324906 329892 324912
rect 329840 322992 329892 322998
rect 329840 322934 329892 322940
rect 329852 240145 329880 322934
rect 331232 307766 331260 375974
rect 333980 368756 334032 368762
rect 333980 368698 334032 368704
rect 333992 314634 334020 368698
rect 335452 368688 335504 368694
rect 335452 368630 335504 368636
rect 335360 364608 335412 364614
rect 335360 364550 335412 364556
rect 334624 348424 334676 348430
rect 334624 348366 334676 348372
rect 334636 324970 334664 348366
rect 334624 324964 334676 324970
rect 334624 324906 334676 324912
rect 333980 314628 334032 314634
rect 333980 314570 334032 314576
rect 333992 313954 334020 314570
rect 333980 313948 334032 313954
rect 333980 313890 334032 313896
rect 331220 307760 331272 307766
rect 331220 307702 331272 307708
rect 331232 307086 331260 307702
rect 331220 307080 331272 307086
rect 331220 307022 331272 307028
rect 333980 301572 334032 301578
rect 333980 301514 334032 301520
rect 333992 300898 334020 301514
rect 333980 300892 334032 300898
rect 333980 300834 334032 300840
rect 330484 298784 330536 298790
rect 330484 298726 330536 298732
rect 330496 297430 330524 298726
rect 330484 297424 330536 297430
rect 330484 297366 330536 297372
rect 331220 295384 331272 295390
rect 331220 295326 331272 295332
rect 329932 282940 329984 282946
rect 329932 282882 329984 282888
rect 329838 240136 329894 240145
rect 329838 240071 329840 240080
rect 329892 240071 329894 240080
rect 329840 240042 329892 240048
rect 329852 240011 329880 240042
rect 329944 231674 329972 282882
rect 330024 264988 330076 264994
rect 330024 264930 330076 264936
rect 329932 231668 329984 231674
rect 329932 231610 329984 231616
rect 329944 219434 329972 231610
rect 330036 227526 330064 264930
rect 330024 227520 330076 227526
rect 330024 227462 330076 227468
rect 329852 219406 329972 219434
rect 328644 202224 328696 202230
rect 328644 202166 328696 202172
rect 328656 148986 328684 202166
rect 328736 196784 328788 196790
rect 328736 196726 328788 196732
rect 328748 154494 328776 196726
rect 328736 154488 328788 154494
rect 328736 154430 328788 154436
rect 328644 148980 328696 148986
rect 328644 148922 328696 148928
rect 328552 143540 328604 143546
rect 328552 143482 328604 143488
rect 329852 142050 329880 219406
rect 329932 207868 329984 207874
rect 329932 207810 329984 207816
rect 329840 142044 329892 142050
rect 329840 141986 329892 141992
rect 329944 128246 329972 207810
rect 330036 153202 330064 227462
rect 331232 226273 331260 295326
rect 331312 270564 331364 270570
rect 331312 270506 331364 270512
rect 331324 233102 331352 270506
rect 332600 263560 332652 263566
rect 332600 263502 332652 263508
rect 332612 262274 332640 263502
rect 332600 262268 332652 262274
rect 332600 262210 332652 262216
rect 332612 237318 332640 262210
rect 332968 237516 333020 237522
rect 332968 237458 333020 237464
rect 332600 237312 332652 237318
rect 332600 237254 332652 237260
rect 331312 233096 331364 233102
rect 331312 233038 331364 233044
rect 331218 226264 331274 226273
rect 331218 226199 331274 226208
rect 330116 193928 330168 193934
rect 330116 193870 330168 193876
rect 330024 153196 330076 153202
rect 330024 153138 330076 153144
rect 330128 151706 330156 193870
rect 330116 151700 330168 151706
rect 330116 151642 330168 151648
rect 329932 128240 329984 128246
rect 329932 128182 329984 128188
rect 328460 109744 328512 109750
rect 328460 109686 328512 109692
rect 327172 108248 327224 108254
rect 327172 108190 327224 108196
rect 325662 104230 325832 104258
rect 325606 104207 325662 104216
rect 325700 104168 325752 104174
rect 325700 104110 325752 104116
rect 324688 98796 324740 98802
rect 324688 98738 324740 98744
rect 324700 94994 324728 98738
rect 324688 94988 324740 94994
rect 324688 94930 324740 94936
rect 324596 93764 324648 93770
rect 324596 93706 324648 93712
rect 324964 82136 325016 82142
rect 324964 82078 325016 82084
rect 324332 16546 324452 16574
rect 324424 480 324452 16546
rect 324976 9654 325004 82078
rect 325712 16574 325740 104110
rect 330484 100020 330536 100026
rect 330484 99962 330536 99968
rect 327724 46232 327776 46238
rect 327724 46174 327776 46180
rect 327736 33114 327764 46174
rect 327724 33108 327776 33114
rect 327724 33050 327776 33056
rect 327736 31822 327764 33050
rect 327080 31816 327132 31822
rect 327080 31758 327132 31764
rect 327724 31816 327776 31822
rect 327724 31758 327776 31764
rect 327092 16574 327120 31758
rect 330496 26217 330524 99962
rect 331232 98666 331260 226199
rect 331324 131034 331352 233038
rect 331496 182844 331548 182850
rect 331496 182786 331548 182792
rect 331404 177608 331456 177614
rect 331404 177550 331456 177556
rect 331416 150346 331444 177550
rect 331508 164150 331536 182786
rect 332876 180328 332928 180334
rect 332876 180270 332928 180276
rect 332692 178968 332744 178974
rect 332692 178910 332744 178916
rect 331496 164144 331548 164150
rect 331496 164086 331548 164092
rect 332048 154624 332100 154630
rect 332048 154566 332100 154572
rect 331404 150340 331456 150346
rect 331404 150282 331456 150288
rect 331862 147792 331918 147801
rect 331862 147727 331918 147736
rect 331312 131028 331364 131034
rect 331312 130970 331364 130976
rect 331220 98660 331272 98666
rect 331220 98602 331272 98608
rect 330482 26208 330538 26217
rect 330482 26143 330538 26152
rect 330496 24993 330524 26143
rect 329838 24984 329894 24993
rect 329838 24919 329894 24928
rect 330482 24984 330538 24993
rect 330482 24919 330538 24928
rect 329104 21412 329156 21418
rect 329104 21354 329156 21360
rect 329116 16574 329144 21354
rect 329852 16574 329880 24919
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 329116 16546 329236 16574
rect 329852 16546 330432 16574
rect 324964 9648 325016 9654
rect 324964 9590 325016 9596
rect 325608 9648 325660 9654
rect 325608 9590 325660 9596
rect 325620 480 325648 9590
rect 323278 354 323390 480
rect 322952 326 323390 354
rect 323278 -960 323390 326
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 354 326384 16546
rect 328012 480 328040 16546
rect 329208 480 329236 16546
rect 330404 480 330432 16546
rect 331876 10402 331904 147727
rect 332060 84182 332088 154566
rect 332506 147792 332562 147801
rect 332506 147727 332562 147736
rect 332520 147694 332548 147727
rect 332508 147688 332560 147694
rect 332508 147630 332560 147636
rect 332704 115870 332732 178910
rect 332784 177472 332836 177478
rect 332784 177414 332836 177420
rect 332796 154562 332824 177414
rect 332888 165510 332916 180270
rect 332876 165504 332928 165510
rect 332876 165446 332928 165452
rect 332784 154556 332836 154562
rect 332784 154498 332836 154504
rect 332692 115864 332744 115870
rect 332692 115806 332744 115812
rect 332980 102134 333008 237458
rect 333992 234433 334020 300834
rect 335268 300144 335320 300150
rect 335268 300086 335320 300092
rect 335280 263634 335308 300086
rect 335268 263628 335320 263634
rect 335268 263570 335320 263576
rect 333978 234424 334034 234433
rect 333978 234359 334034 234368
rect 333980 233164 334032 233170
rect 333980 233106 334032 233112
rect 333992 155242 334020 233106
rect 334716 229764 334768 229770
rect 334716 229706 334768 229712
rect 334072 188420 334124 188426
rect 334072 188362 334124 188368
rect 334084 162858 334112 188362
rect 334164 181620 334216 181626
rect 334164 181562 334216 181568
rect 334176 164218 334204 181562
rect 334164 164212 334216 164218
rect 334164 164154 334216 164160
rect 334072 162852 334124 162858
rect 334072 162794 334124 162800
rect 333980 155236 334032 155242
rect 333980 155178 334032 155184
rect 333244 142180 333296 142186
rect 333244 142122 333296 142128
rect 332968 102128 333020 102134
rect 332968 102070 333020 102076
rect 333256 84862 333284 142122
rect 334624 141432 334676 141438
rect 334624 141374 334676 141380
rect 333244 84856 333296 84862
rect 333244 84798 333296 84804
rect 332048 84176 332100 84182
rect 332048 84118 332100 84124
rect 331956 83496 332008 83502
rect 331956 83438 332008 83444
rect 331968 21418 331996 83438
rect 332048 65680 332100 65686
rect 332048 65622 332100 65628
rect 331956 21412 332008 21418
rect 331956 21354 332008 21360
rect 331864 10396 331916 10402
rect 331864 10338 331916 10344
rect 332060 9586 332088 65622
rect 333244 64320 333296 64326
rect 333244 64262 333296 64268
rect 332598 59936 332654 59945
rect 332598 59871 332654 59880
rect 332612 59362 332640 59871
rect 332600 59356 332652 59362
rect 332600 59298 332652 59304
rect 332048 9580 332100 9586
rect 332048 9522 332100 9528
rect 332060 9314 332088 9522
rect 331588 9308 331640 9314
rect 331588 9250 331640 9256
rect 332048 9308 332100 9314
rect 332048 9250 332100 9256
rect 331600 480 331628 9250
rect 332612 3534 332640 59298
rect 333256 4146 333284 64262
rect 333978 44840 334034 44849
rect 333978 44775 334034 44784
rect 333992 6914 334020 44775
rect 334636 8974 334664 141374
rect 334728 135250 334756 229706
rect 334808 161492 334860 161498
rect 334808 161434 334860 161440
rect 334716 135244 334768 135250
rect 334716 135186 334768 135192
rect 334820 76673 334848 161434
rect 335372 121446 335400 364550
rect 335464 158710 335492 368630
rect 335556 317422 335584 389127
rect 349804 382968 349856 382974
rect 349804 382910 349856 382916
rect 346400 378208 346452 378214
rect 346400 378150 346452 378156
rect 339500 375420 339552 375426
rect 339500 375362 339552 375368
rect 338764 371272 338816 371278
rect 338764 371214 338816 371220
rect 337384 370524 337436 370530
rect 337384 370466 337436 370472
rect 335544 317416 335596 317422
rect 335544 317358 335596 317364
rect 336648 317416 336700 317422
rect 336648 317358 336700 317364
rect 336660 316742 336688 317358
rect 336648 316736 336700 316742
rect 336648 316678 336700 316684
rect 336004 280220 336056 280226
rect 336004 280162 336056 280168
rect 336016 271930 336044 280162
rect 336004 271924 336056 271930
rect 336004 271866 336056 271872
rect 336016 227662 336044 271866
rect 336004 227656 336056 227662
rect 336004 227598 336056 227604
rect 336924 195492 336976 195498
rect 336924 195434 336976 195440
rect 335636 189984 335688 189990
rect 335636 189926 335688 189932
rect 335544 187196 335596 187202
rect 335544 187138 335596 187144
rect 335452 158704 335504 158710
rect 335452 158646 335504 158652
rect 335556 149054 335584 187138
rect 335648 169726 335676 189926
rect 336740 181756 336792 181762
rect 336740 181698 336792 181704
rect 335636 169720 335688 169726
rect 335636 169662 335688 169668
rect 336004 155984 336056 155990
rect 336004 155926 336056 155932
rect 335544 149048 335596 149054
rect 335544 148990 335596 148996
rect 335360 121440 335412 121446
rect 335360 121382 335412 121388
rect 334806 76664 334862 76673
rect 334806 76599 334862 76608
rect 335360 69012 335412 69018
rect 335360 68954 335412 68960
rect 335372 16574 335400 68954
rect 336016 39642 336044 155926
rect 336752 111722 336780 181698
rect 336832 178900 336884 178906
rect 336832 178842 336884 178848
rect 336844 111790 336872 178842
rect 336936 137902 336964 195434
rect 336924 137896 336976 137902
rect 336924 137838 336976 137844
rect 336832 111784 336884 111790
rect 336832 111726 336884 111732
rect 336740 111716 336792 111722
rect 336740 111658 336792 111664
rect 336096 84856 336148 84862
rect 336096 84798 336148 84804
rect 336108 69018 336136 84798
rect 336096 69012 336148 69018
rect 336096 68954 336148 68960
rect 336004 39636 336056 39642
rect 336004 39578 336056 39584
rect 337396 16574 337424 370466
rect 338120 209228 338172 209234
rect 338120 209170 338172 209176
rect 338132 117230 338160 209170
rect 338304 182912 338356 182918
rect 338304 182854 338356 182860
rect 338212 177336 338264 177342
rect 338212 177278 338264 177284
rect 338224 136542 338252 177278
rect 338316 145586 338344 182854
rect 338776 167686 338804 371214
rect 338764 167680 338816 167686
rect 338764 167622 338816 167628
rect 338764 165640 338816 165646
rect 338764 165582 338816 165588
rect 338304 145580 338356 145586
rect 338304 145522 338356 145528
rect 338212 136536 338264 136542
rect 338212 136478 338264 136484
rect 338120 117224 338172 117230
rect 338120 117166 338172 117172
rect 338776 78674 338804 165582
rect 339512 99346 339540 375362
rect 339592 371884 339644 371890
rect 339592 371826 339644 371832
rect 339604 274650 339632 371826
rect 342260 371340 342312 371346
rect 342260 371282 342312 371288
rect 340880 367464 340932 367470
rect 340880 367406 340932 367412
rect 339592 274644 339644 274650
rect 339592 274586 339644 274592
rect 339604 273970 339632 274586
rect 339592 273964 339644 273970
rect 339592 273906 339644 273912
rect 340236 227044 340288 227050
rect 340236 226986 340288 226992
rect 339592 188488 339644 188494
rect 339592 188430 339644 188436
rect 339604 137970 339632 188430
rect 339684 178696 339736 178702
rect 339684 178638 339736 178644
rect 339696 165578 339724 178638
rect 339684 165572 339736 165578
rect 339684 165514 339736 165520
rect 340144 162920 340196 162926
rect 340144 162862 340196 162868
rect 339592 137964 339644 137970
rect 339592 137906 339644 137912
rect 339500 99340 339552 99346
rect 339500 99282 339552 99288
rect 338764 78668 338816 78674
rect 338764 78610 338816 78616
rect 339132 78668 339184 78674
rect 339132 78610 339184 78616
rect 339144 77897 339172 78610
rect 339130 77888 339186 77897
rect 339130 77823 339186 77832
rect 339500 69692 339552 69698
rect 339500 69634 339552 69640
rect 338120 46232 338172 46238
rect 338120 46174 338172 46180
rect 335372 16546 336320 16574
rect 334624 8968 334676 8974
rect 334624 8910 334676 8916
rect 333992 6886 334664 6914
rect 332692 4140 332744 4146
rect 332692 4082 332744 4088
rect 333244 4140 333296 4146
rect 333244 4082 333296 4088
rect 332600 3528 332652 3534
rect 332600 3470 332652 3476
rect 332704 480 332732 4082
rect 333888 3528 333940 3534
rect 333888 3470 333940 3476
rect 333900 480 333928 3470
rect 326774 354 326886 480
rect 326356 326 326886 354
rect 326774 -960 326886 326
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 354 334664 6886
rect 336292 480 336320 16546
rect 337028 16546 337424 16574
rect 338132 16574 338160 46174
rect 338132 16546 338712 16574
rect 337028 15162 337056 16546
rect 337016 15156 337068 15162
rect 337016 15098 337068 15104
rect 335054 354 335166 480
rect 334636 326 335166 354
rect 335054 -960 335166 326
rect 336250 -960 336362 480
rect 337028 354 337056 15098
rect 338684 480 338712 16546
rect 337446 354 337558 480
rect 337028 326 337558 354
rect 337446 -960 337558 326
rect 338642 -960 338754 480
rect 339512 354 339540 69634
rect 340156 48278 340184 162862
rect 340248 117298 340276 226986
rect 340892 147626 340920 367406
rect 342272 267714 342300 371282
rect 343640 368824 343692 368830
rect 343640 368766 343692 368772
rect 342260 267708 342312 267714
rect 342260 267650 342312 267656
rect 342272 267034 342300 267650
rect 342260 267028 342312 267034
rect 342260 266970 342312 266976
rect 340972 229832 341024 229838
rect 340972 229774 341024 229780
rect 340880 147620 340932 147626
rect 340880 147562 340932 147568
rect 340236 117292 340288 117298
rect 340236 117234 340288 117240
rect 340984 117162 341012 229774
rect 342260 225684 342312 225690
rect 342260 225626 342312 225632
rect 341064 193996 341116 194002
rect 341064 193938 341116 193944
rect 340972 117156 341024 117162
rect 340972 117098 341024 117104
rect 341076 110430 341104 193938
rect 341156 181688 341208 181694
rect 341156 181630 341208 181636
rect 341168 114442 341196 181630
rect 342272 122738 342300 225626
rect 342904 211948 342956 211954
rect 342904 211890 342956 211896
rect 342352 186992 342404 186998
rect 342352 186934 342404 186940
rect 342260 122732 342312 122738
rect 342260 122674 342312 122680
rect 342364 118590 342392 186934
rect 342352 118584 342404 118590
rect 342352 118526 342404 118532
rect 341156 114436 341208 114442
rect 341156 114378 341208 114384
rect 341064 110424 341116 110430
rect 341064 110366 341116 110372
rect 342916 106282 342944 211890
rect 342996 176724 343048 176730
rect 342996 176666 343048 176672
rect 342904 106276 342956 106282
rect 342904 106218 342956 106224
rect 342260 86420 342312 86426
rect 342260 86362 342312 86368
rect 340144 48272 340196 48278
rect 340144 48214 340196 48220
rect 340880 47592 340932 47598
rect 340878 47560 340880 47569
rect 340932 47560 340934 47569
rect 340878 47495 340934 47504
rect 342272 16574 342300 86362
rect 343008 86290 343036 176666
rect 343652 142118 343680 368766
rect 345664 361684 345716 361690
rect 345664 361626 345716 361632
rect 343732 228472 343784 228478
rect 343732 228414 343784 228420
rect 343640 142112 343692 142118
rect 343640 142054 343692 142060
rect 343744 115938 343772 228414
rect 343824 192568 343876 192574
rect 343824 192510 343876 192516
rect 343836 149734 343864 192510
rect 345204 185768 345256 185774
rect 345204 185710 345256 185716
rect 345020 183048 345072 183054
rect 345020 182990 345072 182996
rect 344284 158772 344336 158778
rect 344284 158714 344336 158720
rect 343824 149728 343876 149734
rect 343824 149670 343876 149676
rect 343732 115932 343784 115938
rect 343732 115874 343784 115880
rect 343638 96384 343694 96393
rect 343638 96319 343694 96328
rect 343652 95946 343680 96319
rect 343640 95940 343692 95946
rect 343640 95882 343692 95888
rect 342996 86284 343048 86290
rect 342996 86226 343048 86232
rect 342352 41404 342404 41410
rect 342352 41346 342404 41352
rect 342364 41313 342392 41346
rect 342350 41304 342406 41313
rect 342350 41239 342406 41248
rect 342364 40118 342392 41239
rect 342352 40112 342404 40118
rect 342352 40054 342404 40060
rect 342272 16546 342944 16574
rect 342166 11792 342222 11801
rect 342166 11727 342222 11736
rect 340972 8968 341024 8974
rect 340972 8910 341024 8916
rect 339960 8288 340012 8294
rect 339958 8256 339960 8265
rect 340012 8256 340014 8265
rect 339958 8191 340014 8200
rect 339972 6934 340000 8191
rect 339960 6928 340012 6934
rect 339960 6870 340012 6876
rect 340984 480 341012 8910
rect 342180 480 342208 11727
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 354 342944 16546
rect 343652 6914 343680 95882
rect 344296 8226 344324 158714
rect 345032 114510 345060 182990
rect 345110 177304 345166 177313
rect 345110 177239 345166 177248
rect 345124 118658 345152 177239
rect 345216 144906 345244 185710
rect 345676 184346 345704 361626
rect 345664 184340 345716 184346
rect 345664 184282 345716 184288
rect 345296 184272 345348 184278
rect 345296 184214 345348 184220
rect 345308 150414 345336 184214
rect 345296 150408 345348 150414
rect 345296 150350 345348 150356
rect 345664 146328 345716 146334
rect 345664 146270 345716 146276
rect 345204 144900 345256 144906
rect 345204 144842 345256 144848
rect 345112 118652 345164 118658
rect 345112 118594 345164 118600
rect 345020 114504 345072 114510
rect 345020 114446 345072 114452
rect 345018 98696 345074 98705
rect 345018 98631 345074 98640
rect 345032 16574 345060 98631
rect 345676 86358 345704 146270
rect 346412 125594 346440 378150
rect 347780 375488 347832 375494
rect 347780 375430 347832 375436
rect 346492 207052 346544 207058
rect 346492 206994 346544 207000
rect 346504 131102 346532 206994
rect 346584 178764 346636 178770
rect 346584 178706 346636 178712
rect 346596 139398 346624 178706
rect 347044 178084 347096 178090
rect 347044 178026 347096 178032
rect 346584 139392 346636 139398
rect 346584 139334 346636 139340
rect 346492 131096 346544 131102
rect 346492 131038 346544 131044
rect 346400 125588 346452 125594
rect 346400 125530 346452 125536
rect 347056 87650 347084 178026
rect 347792 124098 347820 375430
rect 349160 236020 349212 236026
rect 349160 235962 349212 235968
rect 347872 221536 347924 221542
rect 347872 221478 347924 221484
rect 347884 151774 347912 221478
rect 347962 181384 348018 181393
rect 347962 181319 348018 181328
rect 347872 151768 347924 151774
rect 347872 151710 347924 151716
rect 347780 124092 347832 124098
rect 347780 124034 347832 124040
rect 347976 122806 348004 181319
rect 348424 167680 348476 167686
rect 348424 167622 348476 167628
rect 347964 122800 348016 122806
rect 347964 122742 348016 122748
rect 347044 87644 347096 87650
rect 347044 87586 347096 87592
rect 345664 86352 345716 86358
rect 345664 86294 345716 86300
rect 345754 81424 345810 81433
rect 345754 81359 345756 81368
rect 345808 81359 345810 81368
rect 345756 81330 345808 81336
rect 345768 80102 345796 81330
rect 345756 80096 345808 80102
rect 345756 80038 345808 80044
rect 347044 69828 347096 69834
rect 347044 69770 347096 69776
rect 345032 16546 345336 16574
rect 344284 8220 344336 8226
rect 344284 8162 344336 8168
rect 343652 6886 344600 6914
rect 344572 480 344600 6886
rect 343334 354 343446 480
rect 342916 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 345308 354 345336 16546
rect 347056 4010 347084 69770
rect 348436 46889 348464 167622
rect 349172 113150 349200 235962
rect 349252 180192 349304 180198
rect 349252 180134 349304 180140
rect 349264 124166 349292 180134
rect 349344 176112 349396 176118
rect 349344 176054 349396 176060
rect 349356 129742 349384 176054
rect 349344 129736 349396 129742
rect 349344 129678 349396 129684
rect 349252 124160 349304 124166
rect 349252 124102 349304 124108
rect 349160 113144 349212 113150
rect 349160 113086 349212 113092
rect 349160 49700 349212 49706
rect 349160 49642 349212 49648
rect 347778 46880 347834 46889
rect 347778 46815 347834 46824
rect 348422 46880 348478 46889
rect 348422 46815 348478 46824
rect 347792 16574 347820 46815
rect 349172 16574 349200 49642
rect 347792 16546 348096 16574
rect 349172 16546 349292 16574
rect 347044 4004 347096 4010
rect 347044 3946 347096 3952
rect 347056 3890 347084 3946
rect 346964 3862 347084 3890
rect 346964 480 346992 3862
rect 348068 480 348096 16546
rect 349264 480 349292 16546
rect 349816 4078 349844 382910
rect 350540 367192 350592 367198
rect 350540 367134 350592 367140
rect 350552 97986 350580 367134
rect 351920 363180 351972 363186
rect 351920 363122 351972 363128
rect 351184 185700 351236 185706
rect 351184 185642 351236 185648
rect 350632 177540 350684 177546
rect 350632 177482 350684 177488
rect 350644 128314 350672 177482
rect 350632 128308 350684 128314
rect 350632 128250 350684 128256
rect 350540 97980 350592 97986
rect 350540 97922 350592 97928
rect 349804 4072 349856 4078
rect 349804 4014 349856 4020
rect 350448 4072 350500 4078
rect 350448 4014 350500 4020
rect 350460 480 350488 4014
rect 351196 3942 351224 185642
rect 351932 136610 351960 363122
rect 352564 360528 352616 360534
rect 352564 360470 352616 360476
rect 352012 195356 352064 195362
rect 352012 195298 352064 195304
rect 351920 136604 351972 136610
rect 351920 136546 351972 136552
rect 352024 49706 352052 195298
rect 352576 181626 352604 360470
rect 352656 342916 352708 342922
rect 352656 342858 352708 342864
rect 352668 333266 352696 342858
rect 352656 333260 352708 333266
rect 352656 333202 352708 333208
rect 352564 181620 352616 181626
rect 352564 181562 352616 181568
rect 352656 143608 352708 143614
rect 352656 143550 352708 143556
rect 352668 89078 352696 143550
rect 353312 142118 353340 409838
rect 358820 398880 358872 398886
rect 358820 398822 358872 398828
rect 353944 378208 353996 378214
rect 353944 378150 353996 378156
rect 353956 360369 353984 378150
rect 357440 374196 357492 374202
rect 357440 374138 357492 374144
rect 356704 360868 356756 360874
rect 356704 360810 356756 360816
rect 353390 360360 353446 360369
rect 353390 360295 353446 360304
rect 353942 360360 353998 360369
rect 353942 360295 353998 360304
rect 353404 297430 353432 360295
rect 354678 359544 354734 359553
rect 354678 359479 354734 359488
rect 353392 297424 353444 297430
rect 353392 297366 353444 297372
rect 353944 171148 353996 171154
rect 353944 171090 353996 171096
rect 353300 142112 353352 142118
rect 353300 142054 353352 142060
rect 353312 141438 353340 142054
rect 353300 141432 353352 141438
rect 353300 141374 353352 141380
rect 352656 89072 352708 89078
rect 352656 89014 352708 89020
rect 352564 89004 352616 89010
rect 352564 88946 352616 88952
rect 352012 49700 352064 49706
rect 352012 49642 352064 49648
rect 352576 4146 352604 88946
rect 353956 11830 353984 171090
rect 354036 137284 354088 137290
rect 354036 137226 354088 137232
rect 354048 104174 354076 137226
rect 354692 107642 354720 359479
rect 356060 347064 356112 347070
rect 356060 347006 356112 347012
rect 356072 146266 356100 347006
rect 356060 146260 356112 146266
rect 356060 146202 356112 146208
rect 354680 107636 354732 107642
rect 354680 107578 354732 107584
rect 356716 104854 356744 360810
rect 357452 168366 357480 374138
rect 358084 366036 358136 366042
rect 358084 365978 358136 365984
rect 357532 192500 357584 192506
rect 357532 192442 357584 192448
rect 357440 168360 357492 168366
rect 357440 168302 357492 168308
rect 356796 153264 356848 153270
rect 356796 153206 356848 153212
rect 356704 104848 356756 104854
rect 356704 104790 356756 104796
rect 354036 104168 354088 104174
rect 354036 104110 354088 104116
rect 354036 87644 354088 87650
rect 354036 87586 354088 87592
rect 353944 11824 353996 11830
rect 353944 11766 353996 11772
rect 352564 4140 352616 4146
rect 352564 4082 352616 4088
rect 354048 4010 354076 87586
rect 356808 4826 356836 153206
rect 357544 86426 357572 192442
rect 358096 186998 358124 365978
rect 358084 186992 358136 186998
rect 358084 186934 358136 186940
rect 358084 173936 358136 173942
rect 358084 173878 358136 173884
rect 357532 86420 357584 86426
rect 357532 86362 357584 86368
rect 358096 13734 358124 173878
rect 358832 137970 358860 398822
rect 359462 361992 359518 362001
rect 359462 361927 359518 361936
rect 359476 180198 359504 361927
rect 360844 361888 360896 361894
rect 360844 361830 360896 361836
rect 360200 207732 360252 207738
rect 360200 207674 360252 207680
rect 359464 180192 359516 180198
rect 359464 180134 359516 180140
rect 359464 164280 359516 164286
rect 359464 164222 359516 164228
rect 358820 137964 358872 137970
rect 358820 137906 358872 137912
rect 358832 137290 358860 137906
rect 358820 137284 358872 137290
rect 358820 137226 358872 137232
rect 358176 86964 358228 86970
rect 358176 86906 358228 86912
rect 358188 86426 358216 86906
rect 358176 86420 358228 86426
rect 358176 86362 358228 86368
rect 359476 49638 359504 164222
rect 360212 99385 360240 207674
rect 360856 192506 360884 361830
rect 364260 287094 364288 700726
rect 385684 590708 385736 590714
rect 385684 590650 385736 590656
rect 367100 403028 367152 403034
rect 367100 402970 367152 402976
rect 362960 287088 363012 287094
rect 362960 287030 363012 287036
rect 364248 287088 364300 287094
rect 364248 287030 364300 287036
rect 362972 286346 363000 287030
rect 362960 286340 363012 286346
rect 362960 286282 363012 286288
rect 362958 221504 363014 221513
rect 362958 221439 363014 221448
rect 360844 192500 360896 192506
rect 360844 192442 360896 192448
rect 360844 150476 360896 150482
rect 360844 150418 360896 150424
rect 360198 99376 360254 99385
rect 360198 99311 360254 99320
rect 360212 98705 360240 99311
rect 360198 98696 360254 98705
rect 360198 98631 360254 98640
rect 359464 49632 359516 49638
rect 359464 49574 359516 49580
rect 360856 44878 360884 150418
rect 362972 70378 363000 221439
rect 363604 149116 363656 149122
rect 363604 149058 363656 149064
rect 362960 70372 363012 70378
rect 362960 70314 363012 70320
rect 362972 69698 363000 70314
rect 362960 69692 363012 69698
rect 362960 69634 363012 69640
rect 360844 44872 360896 44878
rect 360844 44814 360896 44820
rect 358084 13728 358136 13734
rect 358084 13670 358136 13676
rect 363616 6798 363644 149058
rect 367112 46238 367140 402970
rect 385696 394806 385724 590650
rect 385684 394800 385736 394806
rect 385684 394742 385736 394748
rect 371884 367396 371936 367402
rect 371884 367338 371936 367344
rect 370504 293276 370556 293282
rect 370504 293218 370556 293224
rect 370516 260166 370544 293218
rect 370504 260160 370556 260166
rect 370504 260102 370556 260108
rect 367744 209160 367796 209166
rect 367744 209102 367796 209108
rect 367756 132462 367784 209102
rect 369860 193860 369912 193866
rect 369860 193802 369912 193808
rect 367836 139460 367888 139466
rect 367836 139402 367888 139408
rect 367744 132456 367796 132462
rect 367744 132398 367796 132404
rect 367848 102814 367876 139402
rect 367836 102808 367888 102814
rect 367836 102750 367888 102756
rect 367836 46912 367888 46918
rect 367836 46854 367888 46860
rect 367848 46238 367876 46854
rect 367100 46232 367152 46238
rect 367100 46174 367152 46180
rect 367836 46232 367888 46238
rect 367836 46174 367888 46180
rect 369872 9654 369900 193802
rect 370504 135312 370556 135318
rect 370504 135254 370556 135260
rect 370516 100026 370544 135254
rect 371896 118658 371924 367338
rect 375932 324964 375984 324970
rect 375932 324906 375984 324912
rect 375944 324358 375972 324906
rect 375932 324352 375984 324358
rect 375932 324294 375984 324300
rect 376668 324352 376720 324358
rect 376668 324294 376720 324300
rect 374644 245676 374696 245682
rect 374644 245618 374696 245624
rect 374656 133890 374684 245618
rect 374644 133884 374696 133890
rect 374644 133826 374696 133832
rect 376680 122806 376708 324294
rect 377404 309800 377456 309806
rect 377404 309742 377456 309748
rect 376668 122800 376720 122806
rect 376668 122742 376720 122748
rect 371884 118652 371936 118658
rect 371884 118594 371936 118600
rect 377416 110430 377444 309742
rect 382924 273964 382976 273970
rect 382924 273906 382976 273912
rect 378784 244316 378836 244322
rect 378784 244258 378836 244264
rect 377404 110424 377456 110430
rect 377404 110366 377456 110372
rect 378796 100706 378824 244258
rect 381544 202156 381596 202162
rect 381544 202098 381596 202104
rect 378784 100700 378836 100706
rect 378784 100642 378836 100648
rect 370504 100020 370556 100026
rect 370504 99962 370556 99968
rect 381556 95169 381584 202098
rect 382936 128314 382964 273906
rect 382924 128308 382976 128314
rect 382924 128250 382976 128256
rect 385696 114510 385724 394742
rect 403624 372700 403676 372706
rect 403624 372642 403676 372648
rect 395344 364540 395396 364546
rect 395344 364482 395396 364488
rect 388444 336048 388496 336054
rect 388444 335990 388496 335996
rect 385684 114504 385736 114510
rect 385684 114446 385736 114452
rect 388456 111790 388484 335990
rect 389824 214736 389876 214742
rect 389824 214678 389876 214684
rect 388444 111784 388496 111790
rect 388444 111726 388496 111732
rect 389836 107642 389864 214678
rect 393964 213240 394016 213246
rect 393964 213182 394016 213188
rect 392584 203584 392636 203590
rect 392584 203526 392636 203532
rect 389824 107636 389876 107642
rect 389824 107578 389876 107584
rect 392596 97986 392624 203526
rect 393976 103494 394004 213182
rect 393964 103488 394016 103494
rect 393964 103430 394016 103436
rect 395356 100638 395384 364482
rect 399484 361820 399536 361826
rect 399484 361762 399536 361768
rect 396724 175976 396776 175982
rect 396724 175918 396776 175924
rect 396736 102134 396764 175918
rect 396724 102128 396776 102134
rect 396724 102070 396776 102076
rect 395344 100632 395396 100638
rect 395344 100574 395396 100580
rect 399496 99278 399524 361762
rect 400864 271924 400916 271930
rect 400864 271866 400916 271872
rect 400876 184278 400904 271866
rect 400864 184272 400916 184278
rect 400864 184214 400916 184220
rect 403636 183530 403664 372642
rect 411904 372632 411956 372638
rect 411904 372574 411956 372580
rect 410524 361616 410576 361622
rect 410524 361558 410576 361564
rect 406384 360392 406436 360398
rect 406384 360334 406436 360340
rect 403624 183524 403676 183530
rect 403624 183466 403676 183472
rect 404268 183524 404320 183530
rect 404268 183466 404320 183472
rect 400864 182300 400916 182306
rect 400864 182242 400916 182248
rect 399484 99272 399536 99278
rect 399484 99214 399536 99220
rect 392584 97980 392636 97986
rect 392584 97922 392636 97928
rect 381542 95160 381598 95169
rect 381542 95095 381598 95104
rect 377404 86284 377456 86290
rect 377404 86226 377456 86232
rect 369860 9648 369912 9654
rect 369860 9590 369912 9596
rect 369872 8974 369900 9590
rect 369860 8968 369912 8974
rect 369860 8910 369912 8916
rect 363604 6792 363656 6798
rect 363604 6734 363656 6740
rect 356796 4820 356848 4826
rect 356796 4762 356848 4768
rect 377416 4078 377444 86226
rect 400876 59362 400904 182242
rect 404280 182238 404308 183466
rect 404268 182232 404320 182238
rect 404268 182174 404320 182180
rect 404280 133210 404308 182174
rect 404268 133204 404320 133210
rect 404268 133146 404320 133152
rect 406396 96626 406424 360334
rect 407764 297424 407816 297430
rect 407764 297366 407816 297372
rect 407776 121446 407804 297366
rect 407764 121440 407816 121446
rect 407764 121382 407816 121388
rect 410536 97918 410564 361558
rect 411916 180266 411944 372574
rect 417424 369980 417476 369986
rect 417424 369922 417476 369928
rect 414664 364472 414716 364478
rect 414664 364414 414716 364420
rect 413284 311160 413336 311166
rect 413284 311102 413336 311108
rect 411904 180260 411956 180266
rect 411904 180202 411956 180208
rect 413296 112946 413324 311102
rect 414676 181694 414704 364414
rect 417436 271930 417464 369922
rect 427820 340196 427872 340202
rect 427820 340138 427872 340144
rect 420920 290488 420972 290494
rect 420920 290430 420972 290436
rect 417424 271924 417476 271930
rect 417424 271866 417476 271872
rect 419540 271924 419592 271930
rect 419540 271866 419592 271872
rect 418804 231872 418856 231878
rect 418804 231814 418856 231820
rect 418816 227730 418844 231814
rect 418804 227724 418856 227730
rect 418804 227666 418856 227672
rect 417424 210452 417476 210458
rect 417424 210394 417476 210400
rect 414664 181688 414716 181694
rect 414664 181630 414716 181636
rect 416778 178664 416834 178673
rect 416778 178599 416834 178608
rect 416792 178090 416820 178599
rect 416780 178084 416832 178090
rect 416780 178026 416832 178032
rect 416778 177032 416834 177041
rect 416778 176967 416834 176976
rect 416792 176730 416820 176967
rect 416780 176724 416832 176730
rect 416780 176666 416832 176672
rect 416778 175264 416834 175273
rect 416778 175199 416834 175208
rect 416792 173942 416820 175199
rect 416780 173936 416832 173942
rect 416780 173878 416832 173884
rect 416778 171864 416834 171873
rect 416778 171799 416834 171808
rect 416792 171154 416820 171799
rect 416780 171148 416832 171154
rect 416780 171090 416832 171096
rect 416778 168464 416834 168473
rect 414664 168428 414716 168434
rect 416778 168399 416780 168408
rect 414664 168370 414716 168376
rect 416832 168399 416834 168408
rect 416780 168370 416832 168376
rect 413284 112940 413336 112946
rect 413284 112882 413336 112888
rect 410524 97912 410576 97918
rect 410524 97854 410576 97860
rect 406384 96620 406436 96626
rect 406384 96562 406436 96568
rect 414676 73098 414704 168370
rect 416778 166832 416834 166841
rect 416778 166767 416834 166776
rect 416792 165646 416820 166767
rect 416780 165640 416832 165646
rect 416780 165582 416832 165588
rect 416778 165064 416834 165073
rect 416778 164999 416834 165008
rect 416792 164286 416820 164999
rect 416780 164280 416832 164286
rect 416780 164222 416832 164228
rect 416778 163432 416834 163441
rect 416778 163367 416834 163376
rect 416792 162926 416820 163367
rect 416780 162920 416832 162926
rect 416780 162862 416832 162868
rect 416778 161800 416834 161809
rect 416778 161735 416834 161744
rect 416792 161498 416820 161735
rect 416780 161492 416832 161498
rect 416780 161434 416832 161440
rect 416778 160032 416834 160041
rect 416778 159967 416834 159976
rect 416792 158778 416820 159967
rect 416780 158772 416832 158778
rect 416780 158714 416832 158720
rect 416778 156632 416834 156641
rect 416778 156567 416834 156576
rect 416792 155990 416820 156567
rect 416780 155984 416832 155990
rect 416780 155926 416832 155932
rect 416778 155000 416834 155009
rect 416778 154935 416834 154944
rect 416792 154630 416820 154935
rect 416780 154624 416832 154630
rect 416780 154566 416832 154572
rect 416780 153264 416832 153270
rect 416778 153232 416780 153241
rect 416832 153232 416834 153241
rect 416778 153167 416834 153176
rect 416778 151600 416834 151609
rect 416778 151535 416834 151544
rect 416792 150482 416820 151535
rect 416780 150476 416832 150482
rect 416780 150418 416832 150424
rect 416778 149832 416834 149841
rect 416778 149767 416834 149776
rect 416792 149122 416820 149767
rect 416780 149116 416832 149122
rect 416780 149058 416832 149064
rect 416778 148200 416834 148209
rect 416778 148135 416834 148144
rect 416792 147694 416820 148135
rect 416780 147688 416832 147694
rect 416780 147630 416832 147636
rect 416778 146568 416834 146577
rect 416778 146503 416834 146512
rect 416792 146334 416820 146503
rect 416780 146328 416832 146334
rect 416780 146270 416832 146276
rect 416778 144800 416834 144809
rect 416778 144735 416834 144744
rect 416792 143614 416820 144735
rect 416780 143608 416832 143614
rect 416780 143550 416832 143556
rect 416870 143168 416926 143177
rect 416870 143103 416926 143112
rect 416884 142186 416912 143103
rect 416872 142180 416924 142186
rect 416872 142122 416924 142128
rect 416780 142112 416832 142118
rect 416780 142054 416832 142060
rect 416792 141409 416820 142054
rect 416778 141400 416834 141409
rect 416778 141335 416834 141344
rect 416778 139768 416834 139777
rect 416778 139703 416834 139712
rect 416792 139466 416820 139703
rect 416780 139460 416832 139466
rect 416780 139402 416832 139408
rect 416778 138000 416834 138009
rect 416778 137935 416780 137944
rect 416832 137935 416834 137944
rect 416780 137906 416832 137912
rect 416778 136368 416834 136377
rect 416778 136303 416834 136312
rect 416792 135318 416820 136303
rect 416780 135312 416832 135318
rect 416780 135254 416832 135260
rect 417332 135244 417384 135250
rect 417332 135186 417384 135192
rect 417344 134609 417372 135186
rect 417330 134600 417386 134609
rect 417330 134535 417386 134544
rect 416780 122800 416832 122806
rect 416778 122768 416780 122777
rect 416832 122768 416834 122777
rect 416778 122703 416834 122712
rect 416780 121440 416832 121446
rect 416780 121382 416832 121388
rect 416792 121145 416820 121382
rect 416778 121136 416834 121145
rect 416778 121071 416834 121080
rect 417436 119377 417464 210394
rect 417516 132456 417568 132462
rect 417516 132398 417568 132404
rect 417528 131345 417556 132398
rect 417514 131336 417570 131345
rect 417514 131271 417570 131280
rect 418712 128308 418764 128314
rect 418712 128250 418764 128256
rect 418724 127945 418752 128250
rect 418710 127936 418766 127945
rect 418710 127871 418766 127880
rect 418816 126177 418844 227666
rect 419356 182844 419408 182850
rect 419356 182786 419408 182792
rect 419262 134600 419318 134609
rect 419262 134535 419318 134544
rect 418802 126168 418858 126177
rect 418802 126103 418858 126112
rect 417422 119368 417478 119377
rect 417422 119303 417478 119312
rect 416780 118652 416832 118658
rect 416780 118594 416832 118600
rect 416792 117745 416820 118594
rect 416778 117736 416834 117745
rect 416778 117671 416834 117680
rect 416780 117292 416832 117298
rect 416780 117234 416832 117240
rect 416792 116113 416820 117234
rect 416778 116104 416834 116113
rect 416778 116039 416834 116048
rect 416780 114504 416832 114510
rect 416780 114446 416832 114452
rect 416792 114345 416820 114446
rect 416778 114336 416834 114345
rect 416778 114271 416834 114280
rect 416780 112940 416832 112946
rect 416780 112882 416832 112888
rect 416792 112713 416820 112882
rect 416778 112704 416834 112713
rect 416778 112639 416834 112648
rect 416780 111784 416832 111790
rect 416780 111726 416832 111732
rect 416792 110945 416820 111726
rect 416778 110936 416834 110945
rect 416778 110871 416834 110880
rect 416780 110424 416832 110430
rect 416780 110366 416832 110372
rect 416792 109313 416820 110366
rect 416778 109304 416834 109313
rect 416778 109239 416834 109248
rect 416780 107636 416832 107642
rect 416780 107578 416832 107584
rect 416792 107545 416820 107578
rect 416778 107536 416834 107545
rect 416778 107471 416834 107480
rect 416780 106276 416832 106282
rect 416780 106218 416832 106224
rect 416792 105913 416820 106218
rect 416778 105904 416834 105913
rect 416778 105839 416834 105848
rect 416780 104848 416832 104854
rect 416780 104790 416832 104796
rect 416792 104145 416820 104790
rect 416778 104136 416834 104145
rect 416778 104071 416834 104080
rect 416780 103488 416832 103494
rect 416780 103430 416832 103436
rect 416792 102513 416820 103430
rect 416778 102504 416834 102513
rect 416778 102439 416834 102448
rect 416780 102128 416832 102134
rect 416780 102070 416832 102076
rect 416792 100881 416820 102070
rect 416778 100872 416834 100881
rect 416778 100807 416834 100816
rect 417424 96824 417476 96830
rect 417424 96766 417476 96772
rect 414664 73092 414716 73098
rect 414664 73034 414716 73040
rect 400864 59356 400916 59362
rect 400864 59298 400916 59304
rect 417436 14482 417464 96766
rect 419276 93158 419304 134535
rect 419368 127945 419396 182786
rect 419448 133884 419500 133890
rect 419448 133826 419500 133832
rect 419460 132977 419488 133826
rect 419446 132968 419502 132977
rect 419446 132903 419502 132912
rect 419354 127936 419410 127945
rect 419354 127871 419410 127880
rect 419264 93152 419316 93158
rect 419264 93094 419316 93100
rect 419460 73166 419488 132903
rect 419552 124545 419580 271866
rect 420932 179466 420960 290430
rect 425060 258120 425112 258126
rect 425060 258062 425112 258068
rect 425072 190454 425100 258062
rect 425072 190426 425376 190454
rect 422944 185700 422996 185706
rect 422944 185642 422996 185648
rect 422956 179466 422984 185642
rect 425348 179466 425376 190426
rect 427832 179466 427860 340138
rect 429212 301510 429240 702782
rect 478524 702778 478552 703520
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 494808 702710 494836 703520
rect 453948 702704 454000 702710
rect 453948 702646 454000 702652
rect 492588 702704 492640 702710
rect 492588 702646 492640 702652
rect 494796 702704 494848 702710
rect 494796 702646 494848 702652
rect 453960 700330 453988 702646
rect 492600 700330 492628 702646
rect 521568 702568 521620 702574
rect 521568 702510 521620 702516
rect 521580 701010 521608 702510
rect 527192 702506 527220 703520
rect 543476 702545 543504 703520
rect 559668 702574 559696 703520
rect 580908 702636 580960 702642
rect 580908 702578 580960 702584
rect 550548 702568 550600 702574
rect 543462 702536 543518 702545
rect 527180 702500 527232 702506
rect 550548 702510 550600 702516
rect 559656 702568 559708 702574
rect 559656 702510 559708 702516
rect 543462 702471 543518 702480
rect 527180 702442 527232 702448
rect 519544 701004 519596 701010
rect 519544 700946 519596 700952
rect 521568 701004 521620 701010
rect 521568 700946 521620 700952
rect 450544 700324 450596 700330
rect 450544 700266 450596 700272
rect 453948 700324 454000 700330
rect 453948 700266 454000 700272
rect 492588 700324 492640 700330
rect 492588 700266 492640 700272
rect 431224 510672 431276 510678
rect 431224 510614 431276 510620
rect 429200 301504 429252 301510
rect 429200 301446 429252 301452
rect 431236 220794 431264 510614
rect 446404 456816 446456 456822
rect 446404 456758 446456 456764
rect 434720 248464 434772 248470
rect 434720 248406 434772 248412
rect 432604 234660 432656 234666
rect 432604 234602 432656 234608
rect 429844 220788 429896 220794
rect 429844 220730 429896 220736
rect 431224 220788 431276 220794
rect 431224 220730 431276 220736
rect 429856 220114 429884 220730
rect 429844 220108 429896 220114
rect 429844 220050 429896 220056
rect 429856 190454 429884 220050
rect 432616 211138 432644 234602
rect 432604 211132 432656 211138
rect 432604 211074 432656 211080
rect 432616 210730 432644 211074
rect 431960 210724 432012 210730
rect 431960 210666 432012 210672
rect 432604 210724 432656 210730
rect 432604 210666 432656 210672
rect 431972 190454 432000 210666
rect 429856 190426 429976 190454
rect 431972 190426 432368 190454
rect 429948 179466 429976 190426
rect 432340 179466 432368 190426
rect 434732 179466 434760 248406
rect 438860 238060 438912 238066
rect 438860 238002 438912 238008
rect 436100 217320 436152 217326
rect 436100 217262 436152 217268
rect 436112 190454 436140 217262
rect 438872 190454 438900 238002
rect 446416 211138 446444 456758
rect 447784 307080 447836 307086
rect 447784 307022 447836 307028
rect 446404 211132 446456 211138
rect 446404 211074 446456 211080
rect 447796 210458 447824 307022
rect 449164 242956 449216 242962
rect 449164 242898 449216 242904
rect 447784 210452 447836 210458
rect 447784 210394 447836 210400
rect 436112 190426 436968 190454
rect 438872 190426 439360 190454
rect 436940 179466 436968 190426
rect 439332 179466 439360 190426
rect 443920 184340 443972 184346
rect 443920 184282 443972 184288
rect 441620 181688 441672 181694
rect 441620 181630 441672 181636
rect 441632 179466 441660 181630
rect 443932 179466 443960 184282
rect 448612 181620 448664 181626
rect 448612 181562 448664 181568
rect 446404 181552 446456 181558
rect 446404 181494 446456 181500
rect 446416 179466 446444 181494
rect 448624 179466 448652 181562
rect 449176 181558 449204 242898
rect 450556 185706 450584 700266
rect 497464 565140 497516 565146
rect 497464 565082 497516 565088
rect 504364 565140 504416 565146
rect 504364 565082 504416 565088
rect 471980 374060 472032 374066
rect 471980 374002 472032 374008
rect 464344 369912 464396 369918
rect 464344 369854 464396 369860
rect 457444 368552 457496 368558
rect 457444 368494 457496 368500
rect 452660 351212 452712 351218
rect 452660 351154 452712 351160
rect 451280 198008 451332 198014
rect 451280 197950 451332 197956
rect 451292 190454 451320 197950
rect 452672 190454 452700 351154
rect 454684 316736 454736 316742
rect 454684 316678 454736 316684
rect 451292 190426 451412 190454
rect 452672 190426 453160 190454
rect 450544 185700 450596 185706
rect 450544 185642 450596 185648
rect 449164 181552 449216 181558
rect 449164 181494 449216 181500
rect 451384 179466 451412 190426
rect 420932 179438 421130 179466
rect 422956 179438 423430 179466
rect 425348 179438 425730 179466
rect 427832 179438 428030 179466
rect 429948 179438 430422 179466
rect 432340 179438 432722 179466
rect 434732 179438 435022 179466
rect 436940 179438 437322 179466
rect 439332 179438 439714 179466
rect 441632 179438 442014 179466
rect 443932 179438 444314 179466
rect 446416 179438 446706 179466
rect 448624 179438 449006 179466
rect 451306 179438 451412 179466
rect 453132 179466 453160 190426
rect 454696 182170 454724 316678
rect 454684 182164 454736 182170
rect 454684 182106 454736 182112
rect 455604 182164 455656 182170
rect 455604 182106 455656 182112
rect 455616 179466 455644 182106
rect 457456 181694 457484 368494
rect 458180 355360 458232 355366
rect 458180 355302 458232 355308
rect 457444 181688 457496 181694
rect 457444 181630 457496 181636
rect 458192 179466 458220 355302
rect 461584 345092 461636 345098
rect 461584 345034 461636 345040
rect 460112 189780 460164 189786
rect 460112 189722 460164 189728
rect 460124 179466 460152 189722
rect 461596 182170 461624 345034
rect 461584 182164 461636 182170
rect 461584 182106 461636 182112
rect 462596 182164 462648 182170
rect 462596 182106 462648 182112
rect 462608 179466 462636 182106
rect 464356 181626 464384 369854
rect 466460 363044 466512 363050
rect 466460 362986 466512 362992
rect 465080 333260 465132 333266
rect 465080 333202 465132 333208
rect 464344 181620 464396 181626
rect 464344 181562 464396 181568
rect 465092 179466 465120 333202
rect 466472 190454 466500 362986
rect 469220 358080 469272 358086
rect 469220 358022 469272 358028
rect 468484 300892 468536 300898
rect 468484 300834 468536 300840
rect 466472 190426 467144 190454
rect 467116 179466 467144 190426
rect 468496 184346 468524 300834
rect 469232 190454 469260 358022
rect 471244 222896 471296 222902
rect 471244 222838 471296 222844
rect 469232 190426 469536 190454
rect 468484 184340 468536 184346
rect 468484 184282 468536 184288
rect 469508 179466 469536 190426
rect 471256 182170 471284 222838
rect 471244 182164 471296 182170
rect 471244 182106 471296 182112
rect 471992 179466 472020 374002
rect 475384 365900 475436 365906
rect 475384 365842 475436 365848
rect 475396 181762 475424 365842
rect 495440 358828 495492 358834
rect 495440 358770 495492 358776
rect 489184 349852 489236 349858
rect 489184 349794 489236 349800
rect 482284 327752 482336 327758
rect 482284 327694 482336 327700
rect 478880 224256 478932 224262
rect 478880 224198 478932 224204
rect 476580 182164 476632 182170
rect 476580 182106 476632 182112
rect 475384 181756 475436 181762
rect 475384 181698 475436 181704
rect 474188 181688 474240 181694
rect 474188 181630 474240 181636
rect 474200 179466 474228 181630
rect 476592 179466 476620 182106
rect 478892 179466 478920 224198
rect 480260 210452 480312 210458
rect 480260 210394 480312 210400
rect 480272 190454 480300 210394
rect 480272 190426 481128 190454
rect 481100 179466 481128 190426
rect 482296 181694 482324 327694
rect 485044 225616 485096 225622
rect 485044 225558 485096 225564
rect 483020 217388 483072 217394
rect 483020 217330 483072 217336
rect 483032 190454 483060 217330
rect 483032 190426 483520 190454
rect 482284 181688 482336 181694
rect 482284 181630 482336 181636
rect 483492 179466 483520 190426
rect 485056 182170 485084 225558
rect 486424 214600 486476 214606
rect 486424 214542 486476 214548
rect 485044 182164 485096 182170
rect 485044 182106 485096 182112
rect 485780 182164 485832 182170
rect 485780 182106 485832 182112
rect 485792 179466 485820 182106
rect 486436 181830 486464 214542
rect 489196 182374 489224 349794
rect 493876 342304 493928 342310
rect 493876 342246 493928 342252
rect 490564 263628 490616 263634
rect 490564 263570 490616 263576
rect 490576 190454 490604 263570
rect 490576 190426 490696 190454
rect 489184 182368 489236 182374
rect 489184 182310 489236 182316
rect 490564 182368 490616 182374
rect 490564 182310 490616 182316
rect 486424 181824 486476 181830
rect 486424 181766 486476 181772
rect 488632 181756 488684 181762
rect 488632 181698 488684 181704
rect 488644 179466 488672 181698
rect 453132 179438 453606 179466
rect 455616 179438 455998 179466
rect 458192 179438 458298 179466
rect 460124 179438 460598 179466
rect 462608 179438 462990 179466
rect 465092 179438 465290 179466
rect 467116 179438 467590 179466
rect 469508 179438 469890 179466
rect 471992 179438 472282 179466
rect 474200 179438 474582 179466
rect 476592 179438 476882 179466
rect 478892 179438 479274 179466
rect 481100 179438 481574 179466
rect 483492 179438 483874 179466
rect 485792 179438 486174 179466
rect 488566 179438 488672 179466
rect 490576 179466 490604 182310
rect 490668 180334 490696 190426
rect 492864 181824 492916 181830
rect 492864 181766 492916 181772
rect 490656 180328 490708 180334
rect 490656 180270 490708 180276
rect 492876 179466 492904 181766
rect 490576 179438 490866 179466
rect 492876 179438 493166 179466
rect 493888 178673 493916 342246
rect 494244 209092 494296 209098
rect 494244 209034 494296 209040
rect 494152 204944 494204 204950
rect 494152 204886 494204 204892
rect 494060 182300 494112 182306
rect 494060 182242 494112 182248
rect 494072 179353 494100 182242
rect 494058 179344 494114 179353
rect 494058 179279 494114 179288
rect 493874 178664 493930 178673
rect 493874 178599 493930 178608
rect 494058 168464 494114 168473
rect 494058 168399 494114 168408
rect 419632 133204 419684 133210
rect 419632 133146 419684 133152
rect 419644 129577 419672 133146
rect 419722 131336 419778 131345
rect 419722 131271 419778 131280
rect 419630 129568 419686 129577
rect 419630 129503 419686 129512
rect 419538 124536 419594 124545
rect 419538 124471 419594 124480
rect 419736 122834 419764 131271
rect 419644 122806 419764 122834
rect 419644 99346 419672 122806
rect 493968 100700 494020 100706
rect 493968 100642 494020 100648
rect 493980 100473 494008 100642
rect 493966 100464 494022 100473
rect 493966 100399 494022 100408
rect 419632 99340 419684 99346
rect 419632 99282 419684 99288
rect 420184 97368 420236 97374
rect 420184 97310 420236 97316
rect 420196 93226 420224 97310
rect 420564 96830 420592 100028
rect 420932 100014 421774 100042
rect 422312 100014 422970 100042
rect 423692 100014 424166 100042
rect 425072 100014 425362 100042
rect 420552 96824 420604 96830
rect 420552 96766 420604 96772
rect 420184 93220 420236 93226
rect 420184 93162 420236 93168
rect 420932 89690 420960 100014
rect 421564 97300 421616 97306
rect 421564 97242 421616 97248
rect 420920 89684 420972 89690
rect 420920 89626 420972 89632
rect 421576 86970 421604 97242
rect 421564 86964 421616 86970
rect 421564 86906 421616 86912
rect 419448 73160 419500 73166
rect 419448 73102 419500 73108
rect 422312 46918 422340 100014
rect 422300 46912 422352 46918
rect 422300 46854 422352 46860
rect 417424 14476 417476 14482
rect 417424 14418 417476 14424
rect 423692 9586 423720 100014
rect 425072 33114 425100 100014
rect 426544 94518 426572 100028
rect 427740 97374 427768 100028
rect 427832 100014 428950 100042
rect 429212 100014 430146 100042
rect 430592 100014 431342 100042
rect 431972 100014 432538 100042
rect 433352 100014 433734 100042
rect 434732 100014 434930 100042
rect 436126 100014 436232 100042
rect 427728 97368 427780 97374
rect 427728 97310 427780 97316
rect 426532 94512 426584 94518
rect 426532 94454 426584 94460
rect 427832 43450 427860 100014
rect 427820 43444 427872 43450
rect 427820 43386 427872 43392
rect 429212 42770 429240 100014
rect 429200 42764 429252 42770
rect 429200 42706 429252 42712
rect 430592 41410 430620 100014
rect 430580 41404 430632 41410
rect 430580 41346 430632 41352
rect 425060 33108 425112 33114
rect 425060 33050 425112 33056
rect 423680 9580 423732 9586
rect 423680 9522 423732 9528
rect 431972 8294 432000 100014
rect 433352 39370 433380 100014
rect 433340 39364 433392 39370
rect 433340 39306 433392 39312
rect 434732 37942 434760 100014
rect 434720 37936 434772 37942
rect 434720 37878 434772 37884
rect 436204 36582 436232 100014
rect 436296 100014 437322 100042
rect 437492 100014 438518 100042
rect 438872 100014 439714 100042
rect 436192 36576 436244 36582
rect 436192 36518 436244 36524
rect 436296 35222 436324 100014
rect 436284 35216 436336 35222
rect 436284 35158 436336 35164
rect 437492 34474 437520 100014
rect 437480 34468 437532 34474
rect 437480 34410 437532 34416
rect 438872 31210 438900 100014
rect 440896 96966 440924 100028
rect 441632 100014 442106 100042
rect 443012 100014 443302 100042
rect 444392 100014 444498 100042
rect 445786 100014 445892 100042
rect 439504 96960 439556 96966
rect 439504 96902 439556 96908
rect 440884 96960 440936 96966
rect 440884 96902 440936 96908
rect 438860 31204 438912 31210
rect 438860 31146 438912 31152
rect 431960 8288 432012 8294
rect 431960 8230 432012 8236
rect 439516 6866 439544 96902
rect 441632 30326 441660 100014
rect 441620 30320 441672 30326
rect 441620 30262 441672 30268
rect 443012 28354 443040 100014
rect 443000 28348 443052 28354
rect 443000 28290 443052 28296
rect 444392 26926 444420 100014
rect 444380 26920 444432 26926
rect 444380 26862 444432 26868
rect 445864 25634 445892 100014
rect 445956 100014 446982 100042
rect 447152 100014 448178 100042
rect 448532 100014 449374 100042
rect 449912 100014 450570 100042
rect 451292 100014 451766 100042
rect 452672 100014 452962 100042
rect 445852 25628 445904 25634
rect 445852 25570 445904 25576
rect 445956 24818 445984 100014
rect 445944 24812 445996 24818
rect 445944 24754 445996 24760
rect 447152 22846 447180 100014
rect 447140 22840 447192 22846
rect 447140 22782 447192 22788
rect 439504 6860 439556 6866
rect 439504 6802 439556 6808
rect 448532 5506 448560 100014
rect 449912 22098 449940 100014
rect 449900 22092 449952 22098
rect 449900 22034 449952 22040
rect 451292 20058 451320 100014
rect 451280 20052 451332 20058
rect 451280 19994 451332 20000
rect 452672 18630 452700 100014
rect 454040 96960 454092 96966
rect 454040 96902 454092 96908
rect 452660 18624 452712 18630
rect 452660 18566 452712 18572
rect 454052 16046 454080 96902
rect 454144 17406 454172 100028
rect 455064 100014 455354 100042
rect 455432 100014 456550 100042
rect 456812 100014 457746 100042
rect 455064 96966 455092 100014
rect 455052 96960 455104 96966
rect 455052 96902 455104 96908
rect 455432 86290 455460 100014
rect 456812 87650 456840 100014
rect 458928 97306 458956 100028
rect 459572 100014 460138 100042
rect 460952 100014 461334 100042
rect 462332 100014 462530 100042
rect 458916 97300 458968 97306
rect 458916 97242 458968 97248
rect 456800 87644 456852 87650
rect 456800 87586 456852 87592
rect 455420 86284 455472 86290
rect 455420 86226 455472 86232
rect 459572 70378 459600 100014
rect 460952 84862 460980 100014
rect 461584 96960 461636 96966
rect 461584 96902 461636 96908
rect 460940 84856 460992 84862
rect 460940 84798 460992 84804
rect 461596 82142 461624 96902
rect 462332 89010 462360 100014
rect 462320 89004 462372 89010
rect 462320 88946 462372 88952
rect 463712 83502 463740 100028
rect 464908 96966 464936 100028
rect 465092 100014 466118 100042
rect 464896 96960 464948 96966
rect 464896 96902 464948 96908
rect 465092 90370 465120 100014
rect 467104 97300 467156 97306
rect 467104 97242 467156 97248
rect 465724 96960 465776 96966
rect 465724 96902 465776 96908
rect 465080 90364 465132 90370
rect 465080 90306 465132 90312
rect 463700 83496 463752 83502
rect 463700 83438 463752 83444
rect 461584 82136 461636 82142
rect 461584 82078 461636 82084
rect 465736 81394 465764 96902
rect 465724 81388 465776 81394
rect 465724 81330 465776 81336
rect 459560 70372 459612 70378
rect 459560 70314 459612 70320
rect 467116 51882 467144 97242
rect 467300 96966 467328 100028
rect 467852 100014 468510 100042
rect 469232 100014 469706 100042
rect 470612 100014 470994 100042
rect 471992 100014 472190 100042
rect 467288 96960 467340 96966
rect 467288 96902 467340 96908
rect 467104 51876 467156 51882
rect 467104 51818 467156 51824
rect 454132 17400 454184 17406
rect 454132 17342 454184 17348
rect 454040 16040 454092 16046
rect 454040 15982 454092 15988
rect 467852 13802 467880 100014
rect 469232 73846 469260 100014
rect 470612 79354 470640 100014
rect 470600 79348 470652 79354
rect 470600 79290 470652 79296
rect 471992 78674 472020 100014
rect 472624 96960 472676 96966
rect 472624 96902 472676 96908
rect 471980 78668 472032 78674
rect 471980 78610 472032 78616
rect 472636 75206 472664 96902
rect 473372 76566 473400 100028
rect 474568 96966 474596 100028
rect 474752 100014 475778 100042
rect 476132 100014 476974 100042
rect 477512 100014 478170 100042
rect 478892 100014 479366 100042
rect 480272 100014 480562 100042
rect 474556 96960 474608 96966
rect 474556 96902 474608 96908
rect 473360 76560 473412 76566
rect 473360 76502 473412 76508
rect 472624 75200 472676 75206
rect 472624 75142 472676 75148
rect 469220 73840 469272 73846
rect 469220 73782 469272 73788
rect 474752 68338 474780 100014
rect 474740 68332 474792 68338
rect 474740 68274 474792 68280
rect 476132 66978 476160 100014
rect 476120 66972 476172 66978
rect 476120 66914 476172 66920
rect 477512 66230 477540 100014
rect 477500 66224 477552 66230
rect 477500 66166 477552 66172
rect 467840 13796 467892 13802
rect 467840 13738 467892 13744
rect 478892 11762 478920 100014
rect 480272 64258 480300 100014
rect 481640 96960 481692 96966
rect 481640 96902 481692 96908
rect 480260 64252 480312 64258
rect 480260 64194 480312 64200
rect 481652 61402 481680 96902
rect 481744 62830 481772 100028
rect 482664 100014 482954 100042
rect 483032 100014 484150 100042
rect 484412 100014 485346 100042
rect 485792 100014 486542 100042
rect 482664 96966 482692 100014
rect 482652 96960 482704 96966
rect 482652 96902 482704 96908
rect 481732 62824 481784 62830
rect 481732 62766 481784 62772
rect 481640 61396 481692 61402
rect 481640 61338 481692 61344
rect 483032 60110 483060 100014
rect 483020 60104 483072 60110
rect 483020 60046 483072 60052
rect 484412 58682 484440 100014
rect 484400 58676 484452 58682
rect 484400 58618 484452 58624
rect 485792 57934 485820 100014
rect 487724 96966 487752 100028
rect 488552 100014 488934 100042
rect 489932 100014 490130 100042
rect 486424 96960 486476 96966
rect 486424 96902 486476 96908
rect 487712 96960 487764 96966
rect 487712 96902 487764 96908
rect 485780 57928 485832 57934
rect 485780 57870 485832 57876
rect 478880 11756 478932 11762
rect 478880 11698 478932 11704
rect 486436 10334 486464 96902
rect 488552 55894 488580 100014
rect 488540 55888 488592 55894
rect 488540 55830 488592 55836
rect 489932 54534 489960 100014
rect 489920 54528 489972 54534
rect 489920 54470 489972 54476
rect 491312 53106 491340 100028
rect 492508 97306 492536 100028
rect 492692 100014 493718 100042
rect 492496 97300 492548 97306
rect 492496 97242 492548 97248
rect 491300 53100 491352 53106
rect 491300 53042 491352 53048
rect 492692 50454 492720 100014
rect 492680 50448 492732 50454
rect 492680 50390 492732 50396
rect 494072 49706 494100 168399
rect 494164 149025 494192 204886
rect 494150 149016 494206 149025
rect 494150 148951 494206 148960
rect 494150 146296 494206 146305
rect 494150 146231 494206 146240
rect 494164 71738 494192 146231
rect 494256 141273 494284 209034
rect 494336 188352 494388 188358
rect 494336 188294 494388 188300
rect 494242 141264 494298 141273
rect 494242 141199 494298 141208
rect 494348 132161 494376 188294
rect 495346 140856 495402 140865
rect 495346 140791 495348 140800
rect 495400 140791 495402 140800
rect 495348 140762 495400 140768
rect 494334 132152 494390 132161
rect 494334 132087 494390 132096
rect 495452 119649 495480 358770
rect 497476 340202 497504 565082
rect 504376 563718 504404 565082
rect 504364 563712 504416 563718
rect 504364 563654 504416 563660
rect 510620 362976 510672 362982
rect 510620 362918 510672 362924
rect 499578 360224 499634 360233
rect 499578 360159 499634 360168
rect 497464 340196 497516 340202
rect 497464 340138 497516 340144
rect 498292 237448 498344 237454
rect 498292 237390 498344 237396
rect 495624 228404 495676 228410
rect 495624 228346 495676 228352
rect 495530 173360 495586 173369
rect 495530 173295 495586 173304
rect 495438 119640 495494 119649
rect 495438 119575 495494 119584
rect 494242 104816 494298 104825
rect 494242 104751 494298 104760
rect 494256 100638 494284 104751
rect 495438 103864 495494 103873
rect 495438 103799 495494 103808
rect 494244 100632 494296 100638
rect 494244 100574 494296 100580
rect 495452 97986 495480 103799
rect 495440 97980 495492 97986
rect 495440 97922 495492 97928
rect 494152 71732 494204 71738
rect 494152 71674 494204 71680
rect 494060 49700 494112 49706
rect 494060 49642 494112 49648
rect 486424 10328 486476 10334
rect 486424 10270 486476 10276
rect 448520 5500 448572 5506
rect 448520 5442 448572 5448
rect 377404 4072 377456 4078
rect 377404 4014 377456 4020
rect 354036 4004 354088 4010
rect 354036 3946 354088 3952
rect 495544 3942 495572 173295
rect 495636 130801 495664 228346
rect 495716 222964 495768 222970
rect 495716 222906 495768 222912
rect 495728 164393 495756 222906
rect 497464 215960 497516 215966
rect 497464 215902 497516 215908
rect 497004 181484 497056 181490
rect 497004 181426 497056 181432
rect 496910 177848 496966 177857
rect 496910 177783 496966 177792
rect 496924 176798 496952 177783
rect 496912 176792 496964 176798
rect 496818 176760 496874 176769
rect 496912 176734 496964 176740
rect 496818 176695 496820 176704
rect 496872 176695 496874 176704
rect 496820 176666 496872 176672
rect 496818 175672 496874 175681
rect 496818 175607 496820 175616
rect 496872 175607 496874 175616
rect 496820 175578 496872 175584
rect 496820 168360 496872 168366
rect 496820 168302 496872 168308
rect 496832 167793 496860 168302
rect 496818 167784 496874 167793
rect 496818 167719 496874 167728
rect 496818 166696 496874 166705
rect 496818 166631 496874 166640
rect 496832 166326 496860 166631
rect 496820 166320 496872 166326
rect 496820 166262 496872 166268
rect 496818 165472 496874 165481
rect 496818 165407 496874 165416
rect 496832 164898 496860 165407
rect 496820 164892 496872 164898
rect 496820 164834 496872 164840
rect 495714 164384 495770 164393
rect 495714 164319 495770 164328
rect 496358 164384 496414 164393
rect 496358 164319 496414 164328
rect 496372 164286 496400 164319
rect 496360 164280 496412 164286
rect 496360 164222 496412 164228
rect 496820 164212 496872 164218
rect 496820 164154 496872 164160
rect 496832 163305 496860 164154
rect 496818 163296 496874 163305
rect 496818 163231 496874 163240
rect 496820 162852 496872 162858
rect 496820 162794 496872 162800
rect 496832 162217 496860 162794
rect 496818 162208 496874 162217
rect 496818 162143 496874 162152
rect 497016 161514 497044 181426
rect 497476 178702 497504 215902
rect 497464 178696 497516 178702
rect 497464 178638 497516 178644
rect 498106 171184 498162 171193
rect 498162 171142 498240 171170
rect 498106 171119 498162 171128
rect 496832 161486 497044 161514
rect 496832 150929 496860 161486
rect 496912 161424 496964 161430
rect 496912 161366 496964 161372
rect 496924 160993 496952 161366
rect 496910 160984 496966 160993
rect 496910 160919 496966 160928
rect 496912 160064 496964 160070
rect 496912 160006 496964 160012
rect 496924 159905 496952 160006
rect 497004 159996 497056 160002
rect 497004 159938 497056 159944
rect 496910 159896 496966 159905
rect 496910 159831 496966 159840
rect 497016 158817 497044 159938
rect 497002 158808 497058 158817
rect 497002 158743 497058 158752
rect 496912 158704 496964 158710
rect 496912 158646 496964 158652
rect 496924 157729 496952 158646
rect 496910 157720 496966 157729
rect 496910 157655 496966 157664
rect 496912 157344 496964 157350
rect 496912 157286 496964 157292
rect 496924 156505 496952 157286
rect 496910 156496 496966 156505
rect 496910 156431 496966 156440
rect 496912 155916 496964 155922
rect 496912 155858 496964 155864
rect 496924 155417 496952 155858
rect 496910 155408 496966 155417
rect 496910 155343 496966 155352
rect 497004 154556 497056 154562
rect 497004 154498 497056 154504
rect 496912 154488 496964 154494
rect 496912 154430 496964 154436
rect 496924 154329 496952 154430
rect 496910 154320 496966 154329
rect 496910 154255 496966 154264
rect 497016 153241 497044 154498
rect 497002 153232 497058 153241
rect 496912 153196 496964 153202
rect 497002 153167 497058 153176
rect 496912 153138 496964 153144
rect 496924 152153 496952 153138
rect 496910 152144 496966 152153
rect 496910 152079 496966 152088
rect 496818 150920 496874 150929
rect 496818 150855 496874 150864
rect 496820 150408 496872 150414
rect 496820 150350 496872 150356
rect 496832 149841 496860 150350
rect 496818 149832 496874 149841
rect 496818 149767 496874 149776
rect 496818 147656 496874 147665
rect 496818 147591 496820 147600
rect 496872 147591 496874 147600
rect 496820 147562 496872 147568
rect 496820 146260 496872 146266
rect 496820 146202 496872 146208
rect 496832 145353 496860 146202
rect 496818 145344 496874 145353
rect 496818 145279 496874 145288
rect 496818 144256 496874 144265
rect 496818 144191 496820 144200
rect 496872 144191 496874 144200
rect 496820 144162 496872 144168
rect 496820 143540 496872 143546
rect 496820 143482 496872 143488
rect 496832 143177 496860 143482
rect 496818 143168 496874 143177
rect 496818 143103 496874 143112
rect 496818 141944 496874 141953
rect 496818 141879 496874 141888
rect 496832 140894 496860 141879
rect 496820 140888 496872 140894
rect 496820 140830 496872 140836
rect 496820 140752 496872 140758
rect 496820 140694 496872 140700
rect 496832 139777 496860 140694
rect 496818 139768 496874 139777
rect 496818 139703 496874 139712
rect 496820 139392 496872 139398
rect 496820 139334 496872 139340
rect 496832 138689 496860 139334
rect 496818 138680 496874 138689
rect 496818 138615 496874 138624
rect 496820 137964 496872 137970
rect 496820 137906 496872 137912
rect 496832 137465 496860 137906
rect 496818 137456 496874 137465
rect 496818 137391 496874 137400
rect 496912 136604 496964 136610
rect 496912 136546 496964 136552
rect 496820 136400 496872 136406
rect 496818 136368 496820 136377
rect 496872 136368 496874 136377
rect 496818 136303 496874 136312
rect 496924 135289 496952 136546
rect 496910 135280 496966 135289
rect 496910 135215 496966 135224
rect 496820 133884 496872 133890
rect 496820 133826 496872 133832
rect 496832 132977 496860 133826
rect 496818 132968 496874 132977
rect 496818 132903 496874 132912
rect 497464 131164 497516 131170
rect 497464 131106 497516 131112
rect 495622 130792 495678 130801
rect 495622 130727 495678 130736
rect 496820 129736 496872 129742
rect 496818 129704 496820 129713
rect 496872 129704 496874 129713
rect 496818 129639 496874 129648
rect 496820 128308 496872 128314
rect 496820 128250 496872 128256
rect 496832 127401 496860 128250
rect 496818 127392 496874 127401
rect 496818 127327 496874 127336
rect 496912 127288 496964 127294
rect 496912 127230 496964 127236
rect 496820 126948 496872 126954
rect 496820 126890 496872 126896
rect 496832 126313 496860 126890
rect 496818 126304 496874 126313
rect 496818 126239 496874 126248
rect 496820 125588 496872 125594
rect 496820 125530 496872 125536
rect 496832 125225 496860 125530
rect 496818 125216 496874 125225
rect 496818 125151 496874 125160
rect 496924 124137 496952 127230
rect 496910 124128 496966 124137
rect 496820 124092 496872 124098
rect 496910 124063 496966 124072
rect 496820 124034 496872 124040
rect 496832 122913 496860 124034
rect 496818 122904 496874 122913
rect 496818 122839 496874 122848
rect 496820 122800 496872 122806
rect 496820 122742 496872 122748
rect 496832 121825 496860 122742
rect 496818 121816 496874 121825
rect 496818 121751 496874 121760
rect 496912 119604 496964 119610
rect 496912 119546 496964 119552
rect 496820 118652 496872 118658
rect 496820 118594 496872 118600
rect 496832 118425 496860 118594
rect 496818 118416 496874 118425
rect 496818 118351 496874 118360
rect 496924 117337 496952 119546
rect 496910 117328 496966 117337
rect 496820 117292 496872 117298
rect 496910 117263 496966 117272
rect 496820 117234 496872 117240
rect 496832 116249 496860 117234
rect 496818 116240 496874 116249
rect 496818 116175 496874 116184
rect 497476 115161 497504 131106
rect 497462 115152 497518 115161
rect 497462 115087 497518 115096
rect 496820 114232 496872 114238
rect 496820 114174 496872 114180
rect 496832 113937 496860 114174
rect 496818 113928 496874 113937
rect 496818 113863 496874 113872
rect 496910 112840 496966 112849
rect 496910 112775 496966 112784
rect 496820 111784 496872 111790
rect 496818 111752 496820 111761
rect 496872 111752 496874 111761
rect 496818 111687 496874 111696
rect 496820 111648 496872 111654
rect 496820 111590 496872 111596
rect 496832 110673 496860 111590
rect 496818 110664 496874 110673
rect 496818 110599 496874 110608
rect 496820 110424 496872 110430
rect 496820 110366 496872 110372
rect 496832 109449 496860 110366
rect 496818 109440 496874 109449
rect 496818 109375 496874 109384
rect 496820 107636 496872 107642
rect 496820 107578 496872 107584
rect 496832 107273 496860 107578
rect 496818 107264 496874 107273
rect 496818 107199 496874 107208
rect 496924 107114 496952 112775
rect 497002 108352 497058 108361
rect 497002 108287 497058 108296
rect 496832 107086 496952 107114
rect 496832 96626 496860 107086
rect 496910 106176 496966 106185
rect 496910 106111 496966 106120
rect 496924 99278 496952 106111
rect 496912 99272 496964 99278
rect 496912 99214 496964 99220
rect 497016 97918 497044 108287
rect 497094 101688 497150 101697
rect 497094 101623 497150 101632
rect 497004 97912 497056 97918
rect 497004 97854 497056 97860
rect 496820 96620 496872 96626
rect 496820 96562 496872 96568
rect 497108 92478 497136 101623
rect 497096 92472 497148 92478
rect 497096 92414 497148 92420
rect 498212 47598 498240 171142
rect 498304 131170 498332 237390
rect 498384 210520 498436 210526
rect 498384 210462 498436 210468
rect 498292 131164 498344 131170
rect 498292 131106 498344 131112
rect 498396 120737 498424 210462
rect 498476 175636 498528 175642
rect 498476 175578 498528 175584
rect 498382 120728 498438 120737
rect 498382 120663 498438 120672
rect 498488 95946 498516 175578
rect 499592 124098 499620 360159
rect 508504 354000 508556 354006
rect 508504 353942 508556 353948
rect 500960 313948 501012 313954
rect 500960 313890 501012 313896
rect 499672 291236 499724 291242
rect 499672 291178 499724 291184
rect 499580 124092 499632 124098
rect 499580 124034 499632 124040
rect 499684 114238 499712 291178
rect 499856 267028 499908 267034
rect 499856 266970 499908 266976
rect 499764 176724 499816 176730
rect 499764 176666 499816 176672
rect 499672 114232 499724 114238
rect 499672 114174 499724 114180
rect 498476 95940 498528 95946
rect 498476 95882 498528 95888
rect 498200 47592 498252 47598
rect 498200 47534 498252 47540
rect 499776 9654 499804 176666
rect 499868 127294 499896 266970
rect 499856 127288 499908 127294
rect 499856 127230 499908 127236
rect 500972 119610 501000 313890
rect 504364 312588 504416 312594
rect 504364 312530 504416 312536
rect 502432 240236 502484 240242
rect 502432 240178 502484 240184
rect 502340 196648 502392 196654
rect 502340 196590 502392 196596
rect 501144 189848 501196 189854
rect 501144 189790 501196 189796
rect 501052 176792 501104 176798
rect 501052 176734 501104 176740
rect 500960 119604 501012 119610
rect 500960 119546 501012 119552
rect 501064 15162 501092 176734
rect 501156 111654 501184 189790
rect 501236 180328 501288 180334
rect 501236 180270 501288 180276
rect 501248 136406 501276 180270
rect 501236 136400 501288 136406
rect 501236 136342 501288 136348
rect 501144 111648 501196 111654
rect 501144 111590 501196 111596
rect 502352 107642 502380 196590
rect 502444 168366 502472 240178
rect 504376 235958 504404 312530
rect 506480 287088 506532 287094
rect 506480 287030 506532 287036
rect 504364 235952 504416 235958
rect 504364 235894 504416 235900
rect 504376 235006 504404 235894
rect 503720 235000 503772 235006
rect 503720 234942 503772 234948
rect 504364 235000 504416 235006
rect 504364 234942 504416 234948
rect 502616 181552 502668 181558
rect 502616 181494 502668 181500
rect 502524 178696 502576 178702
rect 502524 178638 502576 178644
rect 502432 168360 502484 168366
rect 502432 168302 502484 168308
rect 502536 140758 502564 178638
rect 502628 154494 502656 181494
rect 503628 178696 503680 178702
rect 503628 178638 503680 178644
rect 503640 178090 503668 178638
rect 503628 178084 503680 178090
rect 503628 178026 503680 178032
rect 503628 168360 503680 168366
rect 503628 168302 503680 168308
rect 503640 167686 503668 168302
rect 503628 167680 503680 167686
rect 503628 167622 503680 167628
rect 503732 160002 503760 234942
rect 505100 206304 505152 206310
rect 505100 206246 505152 206252
rect 503904 185632 503956 185638
rect 503904 185574 503956 185580
rect 503812 180124 503864 180130
rect 503812 180066 503864 180072
rect 503720 159996 503772 160002
rect 503720 159938 503772 159944
rect 502616 154488 502668 154494
rect 502616 154430 502668 154436
rect 502800 140820 502852 140826
rect 502800 140762 502852 140768
rect 502524 140752 502576 140758
rect 502524 140694 502576 140700
rect 502812 140078 502840 140762
rect 502800 140072 502852 140078
rect 502800 140014 502852 140020
rect 503824 117298 503852 180066
rect 503916 150414 503944 185574
rect 503996 181620 504048 181626
rect 503996 181562 504048 181568
rect 504008 164898 504036 181562
rect 504086 166968 504142 166977
rect 504086 166903 504142 166912
rect 504100 166326 504128 166903
rect 504088 166320 504140 166326
rect 504088 166262 504140 166268
rect 504100 165646 504128 166262
rect 504088 165640 504140 165646
rect 504088 165582 504140 165588
rect 503996 164892 504048 164898
rect 503996 164834 504048 164840
rect 504008 161474 504036 164834
rect 504008 161446 504404 161474
rect 503904 150408 503956 150414
rect 503904 150350 503956 150356
rect 503812 117292 503864 117298
rect 503812 117234 503864 117240
rect 502340 107636 502392 107642
rect 502340 107578 502392 107584
rect 504376 86970 504404 161446
rect 505112 122806 505140 206246
rect 505192 184272 505244 184278
rect 505192 184214 505244 184220
rect 505204 147626 505232 184214
rect 505284 181688 505336 181694
rect 505284 181630 505336 181636
rect 505296 154562 505324 181630
rect 505284 154556 505336 154562
rect 505284 154498 505336 154504
rect 505192 147620 505244 147626
rect 505192 147562 505244 147568
rect 505100 122800 505152 122806
rect 505100 122742 505152 122748
rect 506492 111790 506520 287030
rect 507952 195288 508004 195294
rect 507952 195230 508004 195236
rect 507860 184204 507912 184210
rect 507860 184146 507912 184152
rect 506572 180260 506624 180266
rect 506572 180202 506624 180208
rect 506584 144498 506612 180202
rect 506572 144492 506624 144498
rect 506572 144434 506624 144440
rect 507124 144492 507176 144498
rect 507124 144434 507176 144440
rect 506584 144226 506612 144434
rect 506572 144220 506624 144226
rect 506572 144162 506624 144168
rect 506480 111784 506532 111790
rect 506480 111726 506532 111732
rect 504364 86964 504416 86970
rect 504364 86906 504416 86912
rect 507136 20670 507164 144434
rect 507872 128314 507900 184146
rect 507964 153202 507992 195230
rect 507952 153196 508004 153202
rect 507952 153138 508004 153144
rect 508516 136610 508544 353942
rect 509332 200796 509384 200802
rect 509332 200738 509384 200744
rect 509240 180192 509292 180198
rect 509240 180134 509292 180140
rect 508504 136604 508556 136610
rect 508504 136546 508556 136552
rect 509252 129742 509280 180134
rect 509344 164218 509372 200738
rect 509332 164212 509384 164218
rect 509332 164154 509384 164160
rect 509240 129736 509292 129742
rect 509240 129678 509292 129684
rect 507860 128308 507912 128314
rect 507860 128250 507912 128256
rect 510632 110430 510660 362918
rect 512092 239420 512144 239426
rect 512092 239362 512144 239368
rect 512104 238814 512132 239362
rect 512092 238808 512144 238814
rect 512092 238750 512144 238756
rect 510712 221468 510764 221474
rect 510712 221410 510764 221416
rect 510724 143546 510752 221410
rect 511998 211848 512054 211857
rect 511998 211783 512054 211792
rect 510804 184340 510856 184346
rect 510804 184282 510856 184288
rect 510816 146266 510844 184282
rect 510804 146260 510856 146266
rect 510804 146202 510856 146208
rect 510712 143540 510764 143546
rect 510712 143482 510764 143488
rect 512012 133890 512040 211783
rect 512104 161430 512132 238750
rect 517610 218648 517666 218657
rect 517610 218583 517666 218592
rect 514760 207664 514812 207670
rect 514760 207606 514812 207612
rect 514772 206310 514800 207606
rect 514760 206304 514812 206310
rect 514760 206246 514812 206252
rect 515404 206304 515456 206310
rect 515404 206246 515456 206252
rect 514760 199436 514812 199442
rect 514760 199378 514812 199384
rect 513380 186992 513432 186998
rect 513380 186934 513432 186940
rect 512092 161424 512144 161430
rect 512092 161366 512144 161372
rect 512644 143540 512696 143546
rect 512644 143482 512696 143488
rect 512000 133884 512052 133890
rect 512000 133826 512052 133832
rect 510620 110424 510672 110430
rect 510620 110366 510672 110372
rect 512656 60722 512684 143482
rect 513392 125594 513420 186934
rect 514772 126954 514800 199378
rect 515416 162858 515444 206246
rect 517520 192500 517572 192506
rect 517520 192442 517572 192448
rect 515404 162852 515456 162858
rect 515404 162794 515456 162800
rect 514760 126948 514812 126954
rect 514760 126890 514812 126896
rect 513380 125588 513432 125594
rect 513380 125530 513432 125536
rect 517532 118658 517560 192442
rect 517624 158710 517652 218583
rect 517612 158704 517664 158710
rect 517612 158646 517664 158652
rect 519556 155922 519584 700946
rect 521580 700330 521608 700946
rect 550560 700330 550588 702510
rect 521568 700324 521620 700330
rect 521568 700266 521620 700272
rect 550548 700324 550600 700330
rect 550548 700266 550600 700272
rect 580920 697241 580948 702578
rect 580906 697232 580962 697241
rect 580906 697167 580962 697176
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580264 680400 580316 680406
rect 580264 680342 580316 680348
rect 580276 670721 580304 680342
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 582378 670712 582434 670721
rect 582378 670647 582434 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 579804 634840 579856 634846
rect 579804 634782 579856 634788
rect 579816 630873 579844 634782
rect 579802 630864 579858 630873
rect 579802 630799 579858 630808
rect 580172 618248 580224 618254
rect 580172 618190 580224 618196
rect 580184 617545 580212 618190
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580262 588024 580318 588033
rect 580262 587959 580318 587968
rect 580276 577697 580304 587959
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 580170 564360 580226 564369
rect 580170 564295 580226 564304
rect 580184 563718 580212 564295
rect 580172 563712 580224 563718
rect 580172 563654 580224 563660
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 431254 580212 431559
rect 580172 431248 580224 431254
rect 580172 431190 580224 431196
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 544384 404388 544436 404394
rect 544384 404330 544436 404336
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 520924 376780 520976 376786
rect 520924 376722 520976 376728
rect 520936 218754 520964 376722
rect 521660 276072 521712 276078
rect 521660 276014 521712 276020
rect 520924 218748 520976 218754
rect 520924 218690 520976 218696
rect 519544 155916 519596 155922
rect 519544 155858 519596 155864
rect 520188 140888 520240 140894
rect 520188 140830 520240 140836
rect 517520 118652 517572 118658
rect 517520 118594 517572 118600
rect 520200 100706 520228 140830
rect 520936 139398 520964 218690
rect 521672 140894 521700 276014
rect 536840 240780 536892 240786
rect 536840 240722 536892 240728
rect 536852 240174 536880 240722
rect 536840 240168 536892 240174
rect 536840 240110 536892 240116
rect 525064 165640 525116 165646
rect 525064 165582 525116 165588
rect 535460 165640 535512 165646
rect 535460 165582 535512 165588
rect 521660 140888 521712 140894
rect 521660 140830 521712 140836
rect 520924 139392 520976 139398
rect 520924 139334 520976 139340
rect 520188 100700 520240 100706
rect 520188 100642 520240 100648
rect 512644 60716 512696 60722
rect 512644 60658 512696 60664
rect 525076 46918 525104 165582
rect 530584 164280 530636 164286
rect 530584 164222 530636 164228
rect 530596 127634 530624 164222
rect 535472 164218 535500 165582
rect 535460 164212 535512 164218
rect 535460 164154 535512 164160
rect 536852 160070 536880 240110
rect 543004 167680 543056 167686
rect 543004 167622 543056 167628
rect 536840 160064 536892 160070
rect 536840 160006 536892 160012
rect 530584 127628 530636 127634
rect 530584 127570 530636 127576
rect 525064 46912 525116 46918
rect 525064 46854 525116 46860
rect 507124 20664 507176 20670
rect 507124 20606 507176 20612
rect 501052 15156 501104 15162
rect 501052 15098 501104 15104
rect 499764 9648 499816 9654
rect 499764 9590 499816 9596
rect 543016 6866 543044 167622
rect 544396 158710 544424 404330
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 579632 354006 579660 364346
rect 579620 354000 579672 354006
rect 579620 353942 579672 353948
rect 580262 351928 580318 351937
rect 580262 351863 580318 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580276 312594 580304 351863
rect 580264 312588 580316 312594
rect 580264 312530 580316 312536
rect 580354 312080 580410 312089
rect 580354 312015 580410 312024
rect 580368 300150 580396 312015
rect 580356 300144 580408 300150
rect 580356 300086 580408 300092
rect 580262 298752 580318 298761
rect 580262 298687 580318 298696
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 548524 260160 548576 260166
rect 548524 260102 548576 260108
rect 548536 258738 548564 260102
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258738 580028 258839
rect 548524 258732 548576 258738
rect 548524 258674 548576 258680
rect 579988 258732 580040 258738
rect 579988 258674 580040 258680
rect 544384 158704 544436 158710
rect 544384 158646 544436 158652
rect 548536 137970 548564 258674
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 239426 580212 245511
rect 580276 240786 580304 298687
rect 580264 240780 580316 240786
rect 580264 240722 580316 240728
rect 580172 239420 580224 239426
rect 580172 239362 580224 239368
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580184 231878 580212 232319
rect 580172 231872 580224 231878
rect 580172 231814 580224 231820
rect 579802 219056 579858 219065
rect 579802 218991 579858 219000
rect 579816 218754 579844 218991
rect 579804 218748 579856 218754
rect 579804 218690 579856 218696
rect 580172 206304 580224 206310
rect 580172 206246 580224 206252
rect 580184 205737 580212 206246
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 580368 182850 580396 192471
rect 580356 182844 580408 182850
rect 580356 182786 580408 182792
rect 580264 182232 580316 182238
rect 580264 182174 580316 182180
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580184 178090 580212 179143
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580276 152697 580304 182174
rect 582392 157350 582420 670647
rect 582380 157344 582432 157350
rect 582380 157286 582432 157292
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580172 140072 580224 140078
rect 580172 140014 580224 140020
rect 580184 139369 580212 140014
rect 580170 139360 580226 139369
rect 580170 139295 580226 139304
rect 548524 137964 548576 137970
rect 548524 137906 548576 137912
rect 580172 127628 580224 127634
rect 580172 127570 580224 127576
rect 580184 126041 580212 127570
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580262 112840 580318 112849
rect 580262 112775 580318 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580276 99346 580304 112775
rect 580264 99340 580316 99346
rect 580264 99282 580316 99288
rect 580264 93152 580316 93158
rect 580264 93094 580316 93100
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580276 33153 580304 93094
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 543004 6860 543056 6866
rect 543004 6802 543056 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 351184 3936 351236 3942
rect 351184 3878 351236 3884
rect 351644 3936 351696 3942
rect 351644 3878 351696 3884
rect 495532 3936 495584 3942
rect 495532 3878 495584 3884
rect 351656 480 351684 3878
rect 345726 354 345838 480
rect 345308 326 345838 354
rect 345726 -960 345838 326
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 2778 658180 2780 658200
rect 2780 658180 2832 658200
rect 2832 658180 2834 658200
rect 2778 658144 2834 658180
rect 4066 632032 4122 632088
rect 3514 619112 3570 619168
rect 3422 606056 3478 606112
rect 3422 579944 3478 580000
rect 3238 566888 3294 566944
rect 3330 553832 3386 553888
rect 3146 527856 3202 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3146 501744 3202 501800
rect 3422 475632 3478 475688
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3146 449520 3202 449576
rect 30286 468424 30342 468480
rect 3514 423544 3570 423600
rect 3422 410488 3478 410544
rect 3422 397432 3478 397488
rect 3146 358400 3202 358456
rect 2778 345344 2834 345400
rect 3514 371320 3570 371376
rect 30286 352552 30342 352608
rect 3422 319232 3478 319288
rect 3422 306176 3478 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 3422 241032 3478 241088
rect 1306 224168 1362 224224
rect 3330 214920 3386 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 3238 162832 3294 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 110608 3478 110664
rect 2778 97552 2834 97608
rect 3146 84632 3202 84688
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3514 32408 3570 32464
rect 3422 19352 3478 19408
rect 11058 76472 11114 76528
rect 3422 6432 3478 6488
rect 8206 16496 8262 16552
rect 33782 549208 33838 549264
rect 35714 586336 35770 586392
rect 34426 549208 34482 549264
rect 35622 447752 35678 447808
rect 37094 546352 37150 546408
rect 37186 525680 37242 525736
rect 38382 445576 38438 445632
rect 41326 586744 41382 586800
rect 41142 448432 41198 448488
rect 41142 447752 41198 447808
rect 43810 585384 43866 585440
rect 43718 568520 43774 568576
rect 42614 459448 42670 459504
rect 45190 588104 45246 588160
rect 46570 586608 46626 586664
rect 47950 585520 48006 585576
rect 49330 534112 49386 534168
rect 48962 489776 49018 489832
rect 48962 402192 49018 402248
rect 52182 583888 52238 583944
rect 50802 438776 50858 438832
rect 50986 438776 51042 438832
rect 53562 583752 53618 583808
rect 52366 539436 52422 539472
rect 52366 539416 52368 539436
rect 52368 539416 52420 539436
rect 52420 539416 52422 539436
rect 52182 488552 52238 488608
rect 50986 390768 51042 390824
rect 49606 298832 49662 298888
rect 54850 585248 54906 585304
rect 55034 533568 55090 533624
rect 56414 542952 56470 543008
rect 53746 387932 53802 387968
rect 53746 387912 53748 387932
rect 53748 387912 53800 387932
rect 53800 387912 53802 387932
rect 49606 210296 49662 210352
rect 53562 300056 53618 300112
rect 57610 553424 57666 553480
rect 45558 61512 45614 61568
rect 44270 12960 44326 13016
rect 57794 538056 57850 538112
rect 57886 533840 57942 533896
rect 58990 462168 59046 462224
rect 56230 308352 56286 308408
rect 56230 235184 56286 235240
rect 57794 339360 57850 339416
rect 60554 584024 60610 584080
rect 59358 379480 59414 379536
rect 57794 278840 57850 278896
rect 57518 192480 57574 192536
rect 57794 93744 57850 93800
rect 60738 546352 60794 546408
rect 60738 542988 60740 543008
rect 60740 542988 60792 543008
rect 60792 542988 60794 543008
rect 60738 542952 60794 542988
rect 67546 679088 67602 679144
rect 61382 538736 61438 538792
rect 61382 463528 61438 463584
rect 61382 462304 61438 462360
rect 60554 367104 60610 367160
rect 60462 356632 60518 356688
rect 61842 447208 61898 447264
rect 61382 366968 61438 367024
rect 59358 57160 59414 57216
rect 63038 477556 63094 477592
rect 63038 477536 63040 477556
rect 63040 477536 63092 477556
rect 63092 477536 63094 477556
rect 63130 445984 63186 446040
rect 67454 675688 67510 675744
rect 64694 578176 64750 578232
rect 64234 468424 64290 468480
rect 64234 467916 64236 467936
rect 64236 467916 64288 467936
rect 64288 467916 64290 467936
rect 64234 467880 64290 467916
rect 63222 237224 63278 237280
rect 64510 364384 64566 364440
rect 66074 573960 66130 574016
rect 65982 546080 66038 546136
rect 64786 401668 64842 401704
rect 64786 401648 64788 401668
rect 64788 401648 64840 401668
rect 64840 401648 64842 401668
rect 67638 678136 67694 678192
rect 67638 676368 67694 676424
rect 67638 675144 67694 675200
rect 67638 674328 67694 674384
rect 67730 673784 67786 673840
rect 68742 677048 68798 677104
rect 68650 671744 68706 671800
rect 67638 670928 67694 670984
rect 67638 670248 67694 670304
rect 67730 669568 67786 669624
rect 67822 669296 67878 669352
rect 67822 668208 67878 668264
rect 67638 666848 67694 666904
rect 67730 665488 67786 665544
rect 67638 665236 67694 665272
rect 67638 665216 67640 665236
rect 67640 665216 67692 665236
rect 67692 665216 67694 665236
rect 67730 664128 67786 664184
rect 67638 663876 67694 663912
rect 67638 663856 67640 663876
rect 67640 663856 67692 663876
rect 67692 663856 67694 663876
rect 67638 662904 67694 662960
rect 67638 661408 67694 661464
rect 67730 660048 67786 660104
rect 67638 659640 67694 659696
rect 68558 658824 68614 658880
rect 67638 658688 67694 658744
rect 67730 657328 67786 657384
rect 68190 656648 68246 656704
rect 67638 655968 67694 656024
rect 67638 654780 67640 654800
rect 67640 654780 67692 654800
rect 67692 654780 67694 654800
rect 67638 654744 67694 654780
rect 67730 653248 67786 653304
rect 67914 652704 67970 652760
rect 67638 651888 67694 651944
rect 67638 650020 67640 650040
rect 67640 650020 67692 650040
rect 67692 650020 67694 650040
rect 67638 649984 67694 650020
rect 67638 649168 67694 649224
rect 67730 647808 67786 647864
rect 67638 647284 67694 647320
rect 67638 647264 67640 647284
rect 67640 647264 67692 647284
rect 67692 647264 67694 647284
rect 67638 646448 67694 646504
rect 68558 643728 68614 643784
rect 67730 642368 67786 642424
rect 67638 641824 67694 641880
rect 67730 641008 67786 641064
rect 67638 640464 67694 640520
rect 67638 579264 67694 579320
rect 67730 578176 67786 578232
rect 67454 575184 67510 575240
rect 67638 577768 67694 577824
rect 67730 577224 67786 577280
rect 67638 575728 67694 575784
rect 67638 574504 67694 574560
rect 67730 573960 67786 574016
rect 67638 573824 67694 573880
rect 67730 573280 67786 573336
rect 67638 571648 67694 571704
rect 67638 570968 67694 571024
rect 67730 570288 67786 570344
rect 67638 569064 67694 569120
rect 67822 568948 67878 568984
rect 67822 568928 67824 568948
rect 67824 568928 67876 568948
rect 67876 568928 67878 568948
rect 67638 568268 67694 568304
rect 67638 568248 67640 568268
rect 67640 568248 67692 568268
rect 67692 568248 67694 568268
rect 67638 567704 67694 567760
rect 67638 566344 67694 566400
rect 67638 564984 67694 565040
rect 67638 564848 67694 564904
rect 67638 564168 67694 564224
rect 67730 563624 67786 563680
rect 67638 562300 67640 562320
rect 67640 562300 67692 562320
rect 67692 562300 67694 562320
rect 67638 562264 67694 562300
rect 67638 561448 67694 561504
rect 67730 560904 67786 560960
rect 67638 559544 67694 559600
rect 67730 558048 67786 558104
rect 67638 557504 67694 557560
rect 67822 557368 67878 557424
rect 67638 556824 67694 556880
rect 67638 555328 67694 555384
rect 67730 554784 67786 554840
rect 67914 554648 67970 554704
rect 67638 554104 67694 554160
rect 67638 552644 67640 552664
rect 67640 552644 67692 552664
rect 67692 552644 67694 552664
rect 67638 552608 67694 552644
rect 67638 551964 67640 551984
rect 67640 551964 67692 551984
rect 67692 551964 67694 551984
rect 67638 551928 67694 551964
rect 67638 549344 67694 549400
rect 67730 549208 67786 549264
rect 67638 548564 67640 548584
rect 67640 548564 67692 548584
rect 67692 548564 67694 548584
rect 67638 548528 67694 548564
rect 67638 547168 67694 547224
rect 67638 546508 67694 546544
rect 67638 546488 67640 546508
rect 67640 546488 67692 546508
rect 67692 546488 67694 546508
rect 67638 545148 67694 545184
rect 67638 545128 67640 545148
rect 67640 545128 67692 545148
rect 67692 545128 67694 545148
rect 68926 654744 68982 654800
rect 68834 651344 68890 651400
rect 68650 576544 68706 576600
rect 68190 543768 68246 543824
rect 68558 543768 68614 543824
rect 67638 543224 67694 543280
rect 67730 543088 67786 543144
rect 67638 541184 67694 541240
rect 67638 540504 67694 540560
rect 67730 489096 67786 489152
rect 67638 488008 67694 488064
rect 67638 487872 67694 487928
rect 67730 486512 67786 486568
rect 67638 485852 67694 485888
rect 67638 485832 67640 485852
rect 67640 485832 67692 485852
rect 67692 485832 67694 485852
rect 67638 485152 67694 485208
rect 67638 483928 67694 483984
rect 68006 482432 68062 482488
rect 68098 481480 68154 481536
rect 67638 481072 67694 481128
rect 68098 480528 68154 480584
rect 67638 479712 67694 479768
rect 67546 479168 67602 479224
rect 67638 478216 67694 478272
rect 67638 476448 67694 476504
rect 67638 475632 67694 475688
rect 66166 404368 66222 404424
rect 67454 466792 67510 466848
rect 67362 453328 67418 453384
rect 67730 474952 67786 475008
rect 67638 472640 67694 472696
rect 67730 471044 67732 471064
rect 67732 471044 67784 471064
rect 67784 471044 67786 471064
rect 67730 471008 67786 471044
rect 67638 470212 67694 470248
rect 67638 470192 67640 470212
rect 67640 470192 67692 470212
rect 67692 470192 67694 470212
rect 67730 469648 67786 469704
rect 67638 468832 67694 468888
rect 67638 468152 67694 468208
rect 67730 466112 67786 466168
rect 67638 465568 67694 465624
rect 67638 464752 67694 464808
rect 67730 464208 67786 464264
rect 67638 462712 67694 462768
rect 67638 460164 67640 460184
rect 67640 460164 67692 460184
rect 67692 460164 67694 460184
rect 67638 460128 67694 460164
rect 67730 459312 67786 459368
rect 67638 458768 67694 458824
rect 67638 457444 67640 457464
rect 67640 457444 67692 457464
rect 67692 457444 67694 457464
rect 67638 457408 67694 457444
rect 67638 457272 67694 457328
rect 67730 456184 67786 456240
rect 67638 454552 67694 454608
rect 68006 454028 68062 454064
rect 68006 454008 68008 454028
rect 68008 454008 68060 454028
rect 68060 454008 68062 454028
rect 67638 453192 67694 453248
rect 67638 452548 67640 452568
rect 67640 452548 67692 452568
rect 67692 452548 67694 452568
rect 67638 452512 67694 452548
rect 67638 450744 67694 450800
rect 67730 449112 67786 449168
rect 67638 448468 67640 448488
rect 67640 448468 67692 448488
rect 67692 448468 67694 448488
rect 67638 448432 67694 448468
rect 67638 447208 67694 447264
rect 67638 446392 67694 446448
rect 68466 484608 68522 484664
rect 68926 644544 68982 644600
rect 68650 476992 68706 477048
rect 68190 444216 68246 444272
rect 67638 443808 67694 443864
rect 67730 442448 67786 442504
rect 67638 442312 67694 442368
rect 67638 441088 67694 441144
rect 67638 440952 67694 441008
rect 67638 384784 67694 384840
rect 67638 382472 67694 382528
rect 67638 380840 67694 380896
rect 67546 380296 67602 380352
rect 67914 380704 67970 380760
rect 67638 379888 67694 379944
rect 67638 377032 67694 377088
rect 67638 375536 67694 375592
rect 67638 374620 67640 374640
rect 67640 374620 67692 374640
rect 67692 374620 67694 374640
rect 67638 374584 67694 374620
rect 67730 374448 67786 374504
rect 67730 373224 67786 373280
rect 67638 372408 67694 372464
rect 67454 371728 67510 371784
rect 67638 370368 67694 370424
rect 67638 369688 67694 369744
rect 67638 368500 67640 368520
rect 67640 368500 67692 368520
rect 67692 368500 67694 368520
rect 67638 368464 67694 368500
rect 67638 367004 67640 367024
rect 67640 367004 67692 367024
rect 67692 367004 67694 367024
rect 67638 366968 67694 367004
rect 68834 551384 68890 551440
rect 70398 679768 70454 679824
rect 74538 681808 74594 681864
rect 75182 680448 75238 680504
rect 77114 680312 77170 680368
rect 79322 680448 79378 680504
rect 89166 699760 89222 699816
rect 89074 680584 89130 680640
rect 84842 680448 84898 680504
rect 81622 680312 81678 680368
rect 82082 680312 82138 680368
rect 85486 680312 85542 680368
rect 89718 680448 89774 680504
rect 98550 681808 98606 681864
rect 99286 681808 99342 681864
rect 91926 680312 91982 680368
rect 94870 679632 94926 679688
rect 96802 679632 96858 679688
rect 81898 679496 81954 679552
rect 85762 679496 85818 679552
rect 92938 679496 92994 679552
rect 96158 679496 96214 679552
rect 106922 681808 106978 681864
rect 107566 681808 107622 681864
rect 102506 680448 102562 680504
rect 104806 680312 104862 680368
rect 100666 679632 100722 679688
rect 99378 679496 99434 679552
rect 71778 679360 71834 679416
rect 73618 679360 73674 679416
rect 75458 679360 75514 679416
rect 76194 679360 76250 679416
rect 78126 679360 78182 679416
rect 78862 679360 78918 679416
rect 80150 679360 80206 679416
rect 82726 679360 82782 679416
rect 84474 679360 84530 679416
rect 86498 679360 86554 679416
rect 87142 679360 87198 679416
rect 87786 679360 87842 679416
rect 91466 679360 91522 679416
rect 92754 679360 92810 679416
rect 94226 679360 94282 679416
rect 96158 679360 96214 679416
rect 97354 679360 97410 679416
rect 98550 679360 98606 679416
rect 100022 679360 100078 679416
rect 101310 679360 101366 679416
rect 103334 679768 103390 679824
rect 107658 680448 107714 680504
rect 108394 679632 108450 679688
rect 105818 679496 105874 679552
rect 106922 679496 106978 679552
rect 102598 679360 102654 679416
rect 105634 679360 105690 679416
rect 107106 679360 107162 679416
rect 69202 643184 69258 643240
rect 68834 544448 68890 544504
rect 110418 672560 110474 672616
rect 70766 586336 70822 586392
rect 70398 585112 70454 585168
rect 70214 581168 70270 581224
rect 69294 580624 69350 580680
rect 69662 580624 69718 580680
rect 69846 544312 69902 544368
rect 70398 581168 70454 581224
rect 71962 585520 72018 585576
rect 70950 584024 71006 584080
rect 72238 584024 72294 584080
rect 73342 586744 73398 586800
rect 73342 586336 73398 586392
rect 72698 585520 72754 585576
rect 77390 638832 77446 638888
rect 75734 589192 75790 589248
rect 74630 583888 74686 583944
rect 75274 583752 75330 583808
rect 75642 583752 75698 583808
rect 76746 587832 76802 587888
rect 76010 585384 76066 585440
rect 80978 639784 81034 639840
rect 77482 624416 77538 624472
rect 79966 589192 80022 589248
rect 78678 587696 78734 587752
rect 78678 586608 78734 586664
rect 78218 585112 78274 585168
rect 81438 638832 81494 638888
rect 84290 638832 84346 638888
rect 85578 629856 85634 629912
rect 86958 629856 87014 629912
rect 92386 638832 92442 638888
rect 89350 627136 89406 627192
rect 89626 593408 89682 593464
rect 88246 588512 88302 588568
rect 84290 588240 84346 588296
rect 84106 586472 84162 586528
rect 83278 582392 83334 582448
rect 81898 581984 81954 582040
rect 84014 583752 84070 583808
rect 84014 582392 84070 582448
rect 85394 585384 85450 585440
rect 85118 585112 85174 585168
rect 86222 583752 86278 583808
rect 88890 585112 88946 585168
rect 91006 593272 91062 593328
rect 90270 585112 90326 585168
rect 95882 639648 95938 639704
rect 95146 638696 95202 638752
rect 100298 638832 100354 638888
rect 91098 589328 91154 589384
rect 92386 589328 92442 589384
rect 96434 590008 96490 590064
rect 94962 587152 95018 587208
rect 93766 583752 93822 583808
rect 94134 582528 94190 582584
rect 97262 589872 97318 589928
rect 96526 589192 96582 589248
rect 97170 587832 97226 587888
rect 97078 585112 97134 585168
rect 98734 586336 98790 586392
rect 99102 584024 99158 584080
rect 99102 583752 99158 583808
rect 101310 585520 101366 585576
rect 100574 581848 100630 581904
rect 103426 638832 103482 638888
rect 103150 587424 103206 587480
rect 105450 637608 105506 637664
rect 107382 638560 107438 638616
rect 105542 585520 105598 585576
rect 104622 584024 104678 584080
rect 104438 583888 104494 583944
rect 106094 578176 106150 578232
rect 105634 574368 105690 574424
rect 68926 482568 68982 482624
rect 69110 482568 69166 482624
rect 69018 482432 69074 482488
rect 69202 480528 69258 480584
rect 68926 473728 68982 473784
rect 68926 473320 68982 473376
rect 68742 451832 68798 451888
rect 68742 383424 68798 383480
rect 67638 364284 67640 364304
rect 67640 364284 67692 364304
rect 67692 364284 67694 364304
rect 67638 364248 67694 364284
rect 67638 362616 67694 362672
rect 67638 360712 67694 360768
rect 67730 360168 67786 360224
rect 67638 359624 67694 359680
rect 67546 358128 67602 358184
rect 67638 358028 67640 358048
rect 67640 358028 67692 358048
rect 67692 358028 67694 358048
rect 67638 357992 67694 358028
rect 66166 347692 66168 347712
rect 66168 347692 66220 347712
rect 66220 347692 66222 347712
rect 66166 347656 66222 347692
rect 68006 356904 68062 356960
rect 67730 355544 67786 355600
rect 67638 355136 67694 355192
rect 67546 353776 67602 353832
rect 67638 351736 67694 351792
rect 67638 349172 67694 349208
rect 67638 349152 67640 349172
rect 67640 349152 67692 349172
rect 67692 349152 67694 349172
rect 67638 349036 67694 349072
rect 67638 349016 67640 349036
rect 67640 349016 67692 349036
rect 67692 349016 67694 349036
rect 67638 347692 67640 347712
rect 67640 347692 67692 347712
rect 67692 347692 67694 347712
rect 67638 347656 67694 347692
rect 68926 445440 68982 445496
rect 74538 537376 74594 537432
rect 70858 492768 70914 492824
rect 81622 538056 81678 538112
rect 76470 494672 76526 494728
rect 74998 492768 75054 492824
rect 79690 492768 79746 492824
rect 83462 496032 83518 496088
rect 86958 531936 87014 531992
rect 86222 498752 86278 498808
rect 84842 497392 84898 497448
rect 91926 536696 91982 536752
rect 93674 532072 93730 532128
rect 87372 490048 87428 490104
rect 94042 538736 94098 538792
rect 97814 533296 97870 533352
rect 95054 491444 95056 491464
rect 95056 491444 95108 491464
rect 95108 491444 95110 491464
rect 95054 491408 95110 491444
rect 94134 489912 94190 489968
rect 95790 493312 95846 493368
rect 97078 491272 97134 491328
rect 99194 532208 99250 532264
rect 99654 538056 99710 538112
rect 99378 536696 99434 536752
rect 99470 446528 99526 446584
rect 99654 443808 99710 443864
rect 99746 443672 99802 443728
rect 99378 442312 99434 442368
rect 69202 439048 69258 439104
rect 71042 439048 71098 439104
rect 69110 380296 69166 380352
rect 68926 353096 68982 353152
rect 68926 347248 68982 347304
rect 68834 346332 68836 346352
rect 68836 346332 68888 346352
rect 68888 346332 68890 346352
rect 68834 346296 68890 346332
rect 68650 344936 68706 344992
rect 67638 343712 67694 343768
rect 67638 342896 67694 342952
rect 67454 298832 67510 298888
rect 67454 298288 67510 298344
rect 67454 283328 67510 283384
rect 67454 271904 67510 271960
rect 67362 261568 67418 261624
rect 67362 248648 67418 248704
rect 66074 225528 66130 225584
rect 67454 129240 67510 129296
rect 65522 128016 65578 128072
rect 66166 125160 66222 125216
rect 66074 123528 66130 123584
rect 65154 120808 65210 120864
rect 65982 102312 66038 102368
rect 67362 122576 67418 122632
rect 66074 100680 66130 100736
rect 67454 94832 67510 94888
rect 66074 88168 66130 88224
rect 67914 341672 67970 341728
rect 68742 341672 68798 341728
rect 67638 340992 67694 341048
rect 67638 340176 67694 340232
rect 68926 339904 68982 339960
rect 69202 363296 69258 363352
rect 71686 405728 71742 405784
rect 71962 438776 72018 438832
rect 74630 407496 74686 407552
rect 77298 437280 77354 437336
rect 77758 437280 77814 437336
rect 75182 407496 75238 407552
rect 75182 407088 75238 407144
rect 78862 437416 78918 437472
rect 79690 437416 79746 437472
rect 78862 389816 78918 389872
rect 84198 438912 84254 438968
rect 85486 438912 85542 438968
rect 84290 435920 84346 435976
rect 84842 435920 84898 435976
rect 83002 393896 83058 393952
rect 87602 437452 87604 437472
rect 87604 437452 87656 437472
rect 87656 437452 87658 437472
rect 87602 437416 87658 437452
rect 86222 437280 86278 437336
rect 85670 401648 85726 401704
rect 84934 390632 84990 390688
rect 88246 402192 88302 402248
rect 92570 438640 92626 438696
rect 92386 404912 92442 404968
rect 70950 385600 71006 385656
rect 97722 439864 97778 439920
rect 95146 393896 95202 393952
rect 98366 437824 98422 437880
rect 99470 441088 99526 441144
rect 99286 437824 99342 437880
rect 99286 407768 99342 407824
rect 98642 400832 98698 400888
rect 97998 397432 98054 397488
rect 101310 458088 101366 458144
rect 101126 400288 101182 400344
rect 100022 388320 100078 388376
rect 101954 470192 102010 470248
rect 101586 451152 101642 451208
rect 102414 485288 102470 485344
rect 102138 485172 102194 485208
rect 102138 485152 102140 485172
rect 102140 485152 102192 485172
rect 102192 485152 102194 485172
rect 102138 482568 102194 482624
rect 102782 487192 102838 487248
rect 102138 481072 102194 481128
rect 102230 480528 102286 480584
rect 102138 479848 102194 479904
rect 102138 476992 102194 477048
rect 102322 477128 102378 477184
rect 102230 476448 102286 476504
rect 102138 475632 102194 475688
rect 102138 474952 102194 475008
rect 102230 474272 102286 474328
rect 102138 472912 102194 472968
rect 102138 472232 102194 472288
rect 102138 471552 102194 471608
rect 102138 470872 102194 470928
rect 102138 469512 102194 469568
rect 102138 468832 102194 468888
rect 102138 467472 102194 467528
rect 102230 466928 102286 466984
rect 102230 466112 102286 466168
rect 102322 464888 102378 464944
rect 102138 464208 102194 464264
rect 102138 463392 102194 463448
rect 102138 462032 102194 462088
rect 102230 461488 102286 461544
rect 102138 460672 102194 460728
rect 102138 459992 102194 460048
rect 104806 539824 104862 539880
rect 104162 536832 104218 536888
rect 103426 488572 103482 488608
rect 103426 488552 103428 488572
rect 103428 488552 103480 488572
rect 103480 488552 103482 488572
rect 103426 487872 103482 487928
rect 103334 487328 103390 487384
rect 103334 486512 103390 486568
rect 103426 477672 103482 477728
rect 102138 459312 102194 459368
rect 102230 458768 102286 458824
rect 102874 456068 102930 456104
rect 102874 456048 102876 456068
rect 102876 456048 102928 456068
rect 102928 456048 102930 456068
rect 102230 455368 102286 455424
rect 102138 454688 102194 454744
rect 102874 453348 102930 453384
rect 102874 453328 102876 453348
rect 102876 453328 102928 453348
rect 102928 453328 102930 453348
rect 102138 453192 102194 453248
rect 102322 451968 102378 452024
rect 102138 450608 102194 450664
rect 102874 449268 102930 449304
rect 102874 449248 102876 449268
rect 102876 449248 102928 449268
rect 102928 449248 102930 449268
rect 102138 449112 102194 449168
rect 102230 448432 102286 448488
rect 102138 447888 102194 447944
rect 102598 446528 102654 446584
rect 102506 445712 102562 445768
rect 103242 445168 103298 445224
rect 102230 443672 102286 443728
rect 102874 442992 102930 443048
rect 102046 441632 102102 441688
rect 102598 441088 102654 441144
rect 102046 439728 102102 439784
rect 102230 395256 102286 395312
rect 104070 465568 104126 465624
rect 103610 455912 103666 455968
rect 105450 538056 105506 538112
rect 104806 536832 104862 536888
rect 103426 391176 103482 391232
rect 105542 479032 105598 479088
rect 105818 539552 105874 539608
rect 106922 587832 106978 587888
rect 107566 582664 107622 582720
rect 107014 577632 107070 577688
rect 106922 575048 106978 575104
rect 108026 580216 108082 580272
rect 108670 578720 108726 578776
rect 108118 578196 108174 578232
rect 108118 578176 108120 578196
rect 108120 578176 108172 578196
rect 108172 578176 108174 578196
rect 108946 580916 109002 580952
rect 108946 580896 108948 580916
rect 108948 580896 109000 580916
rect 109000 580896 109002 580916
rect 108946 579572 108948 579592
rect 108948 579572 109000 579592
rect 109000 579572 109002 579592
rect 108946 579536 109002 579572
rect 108946 577516 109002 577552
rect 108946 577496 108948 577516
rect 108948 577496 109000 577516
rect 109000 577496 109002 577516
rect 108762 576680 108818 576736
rect 108670 576172 108672 576192
rect 108672 576172 108724 576192
rect 108724 576172 108726 576192
rect 108670 576136 108726 576172
rect 107106 574640 107162 574696
rect 108946 573980 109002 574016
rect 108946 573960 108948 573980
rect 108948 573960 109000 573980
rect 109000 573960 109002 573980
rect 108946 573280 109002 573336
rect 107382 572736 107438 572792
rect 108578 572736 108634 572792
rect 106370 550976 106426 551032
rect 106738 550976 106794 551032
rect 106278 538056 106334 538112
rect 106922 485968 106978 486024
rect 106186 478896 106242 478952
rect 105542 395392 105598 395448
rect 104162 386960 104218 387016
rect 108302 571920 108358 571976
rect 108026 571376 108082 571432
rect 107474 560496 107530 560552
rect 108026 559000 108082 559056
rect 108026 558456 108082 558512
rect 107750 557776 107806 557832
rect 107658 542816 107714 542872
rect 107566 467880 107622 467936
rect 108946 569200 109002 569256
rect 108946 567840 109002 567896
rect 108854 567296 108910 567352
rect 108946 566500 109002 566536
rect 108946 566480 108948 566500
rect 108948 566480 109000 566500
rect 109000 566480 109002 566500
rect 108946 565836 108948 565856
rect 108948 565836 109000 565856
rect 109000 565836 109002 565856
rect 108946 565800 109002 565836
rect 108854 565256 108910 565312
rect 108946 563760 109002 563816
rect 108946 563080 109002 563136
rect 108854 562400 108910 562456
rect 108946 561060 109002 561096
rect 108946 561040 108948 561060
rect 108948 561040 109000 561060
rect 109000 561040 109002 561060
rect 108946 560496 109002 560552
rect 108946 559680 109002 559736
rect 108946 558320 109002 558376
rect 108946 557132 108948 557152
rect 108948 557132 109000 557152
rect 109000 557132 109002 557152
rect 108946 557096 109002 557132
rect 108302 556688 108358 556744
rect 108854 555600 108910 555656
rect 108946 554376 109002 554432
rect 108946 553696 109002 553752
rect 108302 552880 108358 552936
rect 108946 552200 109002 552256
rect 108026 539960 108082 540016
rect 108946 551520 109002 551576
rect 108854 550160 108910 550216
rect 109314 645904 109370 645960
rect 109590 640464 109646 640520
rect 109498 639784 109554 639840
rect 109406 637608 109462 637664
rect 109682 638832 109738 638888
rect 109130 549888 109186 549944
rect 108946 548936 109002 548992
rect 108946 547440 109002 547496
rect 108762 546896 108818 546952
rect 108946 546080 109002 546136
rect 108854 545400 108910 545456
rect 108946 544720 109002 544776
rect 108854 544040 108910 544096
rect 110510 665760 110566 665816
rect 111798 678680 111854 678736
rect 112350 678000 112406 678056
rect 111798 677320 111854 677376
rect 112718 676640 112774 676696
rect 113086 676232 113142 676288
rect 111982 675960 112038 676016
rect 113086 675416 113142 675472
rect 112074 674600 112130 674656
rect 111798 671744 111854 671800
rect 111798 671200 111854 671256
rect 111798 670520 111854 670576
rect 111798 669332 111800 669352
rect 111800 669332 111852 669352
rect 111852 669332 111854 669352
rect 111798 669296 111854 669332
rect 111982 667120 112038 667176
rect 111798 666596 111854 666632
rect 111798 666576 111800 666596
rect 111800 666576 111852 666596
rect 111852 666576 111854 666596
rect 111798 665236 111854 665272
rect 111798 665216 111800 665236
rect 111800 665216 111852 665236
rect 111852 665216 111854 665236
rect 111798 663856 111854 663912
rect 111798 662496 111854 662552
rect 111154 661136 111210 661192
rect 110602 658436 110658 658472
rect 110602 658416 110604 658436
rect 110604 658416 110656 658436
rect 110656 658416 110658 658436
rect 110602 654200 110658 654256
rect 111798 658960 111854 659016
rect 108946 543496 109002 543552
rect 108854 542000 108910 542056
rect 108946 540776 109002 540832
rect 108394 469240 108450 469296
rect 109130 491272 109186 491328
rect 109682 489912 109738 489968
rect 109038 481480 109094 481536
rect 108854 452512 108910 452568
rect 108946 395256 109002 395312
rect 109682 387912 109738 387968
rect 110510 491136 110566 491192
rect 111890 654880 111946 654936
rect 112718 669840 112774 669896
rect 112350 664400 112406 664456
rect 112350 660320 112406 660376
rect 112534 659796 112590 659832
rect 112534 659776 112536 659796
rect 112536 659776 112588 659796
rect 112588 659776 112590 659796
rect 112534 656940 112590 656976
rect 112534 656920 112536 656940
rect 112536 656920 112588 656940
rect 112588 656920 112590 656940
rect 112350 656240 112406 656296
rect 112534 655596 112536 655616
rect 112536 655596 112588 655616
rect 112588 655596 112590 655616
rect 112534 655560 112590 655596
rect 112074 650800 112130 650856
rect 111982 650120 112038 650176
rect 111982 648080 112038 648136
rect 113086 652840 113142 652896
rect 112534 651480 112590 651536
rect 113086 649440 113142 649496
rect 112994 648760 113050 648816
rect 113086 647400 113142 647456
rect 112994 645360 113050 645416
rect 113086 644680 113142 644736
rect 112810 643456 112866 643512
rect 113086 642640 113142 642696
rect 112626 642116 112682 642152
rect 112626 642096 112628 642116
rect 112628 642096 112680 642116
rect 112680 642096 112682 642116
rect 112902 639920 112958 639976
rect 113178 638560 113234 638616
rect 115294 644408 115350 644464
rect 115202 638560 115258 638616
rect 113454 568520 113510 568576
rect 114466 493312 114522 493368
rect 114466 485016 114522 485072
rect 113178 442448 113234 442504
rect 112626 392536 112682 392592
rect 113914 390768 113970 390824
rect 115202 545128 115258 545184
rect 116122 587288 116178 587344
rect 116214 583888 116270 583944
rect 116398 578176 116454 578232
rect 116306 576172 116308 576192
rect 116308 576172 116360 576192
rect 116360 576172 116362 576192
rect 116306 576136 116362 576172
rect 117134 576136 117190 576192
rect 115846 406272 115902 406328
rect 117594 587424 117650 587480
rect 117226 488416 117282 488472
rect 117226 485696 117282 485752
rect 117410 485016 117466 485072
rect 116398 380840 116454 380896
rect 115938 378528 115994 378584
rect 115478 377440 115534 377496
rect 115294 374584 115350 374640
rect 115478 373088 115534 373144
rect 115294 371864 115350 371920
rect 115294 366968 115350 367024
rect 69662 349832 69718 349888
rect 67638 290808 67694 290864
rect 67638 290128 67694 290184
rect 67638 288768 67694 288824
rect 68650 288088 68706 288144
rect 67638 287408 67694 287464
rect 67822 287000 67878 287056
rect 67730 286728 67786 286784
rect 67638 286048 67694 286104
rect 67638 285368 67694 285424
rect 67638 284416 67694 284472
rect 67638 282104 67694 282160
rect 67638 280336 67694 280392
rect 67730 279792 67786 279848
rect 67638 279248 67694 279304
rect 67638 277616 67694 277672
rect 67822 276936 67878 276992
rect 67638 275848 67694 275904
rect 67638 274896 67694 274952
rect 67730 274488 67786 274544
rect 67638 273536 67694 273592
rect 67638 270952 67694 271008
rect 67730 270816 67786 270872
rect 69018 298288 69074 298344
rect 68834 278568 68890 278624
rect 68742 276528 68798 276584
rect 68742 272176 68798 272232
rect 68190 270136 68246 270192
rect 67730 269728 67786 269784
rect 68558 268776 68614 268832
rect 67638 268368 67694 268424
rect 67638 267028 67694 267064
rect 67638 267008 67640 267028
rect 67640 267008 67692 267028
rect 67692 267008 67694 267028
rect 67730 266872 67786 266928
rect 67638 265376 67694 265432
rect 67730 264968 67786 265024
rect 67730 264152 67786 264208
rect 67638 263644 67640 263664
rect 67640 263644 67692 263664
rect 67692 263644 67694 263664
rect 67638 263608 67694 263644
rect 67638 263508 67640 263528
rect 67640 263508 67692 263528
rect 67692 263508 67694 263528
rect 67638 263472 67694 263508
rect 67638 262268 67694 262304
rect 67638 262248 67640 262268
rect 67640 262248 67692 262268
rect 67692 262248 67694 262268
rect 67730 262148 67732 262168
rect 67732 262148 67784 262168
rect 67784 262148 67786 262168
rect 67730 262112 67786 262148
rect 67638 260788 67640 260808
rect 67640 260788 67692 260808
rect 67692 260788 67694 260808
rect 67638 260752 67694 260788
rect 67730 258576 67786 258632
rect 67638 257896 67694 257952
rect 68006 256808 68062 256864
rect 67638 255332 67694 255368
rect 67638 255312 67640 255332
rect 67640 255312 67692 255332
rect 67692 255312 67694 255332
rect 67730 255212 67732 255232
rect 67732 255212 67784 255232
rect 67784 255212 67786 255232
rect 67730 255176 67786 255212
rect 67638 254768 67694 254824
rect 67638 253852 67640 253872
rect 67640 253852 67692 253872
rect 67692 253852 67694 253872
rect 67638 253816 67694 253852
rect 67638 251776 67694 251832
rect 68558 251368 68614 251424
rect 67730 251132 67732 251152
rect 67732 251132 67784 251152
rect 67784 251132 67786 251152
rect 67730 251096 67786 251132
rect 68466 249872 68522 249928
rect 67638 249056 67694 249112
rect 67730 247696 67786 247752
rect 67638 247152 67694 247208
rect 67730 246336 67786 246392
rect 67638 245792 67694 245848
rect 67638 245248 67694 245304
rect 67638 243752 67694 243808
rect 67730 243616 67786 243672
rect 68650 240896 68706 240952
rect 68742 236544 68798 236600
rect 68834 226888 68890 226944
rect 71686 292340 71688 292360
rect 71688 292340 71740 292360
rect 71740 292340 71742 292360
rect 71686 292304 71742 292340
rect 73250 294480 73306 294536
rect 75182 339904 75238 339960
rect 74630 333240 74686 333296
rect 77390 335996 77392 336016
rect 77392 335996 77444 336016
rect 77444 335996 77446 336016
rect 77390 335960 77446 335996
rect 76654 315288 76710 315344
rect 79690 339360 79746 339416
rect 81622 294616 81678 294672
rect 80702 294480 80758 294536
rect 80978 292576 81034 292632
rect 84842 339360 84898 339416
rect 88982 305632 89038 305688
rect 88706 294752 88762 294808
rect 91282 298696 91338 298752
rect 91282 298152 91338 298208
rect 95790 333920 95846 333976
rect 95790 332560 95846 332616
rect 96526 332560 96582 332616
rect 96526 295976 96582 296032
rect 97814 302776 97870 302832
rect 98734 311072 98790 311128
rect 97906 293120 97962 293176
rect 102046 335280 102102 335336
rect 103610 335144 103666 335200
rect 102046 297336 102102 297392
rect 104806 335144 104862 335200
rect 104162 294480 104218 294536
rect 107658 327664 107714 327720
rect 110234 336776 110290 336832
rect 111246 339632 111302 339688
rect 111798 337320 111854 337376
rect 115938 364248 115994 364304
rect 115846 353232 115902 353288
rect 115662 339768 115718 339824
rect 115754 338000 115810 338056
rect 118698 579672 118754 579728
rect 118882 587152 118938 587208
rect 117594 497392 117650 497448
rect 118790 545128 118846 545184
rect 117594 396616 117650 396672
rect 117502 384920 117558 384976
rect 117410 379480 117466 379536
rect 116674 369960 116730 370016
rect 117318 365200 117374 365256
rect 120262 585248 120318 585304
rect 118790 459584 118846 459640
rect 118790 453192 118846 453248
rect 121734 581576 121790 581632
rect 118514 384920 118570 384976
rect 118606 384240 118662 384296
rect 118606 383560 118662 383616
rect 118606 382220 118662 382256
rect 118606 382200 118608 382220
rect 118608 382200 118660 382220
rect 118660 382200 118662 382220
rect 118606 381556 118608 381576
rect 118608 381556 118660 381576
rect 118660 381556 118662 381576
rect 118606 381520 118662 381556
rect 118330 379480 118386 379536
rect 118606 378800 118662 378856
rect 118054 378156 118056 378176
rect 118056 378156 118108 378176
rect 118108 378156 118110 378176
rect 118054 378120 118110 378156
rect 118238 376760 118294 376816
rect 118606 376080 118662 376136
rect 118146 375400 118202 375456
rect 121458 498228 121514 498264
rect 121458 498208 121460 498228
rect 121460 498208 121512 498228
rect 121512 498208 121514 498228
rect 122930 572736 122986 572792
rect 118606 373360 118662 373416
rect 117870 372716 117872 372736
rect 117872 372716 117924 372736
rect 117924 372716 117926 372736
rect 117870 372680 117926 372716
rect 117778 371320 117834 371376
rect 118606 370640 118662 370696
rect 118606 369960 118662 370016
rect 118422 368600 118478 368656
rect 118606 367920 118662 367976
rect 117778 367240 117834 367296
rect 118146 365880 118202 365936
rect 118054 364520 118110 364576
rect 118146 363160 118202 363216
rect 117962 362480 118018 362536
rect 117686 361800 117742 361856
rect 118606 361120 118662 361176
rect 117962 360168 118018 360224
rect 117594 357040 117650 357096
rect 117778 353640 117834 353696
rect 117410 351600 117466 351656
rect 117502 347656 117558 347712
rect 117318 342080 117374 342136
rect 117410 340756 117412 340776
rect 117412 340756 117464 340776
rect 117464 340756 117466 340776
rect 117410 340720 117466 340756
rect 117318 340040 117374 340096
rect 117778 342760 117834 342816
rect 117226 337864 117282 337920
rect 117226 336776 117282 336832
rect 116674 318008 116730 318064
rect 116582 292032 116638 292088
rect 118606 359760 118662 359816
rect 118146 359080 118202 359136
rect 118606 358400 118662 358456
rect 118606 357040 118662 357096
rect 118606 356360 118662 356416
rect 118514 355680 118570 355736
rect 118606 354356 118608 354376
rect 118608 354356 118660 354376
rect 118660 354356 118662 354376
rect 118606 354320 118662 354356
rect 118606 350920 118662 350976
rect 118606 350240 118662 350296
rect 118606 348880 118662 348936
rect 118514 348200 118570 348256
rect 118606 347520 118662 347576
rect 118514 346160 118570 346216
rect 118606 345480 118662 345536
rect 118606 344800 118662 344856
rect 118606 343440 118662 343496
rect 118514 342080 118570 342136
rect 117134 293256 117190 293312
rect 118974 295160 119030 295216
rect 119342 294752 119398 294808
rect 119710 361528 119766 361584
rect 119710 337864 119766 337920
rect 119526 294616 119582 294672
rect 69202 281288 69258 281344
rect 69110 260208 69166 260264
rect 69202 255856 69258 255912
rect 69110 244296 69166 244352
rect 121550 456068 121606 456104
rect 121550 456048 121552 456068
rect 121552 456048 121604 456068
rect 121604 456048 121606 456068
rect 122838 494672 122894 494728
rect 121550 439320 121606 439376
rect 121734 439320 121790 439376
rect 121550 387812 121552 387832
rect 121552 387812 121604 387832
rect 121604 387812 121606 387832
rect 121550 387776 121606 387812
rect 121458 291760 121514 291816
rect 121550 291080 121606 291136
rect 121458 290400 121514 290456
rect 120814 289720 120870 289776
rect 121550 289040 121606 289096
rect 121458 288380 121514 288416
rect 121458 288360 121460 288380
rect 121460 288360 121512 288380
rect 121512 288360 121514 288380
rect 121550 287680 121606 287736
rect 120722 287000 120778 287056
rect 121550 285640 121606 285696
rect 121458 284960 121514 285016
rect 121550 284280 121606 284336
rect 121458 283600 121514 283656
rect 121458 282940 121514 282976
rect 121458 282920 121460 282940
rect 121460 282920 121512 282940
rect 121512 282920 121514 282940
rect 121458 281580 121514 281616
rect 121458 281560 121460 281580
rect 121460 281560 121512 281580
rect 121512 281560 121514 281580
rect 121550 280880 121606 280936
rect 121458 280220 121514 280256
rect 121458 280200 121460 280220
rect 121460 280200 121512 280220
rect 121512 280200 121514 280220
rect 121550 279520 121606 279576
rect 121458 278840 121514 278896
rect 121550 278160 121606 278216
rect 120814 277480 120870 277536
rect 120722 269320 120778 269376
rect 120170 250960 120226 251016
rect 120630 250960 120686 251016
rect 120078 249600 120134 249656
rect 69846 241576 69902 241632
rect 71778 233144 71834 233200
rect 75826 234368 75882 234424
rect 86130 237088 86186 237144
rect 91742 231784 91798 231840
rect 69018 186904 69074 186960
rect 102046 177656 102102 177712
rect 105726 177656 105782 177712
rect 107566 177656 107622 177712
rect 118606 190984 118662 191040
rect 121458 276800 121514 276856
rect 121458 276120 121514 276176
rect 121550 275440 121606 275496
rect 121458 274780 121514 274816
rect 121458 274760 121460 274780
rect 121460 274760 121512 274780
rect 121512 274760 121514 274780
rect 122746 286320 122802 286376
rect 124310 495508 124366 495544
rect 124310 495488 124312 495508
rect 124312 495488 124364 495508
rect 124364 495488 124366 495508
rect 124126 378700 124128 378720
rect 124128 378700 124180 378720
rect 124180 378700 124182 378720
rect 124126 378664 124182 378700
rect 124402 392536 124458 392592
rect 123574 295160 123630 295216
rect 122194 282240 122250 282296
rect 121550 274080 121606 274136
rect 121458 273400 121514 273456
rect 121458 272720 121514 272776
rect 121458 271360 121514 271416
rect 121550 270000 121606 270056
rect 121458 268640 121514 268696
rect 121458 267960 121514 268016
rect 121550 267280 121606 267336
rect 121458 266600 121514 266656
rect 121550 265920 121606 265976
rect 121458 265240 121514 265296
rect 121550 263880 121606 263936
rect 121458 263200 121514 263256
rect 121458 262520 121514 262576
rect 121458 261876 121460 261896
rect 121460 261876 121512 261896
rect 121512 261876 121514 261896
rect 121458 261840 121514 261876
rect 121550 261160 121606 261216
rect 121458 260480 121514 260536
rect 121458 259800 121514 259856
rect 121642 259120 121698 259176
rect 121550 258440 121606 258496
rect 121550 257760 121606 257816
rect 121458 257080 121514 257136
rect 121458 256400 121514 256456
rect 121550 255720 121606 255776
rect 121458 255040 121514 255096
rect 122102 254360 122158 254416
rect 121458 253680 121514 253736
rect 121550 253000 121606 253056
rect 121458 252320 121514 252376
rect 121458 251640 121514 251696
rect 121458 250280 121514 250336
rect 121550 248920 121606 248976
rect 121458 248240 121514 248296
rect 121550 247560 121606 247616
rect 121550 246880 121606 246936
rect 121458 246200 121514 246256
rect 121458 245520 121514 245576
rect 121550 244840 121606 244896
rect 121458 244160 121514 244216
rect 121458 242820 121514 242856
rect 121458 242800 121460 242820
rect 121460 242800 121512 242820
rect 121512 242800 121514 242820
rect 121550 242120 121606 242176
rect 121458 240760 121514 240816
rect 121458 240080 121514 240136
rect 122286 272040 122342 272096
rect 120722 199280 120778 199336
rect 110694 177656 110750 177712
rect 109958 176976 110014 177032
rect 124310 314628 124366 314664
rect 124310 314608 124312 314628
rect 124312 314608 124364 314628
rect 124364 314608 124366 314628
rect 125966 535472 126022 535528
rect 127070 583752 127126 583808
rect 127254 589872 127310 589928
rect 125598 293256 125654 293312
rect 126242 293120 126298 293176
rect 130106 585384 130162 585440
rect 127622 297336 127678 297392
rect 128726 342216 128782 342272
rect 131210 585112 131266 585168
rect 129922 378664 129978 378720
rect 129738 337320 129794 337376
rect 129922 318008 129978 318064
rect 129922 317364 129924 317384
rect 129924 317364 129976 317384
rect 129976 317364 129978 317384
rect 129922 317328 129978 317364
rect 130290 316104 130346 316160
rect 130474 292032 130530 292088
rect 132866 442312 132922 442368
rect 131762 342216 131818 342272
rect 132590 347656 132646 347712
rect 132498 320184 132554 320240
rect 133878 353368 133934 353424
rect 130474 215872 130530 215928
rect 134522 359216 134578 359272
rect 134154 338000 134210 338056
rect 135166 338000 135222 338056
rect 135166 337320 135222 337376
rect 133786 242120 133842 242176
rect 136914 570696 136970 570752
rect 136822 491136 136878 491192
rect 138110 564984 138166 565040
rect 139490 570560 139546 570616
rect 140962 482976 141018 483032
rect 139306 363568 139362 363624
rect 135994 192616 136050 192672
rect 138018 300092 138020 300112
rect 138020 300092 138072 300112
rect 138072 300092 138074 300112
rect 138018 300056 138074 300092
rect 116950 177656 117006 177712
rect 119710 177656 119766 177712
rect 121182 177656 121238 177712
rect 123298 177656 123354 177712
rect 142250 485016 142306 485072
rect 141054 371320 141110 371376
rect 140870 345616 140926 345672
rect 397458 702616 397514 702672
rect 143538 371320 143594 371376
rect 141422 295976 141478 296032
rect 140870 238584 140926 238640
rect 140870 237360 140926 237416
rect 141514 237360 141570 237416
rect 143446 348472 143502 348528
rect 143722 253136 143778 253192
rect 145194 351056 145250 351112
rect 146206 348336 146262 348392
rect 144918 238584 144974 238640
rect 146482 359352 146538 359408
rect 147218 240760 147274 240816
rect 150530 346296 150586 346352
rect 150530 345616 150586 345672
rect 148414 189624 148470 189680
rect 155222 400288 155278 400344
rect 151818 279384 151874 279440
rect 153198 284824 153254 284880
rect 152554 239808 152610 239864
rect 152646 226208 152702 226264
rect 153842 184184 153898 184240
rect 128266 177656 128322 177712
rect 129462 177656 129518 177712
rect 130934 177656 130990 177712
rect 132406 177656 132462 177712
rect 115846 177112 115902 177168
rect 126058 177112 126114 177168
rect 134706 177112 134762 177168
rect 97814 176704 97870 176760
rect 100666 176704 100722 176760
rect 108118 176704 108174 176760
rect 112258 176704 112314 176760
rect 114374 176704 114430 176760
rect 124494 176704 124550 176760
rect 128174 176704 128230 176760
rect 133142 176724 133198 176760
rect 133142 176704 133144 176724
rect 133144 176704 133196 176724
rect 133196 176704 133198 176724
rect 159454 177384 159510 177440
rect 136086 176740 136088 176760
rect 136088 176740 136140 176760
rect 136140 176740 136142 176760
rect 136086 176704 136142 176740
rect 148230 176704 148286 176760
rect 158902 176704 158958 176760
rect 162306 298152 162362 298208
rect 162306 231648 162362 231704
rect 163594 234368 163650 234424
rect 169022 390768 169078 390824
rect 166446 250416 166502 250472
rect 166354 230424 166410 230480
rect 164882 181600 164938 181656
rect 160834 175888 160890 175944
rect 98366 175344 98422 175400
rect 102046 175344 102102 175400
rect 118422 175344 118478 175400
rect 121918 175344 121974 175400
rect 167642 204856 167698 204912
rect 177302 387912 177358 387968
rect 170402 335960 170458 336016
rect 169022 222808 169078 222864
rect 167734 176976 167790 177032
rect 167642 171536 167698 171592
rect 173254 359352 173310 359408
rect 169114 179968 169170 180024
rect 172426 320204 172482 320240
rect 172426 320184 172428 320204
rect 172428 320184 172480 320204
rect 172480 320184 172482 320204
rect 170586 177248 170642 177304
rect 174542 337320 174598 337376
rect 173162 221448 173218 221504
rect 67638 126248 67694 126304
rect 67638 91024 67694 91080
rect 164882 95104 164938 95160
rect 85578 94696 85634 94752
rect 112350 94696 112406 94752
rect 125414 94696 125470 94752
rect 118238 93608 118294 93664
rect 98550 93472 98606 93528
rect 129462 93472 129518 93528
rect 103334 93200 103390 93256
rect 110142 93200 110198 93256
rect 85118 92384 85174 92440
rect 86774 92384 86830 92440
rect 88982 92384 89038 92440
rect 75366 91160 75422 91216
rect 90546 91704 90602 91760
rect 95054 91704 95110 91760
rect 88062 91160 88118 91216
rect 92386 91160 92442 91216
rect 93766 91160 93822 91216
rect 101862 91432 101918 91488
rect 97906 91296 97962 91352
rect 99194 91296 99250 91352
rect 95146 91160 95202 91216
rect 96526 91160 96582 91216
rect 97814 91160 97870 91216
rect 99286 91160 99342 91216
rect 100206 91160 100262 91216
rect 100574 91160 100630 91216
rect 102046 91296 102102 91352
rect 101954 91160 102010 91216
rect 107750 92384 107806 92440
rect 114374 92384 114430 92440
rect 115478 92384 115534 92440
rect 120354 92404 120410 92440
rect 120354 92384 120356 92404
rect 120356 92384 120408 92404
rect 120408 92384 120410 92404
rect 107290 91296 107346 91352
rect 103426 91160 103482 91216
rect 104438 91160 104494 91216
rect 104806 91160 104862 91216
rect 105542 91160 105598 91216
rect 106094 91160 106150 91216
rect 107566 91160 107622 91216
rect 110234 91296 110290 91352
rect 108946 91160 109002 91216
rect 104806 81368 104862 81424
rect 110326 91160 110382 91216
rect 111246 91160 111302 91216
rect 112442 91160 112498 91216
rect 99286 78512 99342 78568
rect 122102 92384 122158 92440
rect 117134 91296 117190 91352
rect 119894 91296 119950 91352
rect 114466 91160 114522 91216
rect 114926 91160 114982 91216
rect 115846 91160 115902 91216
rect 112442 85448 112498 85504
rect 117226 91160 117282 91216
rect 119986 91160 120042 91216
rect 120630 91160 120686 91216
rect 133142 93472 133198 93528
rect 151726 93472 151782 93528
rect 130750 92384 130806 92440
rect 135166 92384 135222 92440
rect 136086 92384 136142 92440
rect 151634 92384 151690 92440
rect 126518 91704 126574 91760
rect 122838 91432 122894 91488
rect 122746 91160 122802 91216
rect 123298 91160 123354 91216
rect 123942 91160 123998 91216
rect 124770 91160 124826 91216
rect 126886 91160 126942 91216
rect 127622 91160 127678 91216
rect 132406 91160 132462 91216
rect 151450 91160 151506 91216
rect 153014 91432 153070 91488
rect 79322 51720 79378 51776
rect 81438 26832 81494 26888
rect 106278 25472 106334 25528
rect 167918 111732 167920 111752
rect 167920 111732 167972 111752
rect 167972 111732 167974 111752
rect 167918 111696 167974 111732
rect 167734 110064 167790 110120
rect 167642 93880 167698 93936
rect 168102 108704 168158 108760
rect 175186 181328 175242 181384
rect 176198 233008 176254 233064
rect 182914 181600 182970 181656
rect 184386 238448 184442 238504
rect 187054 177384 187110 177440
rect 187054 82184 187110 82240
rect 188526 331200 188582 331256
rect 188434 184184 188490 184240
rect 188526 82048 188582 82104
rect 171966 3440 172022 3496
rect 209042 379480 209098 379536
rect 192574 93744 192630 93800
rect 195242 360304 195298 360360
rect 206466 365744 206522 365800
rect 198186 360168 198242 360224
rect 198094 358264 198150 358320
rect 198002 353640 198058 353696
rect 197358 349560 197414 349616
rect 197358 347384 197414 347440
rect 198002 342624 198058 342680
rect 197358 340584 197414 340640
rect 197358 337864 197414 337920
rect 197358 335824 197414 335880
rect 197358 331744 197414 331800
rect 197358 329024 197414 329080
rect 197358 327140 197414 327176
rect 197358 327120 197360 327140
rect 197360 327120 197412 327140
rect 197412 327120 197414 327140
rect 197358 322360 197414 322416
rect 197358 320204 197414 320240
rect 197358 320184 197360 320204
rect 197360 320184 197412 320204
rect 197412 320184 197414 320204
rect 196806 309304 196862 309360
rect 197358 315424 197414 315480
rect 197358 313384 197414 313440
rect 197358 311344 197414 311400
rect 197266 306584 197322 306640
rect 197358 304544 197414 304600
rect 197358 302504 197414 302560
rect 198278 356360 198334 356416
rect 198278 351464 198334 351520
rect 198186 344664 198242 344720
rect 198094 324944 198150 325000
rect 199014 333784 199070 333840
rect 198646 318144 198702 318200
rect 197450 301280 197506 301336
rect 198002 301280 198058 301336
rect 197450 300872 197506 300928
rect 197358 299920 197414 299976
rect 197358 297744 197414 297800
rect 197450 295704 197506 295760
rect 197450 293664 197506 293720
rect 197450 290944 197506 291000
rect 197450 288904 197506 288960
rect 197450 286864 197506 286920
rect 197450 284144 197506 284200
rect 197450 282104 197506 282160
rect 197450 280200 197506 280256
rect 197450 277500 197506 277536
rect 197450 277480 197452 277500
rect 197452 277480 197504 277500
rect 197504 277480 197506 277500
rect 197358 275304 197414 275360
rect 197358 273284 197414 273320
rect 197358 273264 197360 273284
rect 197360 273264 197412 273284
rect 197412 273264 197414 273284
rect 197358 271224 197414 271280
rect 197358 268504 197414 268560
rect 197358 266464 197414 266520
rect 197358 264424 197414 264480
rect 197358 261704 197414 261760
rect 197358 259664 197414 259720
rect 197358 257624 197414 257680
rect 197358 255584 197414 255640
rect 197358 252864 197414 252920
rect 197358 248804 197414 248840
rect 197358 248784 197360 248804
rect 197360 248784 197412 248804
rect 197412 248784 197414 248804
rect 197358 246200 197414 246256
rect 197174 239400 197230 239456
rect 198646 271224 198702 271280
rect 198462 242120 198518 242176
rect 198094 177384 198150 177440
rect 217966 362344 218022 362400
rect 223486 362208 223542 362264
rect 227718 363024 227774 363080
rect 231858 394712 231914 394768
rect 253202 389272 253258 389328
rect 247038 364384 247094 364440
rect 248970 361664 249026 361720
rect 249706 361684 249762 361720
rect 249706 361664 249708 361684
rect 249708 361664 249760 361684
rect 249760 361664 249762 361684
rect 261850 364520 261906 364576
rect 274730 361936 274786 361992
rect 274730 361528 274786 361584
rect 285034 363160 285090 363216
rect 291474 360168 291530 360224
rect 293222 360440 293278 360496
rect 300122 361800 300178 361856
rect 304354 360168 304410 360224
rect 271970 359488 272026 359544
rect 317050 359488 317106 359544
rect 199658 358808 199714 358864
rect 319350 358808 319406 358864
rect 319350 356360 319406 356416
rect 319902 361800 319958 361856
rect 198922 313384 198978 313440
rect 201406 239808 201462 239864
rect 198278 91568 198334 91624
rect 204902 239400 204958 239456
rect 207662 237904 207718 237960
rect 206282 181464 206338 181520
rect 206466 181464 206522 181520
rect 211618 235184 211674 235240
rect 209134 191120 209190 191176
rect 209042 184184 209098 184240
rect 207662 93744 207718 93800
rect 215942 227024 215998 227080
rect 214562 178608 214618 178664
rect 213918 176160 213974 176216
rect 213918 175072 213974 175128
rect 214010 174664 214066 174720
rect 213918 173712 213974 173768
rect 214010 173304 214066 173360
rect 213918 172352 213974 172408
rect 214102 171944 214158 172000
rect 213918 171012 213974 171048
rect 213918 170992 213920 171012
rect 213920 170992 213972 171012
rect 213972 170992 213974 171012
rect 214010 170720 214066 170776
rect 214654 169360 214710 169416
rect 213918 168292 213974 168328
rect 213918 168272 213920 168292
rect 213920 168272 213972 168292
rect 213972 168272 213974 168292
rect 214010 168000 214066 168056
rect 213918 166912 213974 166968
rect 214102 166640 214158 166696
rect 214010 166096 214066 166152
rect 213918 165280 213974 165336
rect 214010 164736 214066 164792
rect 213918 163376 213974 163432
rect 213918 162732 213920 162752
rect 213920 162732 213972 162752
rect 213972 162732 213974 162752
rect 213918 162696 213974 162732
rect 214010 162016 214066 162072
rect 213918 161372 213920 161392
rect 213920 161372 213972 161392
rect 213972 161372 213974 161392
rect 213918 161336 213974 161372
rect 214010 160792 214066 160848
rect 213918 159840 213974 159896
rect 214010 159432 214066 159488
rect 213918 157392 213974 157448
rect 213918 157292 213920 157312
rect 213920 157292 213972 157312
rect 213972 157292 213974 157312
rect 213918 157256 213974 157292
rect 214010 156848 214066 156904
rect 213918 155916 213974 155952
rect 213918 155896 213920 155916
rect 213920 155896 213972 155916
rect 213972 155896 213974 155916
rect 214010 155352 214066 155408
rect 213918 153856 213974 153912
rect 213366 153176 213422 153232
rect 214010 152632 214066 152688
rect 213918 151952 213974 152008
rect 214010 150864 214066 150920
rect 213918 150592 213974 150648
rect 214010 150048 214066 150104
rect 213918 149504 213974 149560
rect 214930 169632 214986 169688
rect 215022 151816 215078 151872
rect 214746 148824 214802 148880
rect 214562 148008 214618 148064
rect 214010 146648 214066 146704
rect 213918 146396 213974 146432
rect 213918 146376 213920 146396
rect 213920 146376 213972 146396
rect 213972 146376 213974 146396
rect 213918 145288 213974 145344
rect 214010 143928 214066 143984
rect 213918 143520 213974 143576
rect 214010 142704 214066 142760
rect 213918 142296 213974 142352
rect 214010 141344 214066 141400
rect 213918 140820 213974 140856
rect 213918 140800 213920 140820
rect 213920 140800 213972 140820
rect 213972 140800 213974 140820
rect 213918 139984 213974 140040
rect 213918 138760 213974 138816
rect 214010 137400 214066 137456
rect 213918 136740 213974 136776
rect 213918 136720 213920 136740
rect 213920 136720 213972 136740
rect 213972 136720 213974 136740
rect 213918 136040 213974 136096
rect 214010 134272 214066 134328
rect 213918 134000 213974 134056
rect 213918 132932 213974 132968
rect 213918 132912 213920 132932
rect 213920 132912 213972 132932
rect 213972 132912 213974 132932
rect 213918 132776 213974 132832
rect 213918 131416 213974 131472
rect 214010 130056 214066 130112
rect 213918 129820 213920 129840
rect 213920 129820 213972 129840
rect 213972 129820 213974 129840
rect 213918 129784 213974 129820
rect 213918 128832 213974 128888
rect 214010 127472 214066 127528
rect 213918 127064 213974 127120
rect 214010 126112 214066 126168
rect 213918 125704 213974 125760
rect 214010 124752 214066 124808
rect 213918 124344 213974 124400
rect 214010 123528 214066 123584
rect 213918 123120 213974 123176
rect 214010 122168 214066 122224
rect 213918 121508 213974 121544
rect 213918 121488 213920 121508
rect 213920 121488 213972 121508
rect 213972 121488 213974 121508
rect 214010 120808 214066 120864
rect 213918 120148 213974 120184
rect 213918 120128 213920 120148
rect 213920 120128 213972 120148
rect 213972 120128 213974 120148
rect 214010 119584 214066 119640
rect 213458 119040 213514 119096
rect 213918 118904 213974 118960
rect 214010 117544 214066 117600
rect 213918 117272 213974 117328
rect 214010 116184 214066 116240
rect 213918 115912 213974 115968
rect 213918 114960 213974 115016
rect 214010 113600 214066 113656
rect 213918 113212 213974 113248
rect 213918 113192 213920 113212
rect 213920 113192 213972 113212
rect 213972 113192 213974 113212
rect 214010 112240 214066 112296
rect 213918 111868 213920 111888
rect 213920 111868 213972 111888
rect 213972 111868 213974 111888
rect 213918 111832 213974 111868
rect 214010 110880 214066 110936
rect 213918 110508 213920 110528
rect 213920 110508 213972 110528
rect 213972 110508 213974 110528
rect 213918 110472 213974 110508
rect 214010 109656 214066 109712
rect 213918 109132 213974 109168
rect 213918 109112 213920 109132
rect 213920 109112 213972 109132
rect 213972 109112 213974 109132
rect 214010 108296 214066 108352
rect 213918 107888 213974 107944
rect 214010 106936 214066 106992
rect 213918 106528 213974 106584
rect 214010 105712 214066 105768
rect 213918 105032 213974 105088
rect 213918 103672 213974 103728
rect 213918 102448 213974 102504
rect 214010 101224 214066 101280
rect 213918 101088 213974 101144
rect 214010 99728 214066 99784
rect 213918 99456 213974 99512
rect 214010 98368 214066 98424
rect 213918 97996 213920 98016
rect 213920 97996 213972 98016
rect 213972 97996 213974 98016
rect 213918 97960 213974 97996
rect 214746 144880 214802 144936
rect 214654 139576 214710 139632
rect 214654 138080 214710 138136
rect 214838 102312 214894 102368
rect 214654 100000 214710 100056
rect 214654 97008 214710 97064
rect 214746 95784 214802 95840
rect 227074 235864 227130 235920
rect 232502 180104 232558 180160
rect 224222 175888 224278 175944
rect 244462 238448 244518 238504
rect 240966 185544 241022 185600
rect 240874 178744 240930 178800
rect 243542 178880 243598 178936
rect 245106 176024 245162 176080
rect 248050 175788 248052 175808
rect 248052 175788 248104 175808
rect 248104 175788 248106 175808
rect 248050 175752 248106 175788
rect 252834 238756 252836 238776
rect 252836 238756 252888 238776
rect 252888 238756 252890 238776
rect 252834 238720 252890 238756
rect 249154 175208 249210 175264
rect 249246 172760 249302 172816
rect 249338 171400 249394 171456
rect 249154 161472 249210 161528
rect 250258 169496 250314 169552
rect 251914 228248 251970 228304
rect 252006 225528 252062 225584
rect 252006 188264 252062 188320
rect 252466 174664 252522 174720
rect 252466 173712 252522 173768
rect 252466 172352 252522 172408
rect 252374 171808 252430 171864
rect 252466 170856 252522 170912
rect 252374 170448 252430 170504
rect 252466 170040 252522 170096
rect 252466 168136 252522 168192
rect 251454 160112 251510 160168
rect 251362 159160 251418 159216
rect 252374 167184 252430 167240
rect 252466 166660 252522 166696
rect 252466 166640 252468 166660
rect 252468 166640 252520 166660
rect 252520 166640 252522 166660
rect 252374 166232 252430 166288
rect 252466 165688 252522 165744
rect 252466 165280 252522 165336
rect 252374 164736 252430 164792
rect 252466 163920 252522 163976
rect 252374 162968 252430 163024
rect 252466 162424 252522 162480
rect 252374 162016 252430 162072
rect 252466 160520 252522 160576
rect 252466 159568 252522 159624
rect 252374 158208 252430 158264
rect 252466 157800 252522 157856
rect 252466 157292 252468 157312
rect 252468 157292 252520 157312
rect 252520 157292 252522 157312
rect 252466 157256 252522 157292
rect 251546 156848 251602 156904
rect 251178 156304 251234 156360
rect 252374 155896 252430 155952
rect 250074 155352 250130 155408
rect 252466 154944 252522 155000
rect 252466 154400 252522 154456
rect 251454 153312 251510 153368
rect 252466 153076 252468 153096
rect 252468 153076 252520 153096
rect 252520 153076 252522 153096
rect 252466 153040 252522 153076
rect 252374 152632 252430 152688
rect 252282 152088 252338 152144
rect 252834 169088 252890 169144
rect 252742 164328 252798 164384
rect 252650 151680 252706 151736
rect 252466 151136 252522 151192
rect 251454 150728 251510 150784
rect 249890 149776 249946 149832
rect 251362 149232 251418 149288
rect 251362 146512 251418 146568
rect 249798 139440 249854 139496
rect 216678 114552 216734 114608
rect 242898 10920 242954 10976
rect 243542 10920 243598 10976
rect 240506 3984 240562 4040
rect 242990 3304 243046 3360
rect 251178 125704 251234 125760
rect 251730 118768 251786 118824
rect 252466 150184 252522 150240
rect 252466 148824 252522 148880
rect 252374 148280 252430 148336
rect 252466 147464 252522 147520
rect 252098 146920 252154 146976
rect 252466 145560 252522 145616
rect 252374 145016 252430 145072
rect 252466 144064 252522 144120
rect 252374 143656 252430 143712
rect 252466 143112 252522 143168
rect 252374 142704 252430 142760
rect 253202 140800 253258 140856
rect 252466 139848 252522 139904
rect 252466 138488 252522 138544
rect 252466 136720 252522 136776
rect 252466 136584 252522 136640
rect 252282 136176 252338 136232
rect 252374 135632 252430 135688
rect 252190 135224 252246 135280
rect 252466 134680 252522 134736
rect 252374 134272 252430 134328
rect 252466 133728 252522 133784
rect 252282 133320 252338 133376
rect 252374 132776 252430 132832
rect 252466 132388 252522 132424
rect 252466 132368 252468 132388
rect 252468 132368 252520 132388
rect 252520 132368 252522 132388
rect 252282 131824 252338 131880
rect 252374 131416 252430 131472
rect 252466 130872 252522 130928
rect 252374 130464 252430 130520
rect 252466 130056 252522 130112
rect 252282 129104 252338 129160
rect 252466 129512 252522 129568
rect 252374 128560 252430 128616
rect 252282 128172 252338 128208
rect 252282 128152 252284 128172
rect 252284 128152 252336 128172
rect 252336 128152 252338 128172
rect 252098 125296 252154 125352
rect 252466 127608 252522 127664
rect 252374 127200 252430 127256
rect 252466 126656 252522 126712
rect 252466 126248 252522 126304
rect 252190 123936 252246 123992
rect 252466 124752 252522 124808
rect 252374 124344 252430 124400
rect 252466 123392 252522 123448
rect 252282 122984 252338 123040
rect 252466 122440 252522 122496
rect 252374 122032 252430 122088
rect 252282 121488 252338 121544
rect 251914 121080 251970 121136
rect 252466 120536 252522 120592
rect 252466 120128 252522 120184
rect 252466 119584 252522 119640
rect 251822 117272 251878 117328
rect 251730 107888 251786 107944
rect 251730 106528 251786 106584
rect 251362 101768 251418 101824
rect 251822 100816 251878 100872
rect 252466 119176 252522 119232
rect 252466 118224 252522 118280
rect 252374 117816 252430 117872
rect 252374 116864 252430 116920
rect 252466 116320 252522 116376
rect 252282 115912 252338 115968
rect 252466 115368 252522 115424
rect 252374 114960 252430 115016
rect 252466 114008 252522 114064
rect 252374 113464 252430 113520
rect 252098 113056 252154 113112
rect 252282 111716 252338 111752
rect 252282 111696 252284 111716
rect 252284 111696 252336 111716
rect 252336 111696 252338 111716
rect 252466 112648 252522 112704
rect 252466 112104 252522 112160
rect 252374 111152 252430 111208
rect 252466 110744 252522 110800
rect 252466 110236 252468 110256
rect 252468 110236 252520 110256
rect 252520 110236 252522 110256
rect 252466 110200 252522 110236
rect 252374 109792 252430 109848
rect 252282 109248 252338 109304
rect 252466 108840 252522 108896
rect 252190 108296 252246 108352
rect 252466 107480 252522 107536
rect 252098 106936 252154 106992
rect 252466 105984 252522 106040
rect 252374 105576 252430 105632
rect 252282 105032 252338 105088
rect 252282 104080 252338 104136
rect 252466 104624 252522 104680
rect 252374 103672 252430 103728
rect 252466 103128 252522 103184
rect 252466 102720 252522 102776
rect 252374 102176 252430 102232
rect 251914 98504 251970 98560
rect 252466 101360 252522 101416
rect 252466 100408 252522 100464
rect 252374 99864 252430 99920
rect 252282 99456 252338 99512
rect 252466 98912 252522 98968
rect 252190 97960 252246 98016
rect 252466 97552 252522 97608
rect 251178 96192 251234 96248
rect 251362 82184 251418 82240
rect 249246 19896 249302 19952
rect 252466 96600 252522 96656
rect 253478 141752 253534 141808
rect 253478 140936 253534 140992
rect 257434 145560 257490 145616
rect 265622 233008 265678 233064
rect 259642 176024 259698 176080
rect 259458 60696 259514 60752
rect 261482 84768 261538 84824
rect 260194 79328 260250 79384
rect 260194 62056 260250 62112
rect 260194 60696 260250 60752
rect 271878 195200 271934 195256
rect 267738 20576 267794 20632
rect 268474 20576 268530 20632
rect 271878 61512 271934 61568
rect 273350 148280 273406 148336
rect 273166 61512 273222 61568
rect 276018 76608 276074 76664
rect 276662 29552 276718 29608
rect 279422 181464 279478 181520
rect 278042 29552 278098 29608
rect 280802 62736 280858 62792
rect 289450 233144 289506 233200
rect 293222 234504 293278 234560
rect 287702 211928 287758 211984
rect 284298 46824 284354 46880
rect 285218 61376 285274 61432
rect 285218 46824 285274 46880
rect 305642 238584 305698 238640
rect 299202 231784 299258 231840
rect 289082 75112 289138 75168
rect 307390 175208 307446 175264
rect 307298 173576 307354 173632
rect 306746 172216 306802 172272
rect 307114 171808 307170 171864
rect 307574 174800 307630 174856
rect 307482 174392 307538 174448
rect 307666 174004 307722 174040
rect 307666 173984 307668 174004
rect 307668 173984 307720 174004
rect 307720 173984 307722 174004
rect 307482 173168 307538 173224
rect 307666 172644 307722 172680
rect 307666 172624 307668 172644
rect 307668 172624 307720 172644
rect 307720 172624 307722 172644
rect 307666 171400 307722 171456
rect 306562 168816 306618 168872
rect 306562 166368 306618 166424
rect 306746 170992 306802 171048
rect 306930 170584 306986 170640
rect 306746 166776 306802 166832
rect 307666 170176 307722 170232
rect 307482 169788 307538 169824
rect 307482 169768 307484 169788
rect 307484 169768 307536 169788
rect 307536 169768 307538 169788
rect 307574 169224 307630 169280
rect 307666 168444 307668 168464
rect 307668 168444 307720 168464
rect 307720 168444 307722 168464
rect 307666 168408 307722 168444
rect 307298 168000 307354 168056
rect 307574 167592 307630 167648
rect 307482 165824 307538 165880
rect 307206 165416 307262 165472
rect 307022 165008 307078 165064
rect 306930 163784 306986 163840
rect 305642 162968 305698 163024
rect 306930 162968 306986 163024
rect 304354 149640 304410 149696
rect 303158 143928 303214 143984
rect 306562 161200 306618 161256
rect 306930 159976 306986 160032
rect 306746 158208 306802 158264
rect 306562 156984 306618 157040
rect 306562 155624 306618 155680
rect 306654 153584 306710 153640
rect 305826 150592 305882 150648
rect 305734 118768 305790 118824
rect 305642 109248 305698 109304
rect 304354 3440 304410 3496
rect 306746 150184 306802 150240
rect 306930 148416 306986 148472
rect 306746 146784 306802 146840
rect 306930 144200 306986 144256
rect 306562 142976 306618 143032
rect 306562 142024 306618 142080
rect 307114 164192 307170 164248
rect 307666 167184 307722 167240
rect 307666 164600 307722 164656
rect 307390 163376 307446 163432
rect 307666 162968 307722 163024
rect 307482 162424 307538 162480
rect 307574 162016 307630 162072
rect 307666 161608 307722 161664
rect 307574 160792 307630 160848
rect 307666 160384 307722 160440
rect 307574 159568 307630 159624
rect 307666 159024 307722 159080
rect 307390 158616 307446 158672
rect 307114 157392 307170 157448
rect 307298 154808 307354 154864
rect 307298 154400 307354 154456
rect 307482 157800 307538 157856
rect 307574 156576 307630 156632
rect 307666 156168 307722 156224
rect 307666 155216 307722 155272
rect 307574 153992 307630 154048
rect 307666 153176 307722 153232
rect 307482 152632 307538 152688
rect 307574 152224 307630 152280
rect 307114 142432 307170 142488
rect 306562 139032 306618 139088
rect 306562 136584 306618 136640
rect 306562 134816 306618 134872
rect 307022 134000 307078 134056
rect 306562 133592 306618 133648
rect 306930 133184 306986 133240
rect 306562 131008 306618 131064
rect 306930 130600 306986 130656
rect 306930 129240 306986 129296
rect 305918 123256 305974 123312
rect 305826 108296 305882 108352
rect 306562 118632 306618 118688
rect 306746 116592 306802 116648
rect 306930 112648 306986 112704
rect 306746 110200 306802 110256
rect 306746 109248 306802 109304
rect 306930 109248 306986 109304
rect 306930 105848 306986 105904
rect 306930 104624 306986 104680
rect 306562 101224 306618 101280
rect 306930 100816 306986 100872
rect 306562 100408 306618 100464
rect 306930 98640 306986 98696
rect 307666 151816 307722 151872
rect 307574 151408 307630 151464
rect 307666 151000 307722 151056
rect 307666 149776 307722 149832
rect 307574 149232 307630 149288
rect 307574 148824 307630 148880
rect 307666 148008 307722 148064
rect 307390 147600 307446 147656
rect 307298 139576 307354 139632
rect 307298 138624 307354 138680
rect 307206 136992 307262 137048
rect 307114 114008 307170 114064
rect 307298 135224 307354 135280
rect 307574 147192 307630 147248
rect 307666 146396 307722 146432
rect 307666 146376 307668 146396
rect 307668 146376 307720 146396
rect 307720 146376 307722 146396
rect 307666 145832 307722 145888
rect 307574 145424 307630 145480
rect 307666 144608 307722 144664
rect 307574 143792 307630 143848
rect 307666 143384 307722 143440
rect 307574 141616 307630 141672
rect 307482 141208 307538 141264
rect 307666 140820 307722 140856
rect 307666 140800 307668 140820
rect 307668 140800 307720 140820
rect 307720 140800 307722 140820
rect 307298 132640 307354 132696
rect 307574 140392 307630 140448
rect 307666 139984 307722 140040
rect 307666 138216 307722 138272
rect 307666 137808 307722 137864
rect 307574 136176 307630 136232
rect 307666 135632 307722 135688
rect 307482 132232 307538 132288
rect 307574 131824 307630 131880
rect 307666 131416 307722 131472
rect 307482 129784 307538 129840
rect 307666 128832 307722 128888
rect 307574 128424 307630 128480
rect 307574 128016 307630 128072
rect 307666 127200 307722 127256
rect 307482 126792 307538 126848
rect 307574 126384 307630 126440
rect 307666 125840 307722 125896
rect 307482 125432 307538 125488
rect 307298 124208 307354 124264
rect 307574 125024 307630 125080
rect 307666 124616 307722 124672
rect 307574 123800 307630 123856
rect 307666 122984 307722 123040
rect 307482 122440 307538 122496
rect 307666 122032 307722 122088
rect 307574 121624 307630 121680
rect 307482 121216 307538 121272
rect 307666 120808 307722 120864
rect 307574 120400 307630 120456
rect 307482 119992 307538 120048
rect 307574 119584 307630 119640
rect 307666 119040 307722 119096
rect 307574 118768 307630 118824
rect 307574 117816 307630 117872
rect 307666 117408 307722 117464
rect 307574 117000 307630 117056
rect 307666 116184 307722 116240
rect 307482 115640 307538 115696
rect 307574 115232 307630 115288
rect 307666 114824 307722 114880
rect 307666 114416 307722 114472
rect 307574 113600 307630 113656
rect 307666 113212 307722 113248
rect 307666 113192 307668 113212
rect 307668 113192 307720 113212
rect 307720 113192 307722 113212
rect 307666 111868 307668 111888
rect 307668 111868 307720 111888
rect 307720 111868 307722 111888
rect 307666 111832 307722 111868
rect 307482 111424 307538 111480
rect 307574 111016 307630 111072
rect 307666 110608 307722 110664
rect 307666 109792 307722 109848
rect 307574 108840 307630 108896
rect 307666 108024 307722 108080
rect 307666 107616 307722 107672
rect 307574 107208 307630 107264
rect 307482 106800 307538 106856
rect 307666 106392 307722 106448
rect 307482 105440 307538 105496
rect 307666 105032 307722 105088
rect 307574 104216 307630 104272
rect 307666 103808 307722 103864
rect 307574 103400 307630 103456
rect 307666 102448 307722 102504
rect 307666 102040 307722 102096
rect 307574 101632 307630 101688
rect 307574 100000 307630 100056
rect 307666 99592 307722 99648
rect 307574 99048 307630 99104
rect 307666 98232 307722 98288
rect 307482 97824 307538 97880
rect 307666 96600 307722 96656
rect 308494 178064 308550 178120
rect 308494 123392 308550 123448
rect 307666 96192 307722 96248
rect 309138 112240 309194 112296
rect 316038 178064 316094 178120
rect 316406 178064 316462 178120
rect 319350 242528 319406 242584
rect 320270 345480 320326 345536
rect 320270 248784 320326 248840
rect 320362 246744 320418 246800
rect 321742 359352 321798 359408
rect 321650 359080 321706 359136
rect 321558 352144 321614 352200
rect 322846 354356 322848 354376
rect 322848 354356 322900 354376
rect 322900 354356 322902 354376
rect 322846 354320 322902 354356
rect 322202 352144 322258 352200
rect 322662 350104 322718 350160
rect 321834 347384 321890 347440
rect 322294 347384 322350 347440
rect 322478 343304 322534 343360
rect 322846 341400 322902 341456
rect 322478 336676 322480 336696
rect 322480 336676 322532 336696
rect 322532 336676 322534 336696
rect 322478 336640 322534 336676
rect 321742 334620 321798 334656
rect 321742 334600 321744 334620
rect 321744 334600 321796 334620
rect 321796 334600 321798 334620
rect 321650 331744 321706 331800
rect 322202 331764 322258 331800
rect 322202 331744 322204 331764
rect 322204 331744 322256 331764
rect 322256 331744 322258 331764
rect 322202 329840 322258 329896
rect 322846 327700 322848 327720
rect 322848 327700 322900 327720
rect 322900 327700 322902 327720
rect 322846 327664 322902 327700
rect 322754 324964 322810 325000
rect 322754 324944 322756 324964
rect 322756 324944 322808 324964
rect 322808 324944 322810 324964
rect 322478 322940 322480 322960
rect 322480 322940 322532 322960
rect 322532 322940 322534 322960
rect 322478 322904 322534 322940
rect 322202 320864 322258 320920
rect 322846 318844 322902 318880
rect 322846 318824 322848 318844
rect 322848 318824 322900 318844
rect 322900 318824 322902 318844
rect 322478 316240 322534 316296
rect 322478 314200 322534 314256
rect 322846 312044 322902 312080
rect 322846 312024 322848 312044
rect 322848 312024 322900 312044
rect 322900 312024 322902 312044
rect 322478 309440 322534 309496
rect 322478 307400 322534 307456
rect 322478 305224 322534 305280
rect 322478 303184 322534 303240
rect 322846 300600 322902 300656
rect 322478 298560 322534 298616
rect 322478 296384 322534 296440
rect 322846 293664 322902 293720
rect 322846 291624 322902 291680
rect 322846 289584 322902 289640
rect 321558 286864 321614 286920
rect 322202 284960 322258 285016
rect 322478 282940 322534 282976
rect 322478 282920 322480 282940
rect 322480 282920 322532 282940
rect 322532 282920 322534 282940
rect 322478 280744 322534 280800
rect 322202 278024 322258 278080
rect 321650 255584 321706 255640
rect 321742 242528 321798 242584
rect 321742 239944 321798 240000
rect 322846 276020 322848 276040
rect 322848 276020 322900 276040
rect 322900 276020 322902 276040
rect 322846 275984 322902 276020
rect 322386 274080 322442 274136
rect 322846 271224 322902 271280
rect 322846 269184 322902 269240
rect 322478 267280 322534 267336
rect 322478 265104 322534 265160
rect 322478 262384 322534 262440
rect 322570 260344 322626 260400
rect 322478 251504 322534 251560
rect 322846 244704 322902 244760
rect 318614 176160 318670 176216
rect 321466 176024 321522 176080
rect 321374 175752 321430 175808
rect 321374 173712 321430 173768
rect 321282 169632 321338 169688
rect 321650 162152 321706 162208
rect 321834 172624 321890 172680
rect 323030 338680 323086 338736
rect 322938 160792 322994 160848
rect 335542 389136 335598 389192
rect 324502 353368 324558 353424
rect 324410 311752 324466 311808
rect 323674 237224 323730 237280
rect 324410 258304 324466 258360
rect 323214 174664 323270 174720
rect 325054 237088 325110 237144
rect 324962 181464 325018 181520
rect 324410 173984 324466 174040
rect 324318 168544 324374 168600
rect 324318 167728 324374 167784
rect 324318 165416 324374 165472
rect 324410 164736 324466 164792
rect 324318 163920 324374 163976
rect 324410 163104 324466 163160
rect 324318 162424 324374 162480
rect 323122 159296 323178 159352
rect 324318 158516 324320 158536
rect 324320 158516 324372 158536
rect 324372 158516 324374 158536
rect 324318 158480 324374 158516
rect 324410 157800 324466 157856
rect 324318 156304 324374 156360
rect 323030 154672 323086 154728
rect 324318 153992 324374 154048
rect 324410 153176 324466 153232
rect 324318 152360 324374 152416
rect 324318 151700 324374 151736
rect 324318 151680 324320 151700
rect 324320 151680 324372 151700
rect 324372 151680 324374 151700
rect 324410 150864 324466 150920
rect 324318 150048 324374 150104
rect 324410 149368 324466 149424
rect 324318 148552 324374 148608
rect 324410 147736 324466 147792
rect 324318 147056 324374 147112
rect 324318 146260 324374 146296
rect 324318 146240 324320 146260
rect 324320 146240 324372 146260
rect 324372 146240 324374 146260
rect 324318 144744 324374 144800
rect 324410 143112 324466 143168
rect 324318 142432 324374 142488
rect 324318 141616 324374 141672
rect 324410 140800 324466 140856
rect 324318 138488 324374 138544
rect 324318 137844 324320 137864
rect 324320 137844 324372 137864
rect 324372 137844 324374 137864
rect 324318 137808 324374 137844
rect 324410 136992 324466 137048
rect 324318 136312 324374 136368
rect 324410 135496 324466 135552
rect 323490 134136 323546 134192
rect 323490 133864 323546 133920
rect 321742 133728 321798 133784
rect 324318 130872 324374 130928
rect 324410 130056 324466 130112
rect 321558 129648 321614 129704
rect 324318 128560 324374 128616
rect 324318 127744 324374 127800
rect 324410 127064 324466 127120
rect 324594 176160 324650 176216
rect 324594 170856 324650 170912
rect 324594 145424 324650 145480
rect 324502 126248 324558 126304
rect 324318 125468 324320 125488
rect 324320 125468 324372 125488
rect 324372 125468 324374 125488
rect 324318 125432 324374 125468
rect 324410 124752 324466 124808
rect 324318 123936 324374 123992
rect 324410 123120 324466 123176
rect 324318 122440 324374 122496
rect 324410 121624 324466 121680
rect 325606 160112 325662 160168
rect 327078 239980 327080 240000
rect 327080 239980 327132 240000
rect 327132 239980 327134 240000
rect 327078 239944 327134 239980
rect 327262 234232 327318 234288
rect 327446 234232 327502 234288
rect 324962 120808 325018 120864
rect 324318 120128 324374 120184
rect 324318 119312 324374 119368
rect 324318 118532 324320 118552
rect 324320 118532 324372 118552
rect 324372 118532 324374 118552
rect 324318 118496 324374 118532
rect 324410 117816 324466 117872
rect 324318 117000 324374 117056
rect 324410 116320 324466 116376
rect 324318 115504 324374 115560
rect 324410 114688 324466 114744
rect 324318 114008 324374 114064
rect 324410 113192 324466 113248
rect 324318 112376 324374 112432
rect 324318 111732 324320 111752
rect 324320 111732 324372 111752
rect 324372 111732 324374 111752
rect 324318 111696 324374 111732
rect 324410 110880 324466 110936
rect 324502 110064 324558 110120
rect 324318 109384 324374 109440
rect 324318 107752 324374 107808
rect 324318 107072 324374 107128
rect 322938 106256 322994 106312
rect 321834 105032 321890 105088
rect 321650 102720 321706 102776
rect 321558 99592 321614 99648
rect 321742 102176 321798 102232
rect 321466 95784 321522 95840
rect 324410 104760 324466 104816
rect 324594 108568 324650 108624
rect 324318 101632 324374 101688
rect 324318 99340 324374 99376
rect 324318 99320 324320 99340
rect 324320 99320 324372 99340
rect 324372 99320 324374 99340
rect 324502 100816 324558 100872
rect 324410 97824 324466 97880
rect 324318 97008 324374 97064
rect 308494 40568 308550 40624
rect 316038 81368 316094 81424
rect 316130 43424 316186 43480
rect 317326 43444 317382 43480
rect 317326 43424 317328 43444
rect 317328 43424 317380 43444
rect 317380 43424 317382 43444
rect 325606 104216 325662 104272
rect 325882 132368 325938 132424
rect 329838 240100 329894 240136
rect 329838 240080 329840 240100
rect 329840 240080 329892 240100
rect 329892 240080 329894 240100
rect 331218 226208 331274 226264
rect 331862 147736 331918 147792
rect 330482 26152 330538 26208
rect 329838 24928 329894 24984
rect 330482 24928 330538 24984
rect 332506 147736 332562 147792
rect 333978 234368 334034 234424
rect 332598 59880 332654 59936
rect 333978 44784 334034 44840
rect 334806 76608 334862 76664
rect 339130 77832 339186 77888
rect 340878 47540 340880 47560
rect 340880 47540 340932 47560
rect 340932 47540 340934 47560
rect 340878 47504 340934 47540
rect 343638 96328 343694 96384
rect 342350 41248 342406 41304
rect 342166 11736 342222 11792
rect 339958 8236 339960 8256
rect 339960 8236 340012 8256
rect 340012 8236 340014 8256
rect 339958 8200 340014 8236
rect 345110 177248 345166 177304
rect 345018 98640 345074 98696
rect 347962 181328 348018 181384
rect 345754 81388 345810 81424
rect 345754 81368 345756 81388
rect 345756 81368 345808 81388
rect 345808 81368 345810 81388
rect 347778 46824 347834 46880
rect 348422 46824 348478 46880
rect 353390 360304 353446 360360
rect 353942 360304 353998 360360
rect 354678 359488 354734 359544
rect 359462 361936 359518 361992
rect 362958 221448 363014 221504
rect 360198 99320 360254 99376
rect 360198 98640 360254 98696
rect 381542 95104 381598 95160
rect 416778 178608 416834 178664
rect 416778 176976 416834 177032
rect 416778 175208 416834 175264
rect 416778 171808 416834 171864
rect 416778 168428 416834 168464
rect 416778 168408 416780 168428
rect 416780 168408 416832 168428
rect 416832 168408 416834 168428
rect 416778 166776 416834 166832
rect 416778 165008 416834 165064
rect 416778 163376 416834 163432
rect 416778 161744 416834 161800
rect 416778 159976 416834 160032
rect 416778 156576 416834 156632
rect 416778 154944 416834 155000
rect 416778 153212 416780 153232
rect 416780 153212 416832 153232
rect 416832 153212 416834 153232
rect 416778 153176 416834 153212
rect 416778 151544 416834 151600
rect 416778 149776 416834 149832
rect 416778 148144 416834 148200
rect 416778 146512 416834 146568
rect 416778 144744 416834 144800
rect 416870 143112 416926 143168
rect 416778 141344 416834 141400
rect 416778 139712 416834 139768
rect 416778 137964 416834 138000
rect 416778 137944 416780 137964
rect 416780 137944 416832 137964
rect 416832 137944 416834 137964
rect 416778 136312 416834 136368
rect 417330 134544 417386 134600
rect 416778 122748 416780 122768
rect 416780 122748 416832 122768
rect 416832 122748 416834 122768
rect 416778 122712 416834 122748
rect 416778 121080 416834 121136
rect 417514 131280 417570 131336
rect 418710 127880 418766 127936
rect 419262 134544 419318 134600
rect 418802 126112 418858 126168
rect 417422 119312 417478 119368
rect 416778 117680 416834 117736
rect 416778 116048 416834 116104
rect 416778 114280 416834 114336
rect 416778 112648 416834 112704
rect 416778 110880 416834 110936
rect 416778 109248 416834 109304
rect 416778 107480 416834 107536
rect 416778 105848 416834 105904
rect 416778 104080 416834 104136
rect 416778 102448 416834 102504
rect 416778 100816 416834 100872
rect 419446 132912 419502 132968
rect 419354 127880 419410 127936
rect 543462 702480 543518 702536
rect 494058 179288 494114 179344
rect 493874 178608 493930 178664
rect 494058 168408 494114 168464
rect 419722 131280 419778 131336
rect 419630 129512 419686 129568
rect 419538 124480 419594 124536
rect 493966 100408 494022 100464
rect 494150 148960 494206 149016
rect 494150 146240 494206 146296
rect 494242 141208 494298 141264
rect 495346 140820 495402 140856
rect 495346 140800 495348 140820
rect 495348 140800 495400 140820
rect 495400 140800 495402 140820
rect 494334 132096 494390 132152
rect 499578 360168 499634 360224
rect 495530 173304 495586 173360
rect 495438 119584 495494 119640
rect 494242 104760 494298 104816
rect 495438 103808 495494 103864
rect 496910 177792 496966 177848
rect 496818 176724 496874 176760
rect 496818 176704 496820 176724
rect 496820 176704 496872 176724
rect 496872 176704 496874 176724
rect 496818 175636 496874 175672
rect 496818 175616 496820 175636
rect 496820 175616 496872 175636
rect 496872 175616 496874 175636
rect 496818 167728 496874 167784
rect 496818 166640 496874 166696
rect 496818 165416 496874 165472
rect 495714 164328 495770 164384
rect 496358 164328 496414 164384
rect 496818 163240 496874 163296
rect 496818 162152 496874 162208
rect 498106 171128 498162 171184
rect 496910 160928 496966 160984
rect 496910 159840 496966 159896
rect 497002 158752 497058 158808
rect 496910 157664 496966 157720
rect 496910 156440 496966 156496
rect 496910 155352 496966 155408
rect 496910 154264 496966 154320
rect 497002 153176 497058 153232
rect 496910 152088 496966 152144
rect 496818 150864 496874 150920
rect 496818 149776 496874 149832
rect 496818 147620 496874 147656
rect 496818 147600 496820 147620
rect 496820 147600 496872 147620
rect 496872 147600 496874 147620
rect 496818 145288 496874 145344
rect 496818 144220 496874 144256
rect 496818 144200 496820 144220
rect 496820 144200 496872 144220
rect 496872 144200 496874 144220
rect 496818 143112 496874 143168
rect 496818 141888 496874 141944
rect 496818 139712 496874 139768
rect 496818 138624 496874 138680
rect 496818 137400 496874 137456
rect 496818 136348 496820 136368
rect 496820 136348 496872 136368
rect 496872 136348 496874 136368
rect 496818 136312 496874 136348
rect 496910 135224 496966 135280
rect 496818 132912 496874 132968
rect 495622 130736 495678 130792
rect 496818 129684 496820 129704
rect 496820 129684 496872 129704
rect 496872 129684 496874 129704
rect 496818 129648 496874 129684
rect 496818 127336 496874 127392
rect 496818 126248 496874 126304
rect 496818 125160 496874 125216
rect 496910 124072 496966 124128
rect 496818 122848 496874 122904
rect 496818 121760 496874 121816
rect 496818 118360 496874 118416
rect 496910 117272 496966 117328
rect 496818 116184 496874 116240
rect 497462 115096 497518 115152
rect 496818 113872 496874 113928
rect 496910 112784 496966 112840
rect 496818 111732 496820 111752
rect 496820 111732 496872 111752
rect 496872 111732 496874 111752
rect 496818 111696 496874 111732
rect 496818 110608 496874 110664
rect 496818 109384 496874 109440
rect 496818 107208 496874 107264
rect 497002 108296 497058 108352
rect 496910 106120 496966 106176
rect 497094 101632 497150 101688
rect 498382 120672 498438 120728
rect 504086 166912 504142 166968
rect 511998 211792 512054 211848
rect 517610 218592 517666 218648
rect 580906 697176 580962 697232
rect 580170 683848 580226 683904
rect 580262 670656 580318 670712
rect 582378 670656 582434 670712
rect 580170 644000 580226 644056
rect 579802 630808 579858 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580262 587968 580318 588024
rect 580262 577632 580318 577688
rect 580170 564304 580226 564360
rect 580170 537784 580226 537840
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579618 365064 579674 365120
rect 580262 351872 580318 351928
rect 580170 325216 580226 325272
rect 580354 312024 580410 312080
rect 580262 298696 580318 298752
rect 580170 272176 580226 272232
rect 579986 258848 580042 258904
rect 580170 245520 580226 245576
rect 580170 232328 580226 232384
rect 579802 219000 579858 219056
rect 580170 205672 580226 205728
rect 580354 192480 580410 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580262 152632 580318 152688
rect 580170 139304 580226 139360
rect 580170 125976 580226 126032
rect 580262 112784 580318 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580262 33088 580318 33144
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect 81014 702612 81020 702676
rect 81084 702674 81090 702676
rect 397453 702674 397519 702677
rect 81084 702672 397519 702674
rect 81084 702616 397458 702672
rect 397514 702616 397519 702672
rect 81084 702614 397519 702616
rect 81084 702612 81090 702614
rect 397453 702611 397519 702614
rect 68870 702476 68876 702540
rect 68940 702538 68946 702540
rect 543457 702538 543523 702541
rect 68940 702536 543523 702538
rect 68940 702480 543462 702536
rect 543518 702480 543523 702536
rect 68940 702478 543523 702480
rect 68940 702476 68946 702478
rect 543457 702475 543523 702478
rect 89161 699818 89227 699821
rect 89294 699818 89300 699820
rect 89161 699816 89300 699818
rect 89161 699760 89166 699816
rect 89222 699760 89300 699816
rect 89161 699758 89300 699760
rect 89161 699755 89227 699758
rect 89294 699756 89300 699758
rect 89364 699756 89370 699820
rect -960 697220 480 697460
rect 580901 697234 580967 697237
rect 583520 697234 584960 697324
rect 580901 697232 584960 697234
rect 580901 697176 580906 697232
rect 580962 697176 584960 697232
rect 580901 697174 584960 697176
rect 580901 697171 580967 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect 70894 681804 70900 681868
rect 70964 681866 70970 681868
rect 74533 681866 74599 681869
rect 70964 681864 74599 681866
rect 70964 681808 74538 681864
rect 74594 681808 74599 681864
rect 70964 681806 74599 681808
rect 70964 681804 70970 681806
rect 74533 681803 74599 681806
rect 98545 681866 98611 681869
rect 99281 681866 99347 681869
rect 98545 681864 99347 681866
rect 98545 681808 98550 681864
rect 98606 681808 99286 681864
rect 99342 681808 99347 681864
rect 98545 681806 99347 681808
rect 98545 681803 98611 681806
rect 99281 681803 99347 681806
rect 106917 681866 106983 681869
rect 107561 681866 107627 681869
rect 106917 681864 107627 681866
rect 106917 681808 106922 681864
rect 106978 681808 107566 681864
rect 107622 681808 107627 681864
rect 106917 681806 107627 681808
rect 106917 681803 106983 681806
rect 107561 681803 107627 681806
rect 84694 680580 84700 680644
rect 84764 680642 84770 680644
rect 89069 680642 89135 680645
rect 84764 680640 89135 680642
rect 84764 680584 89074 680640
rect 89130 680584 89135 680640
rect 84764 680582 89135 680584
rect 84764 680580 84770 680582
rect 89069 680579 89135 680582
rect 72918 680444 72924 680508
rect 72988 680506 72994 680508
rect 75177 680506 75243 680509
rect 72988 680504 75243 680506
rect 72988 680448 75182 680504
rect 75238 680448 75243 680504
rect 72988 680446 75243 680448
rect 72988 680444 72994 680446
rect 75177 680443 75243 680446
rect 77150 680444 77156 680508
rect 77220 680506 77226 680508
rect 79317 680506 79383 680509
rect 77220 680504 79383 680506
rect 77220 680448 79322 680504
rect 79378 680448 79383 680504
rect 77220 680446 79383 680448
rect 77220 680444 77226 680446
rect 79317 680443 79383 680446
rect 82486 680444 82492 680508
rect 82556 680506 82562 680508
rect 84837 680506 84903 680509
rect 82556 680504 84903 680506
rect 82556 680448 84842 680504
rect 84898 680448 84903 680504
rect 82556 680446 84903 680448
rect 82556 680444 82562 680446
rect 84837 680443 84903 680446
rect 86718 680444 86724 680508
rect 86788 680506 86794 680508
rect 89713 680506 89779 680509
rect 86788 680504 89779 680506
rect 86788 680448 89718 680504
rect 89774 680448 89779 680504
rect 86788 680446 89779 680448
rect 86788 680444 86794 680446
rect 89713 680443 89779 680446
rect 99046 680444 99052 680508
rect 99116 680506 99122 680508
rect 102501 680506 102567 680509
rect 99116 680504 102567 680506
rect 99116 680448 102506 680504
rect 102562 680448 102567 680504
rect 99116 680446 102567 680448
rect 99116 680444 99122 680446
rect 102501 680443 102567 680446
rect 104566 680444 104572 680508
rect 104636 680506 104642 680508
rect 107653 680506 107719 680509
rect 104636 680504 107719 680506
rect 104636 680448 107658 680504
rect 107714 680448 107719 680504
rect 104636 680446 107719 680448
rect 104636 680444 104642 680446
rect 107653 680443 107719 680446
rect 75126 680308 75132 680372
rect 75196 680370 75202 680372
rect 77109 680370 77175 680373
rect 75196 680368 77175 680370
rect 75196 680312 77114 680368
rect 77170 680312 77175 680368
rect 75196 680310 77175 680312
rect 75196 680308 75202 680310
rect 77109 680307 77175 680310
rect 78254 680308 78260 680372
rect 78324 680370 78330 680372
rect 81617 680370 81683 680373
rect 82077 680370 82143 680373
rect 78324 680368 82143 680370
rect 78324 680312 81622 680368
rect 81678 680312 82082 680368
rect 82138 680312 82143 680368
rect 78324 680310 82143 680312
rect 78324 680308 78330 680310
rect 81617 680307 81683 680310
rect 82077 680307 82143 680310
rect 82670 680308 82676 680372
rect 82740 680370 82746 680372
rect 85481 680370 85547 680373
rect 82740 680368 85547 680370
rect 82740 680312 85486 680368
rect 85542 680312 85547 680368
rect 82740 680310 85547 680312
rect 82740 680308 82746 680310
rect 85481 680307 85547 680310
rect 88926 680308 88932 680372
rect 88996 680370 89002 680372
rect 91921 680370 91987 680373
rect 88996 680368 91987 680370
rect 88996 680312 91926 680368
rect 91982 680312 91987 680368
rect 88996 680310 91987 680312
rect 88996 680308 89002 680310
rect 91921 680307 91987 680310
rect 101990 680308 101996 680372
rect 102060 680370 102066 680372
rect 104801 680370 104867 680373
rect 102060 680368 104867 680370
rect 102060 680312 104806 680368
rect 104862 680312 104867 680368
rect 102060 680310 104867 680312
rect 102060 680308 102066 680310
rect 104801 680307 104867 680310
rect 70393 679828 70459 679829
rect 70342 679826 70348 679828
rect 70302 679766 70348 679826
rect 70412 679824 70459 679828
rect 70454 679768 70459 679824
rect 70342 679764 70348 679766
rect 70412 679764 70459 679768
rect 100518 679764 100524 679828
rect 100588 679826 100594 679828
rect 103329 679826 103395 679829
rect 100588 679824 103395 679826
rect 100588 679768 103334 679824
rect 103390 679768 103395 679824
rect 100588 679766 103395 679768
rect 100588 679764 100594 679766
rect 70393 679763 70459 679764
rect 103329 679763 103395 679766
rect 92238 679628 92244 679692
rect 92308 679690 92314 679692
rect 94865 679690 94931 679693
rect 92308 679688 94931 679690
rect 92308 679632 94870 679688
rect 94926 679632 94931 679688
rect 92308 679630 94931 679632
rect 92308 679628 92314 679630
rect 94865 679627 94931 679630
rect 94998 679628 95004 679692
rect 95068 679690 95074 679692
rect 96797 679690 96863 679693
rect 95068 679688 96863 679690
rect 95068 679632 96802 679688
rect 96858 679632 96863 679688
rect 95068 679630 96863 679632
rect 95068 679628 95074 679630
rect 96797 679627 96863 679630
rect 97758 679628 97764 679692
rect 97828 679690 97834 679692
rect 100661 679690 100727 679693
rect 97828 679688 100727 679690
rect 97828 679632 100666 679688
rect 100722 679632 100727 679688
rect 97828 679630 100727 679632
rect 97828 679628 97834 679630
rect 100661 679627 100727 679630
rect 104750 679628 104756 679692
rect 104820 679690 104826 679692
rect 108389 679690 108455 679693
rect 104820 679688 108455 679690
rect 104820 679632 108394 679688
rect 108450 679632 108455 679688
rect 104820 679630 108455 679632
rect 104820 679628 104826 679630
rect 108389 679627 108455 679630
rect 79174 679492 79180 679556
rect 79244 679554 79250 679556
rect 81893 679554 81959 679557
rect 79244 679552 81959 679554
rect 79244 679496 81898 679552
rect 81954 679496 81959 679552
rect 79244 679494 81959 679496
rect 79244 679492 79250 679494
rect 81893 679491 81959 679494
rect 83958 679492 83964 679556
rect 84028 679554 84034 679556
rect 85757 679554 85823 679557
rect 84028 679552 85823 679554
rect 84028 679496 85762 679552
rect 85818 679496 85823 679552
rect 84028 679494 85823 679496
rect 84028 679492 84034 679494
rect 85757 679491 85823 679494
rect 90950 679492 90956 679556
rect 91020 679554 91026 679556
rect 92933 679554 92999 679557
rect 91020 679552 92999 679554
rect 91020 679496 92938 679552
rect 92994 679496 92999 679552
rect 91020 679494 92999 679496
rect 91020 679492 91026 679494
rect 92933 679491 92999 679494
rect 93710 679492 93716 679556
rect 93780 679554 93786 679556
rect 96153 679554 96219 679557
rect 93780 679552 96219 679554
rect 93780 679496 96158 679552
rect 96214 679496 96219 679552
rect 93780 679494 96219 679496
rect 93780 679492 93786 679494
rect 96153 679491 96219 679494
rect 96470 679492 96476 679556
rect 96540 679554 96546 679556
rect 99373 679554 99439 679557
rect 96540 679552 99439 679554
rect 96540 679496 99378 679552
rect 99434 679496 99439 679552
rect 96540 679494 99439 679496
rect 96540 679492 96546 679494
rect 99373 679491 99439 679494
rect 103278 679492 103284 679556
rect 103348 679554 103354 679556
rect 105813 679554 105879 679557
rect 103348 679552 105879 679554
rect 103348 679496 105818 679552
rect 105874 679496 105879 679552
rect 103348 679494 105879 679496
rect 103348 679492 103354 679494
rect 105813 679491 105879 679494
rect 106774 679492 106780 679556
rect 106844 679554 106850 679556
rect 106917 679554 106983 679557
rect 106844 679552 106983 679554
rect 106844 679496 106922 679552
rect 106978 679496 106983 679552
rect 106844 679494 106983 679496
rect 106844 679492 106850 679494
rect 106917 679491 106983 679494
rect 71773 679420 71839 679421
rect 71773 679416 71820 679420
rect 71884 679418 71890 679420
rect 67541 679146 67607 679149
rect 70166 679146 70226 679388
rect 71773 679360 71778 679416
rect 71773 679356 71820 679360
rect 71884 679358 71930 679418
rect 71884 679356 71890 679358
rect 73102 679356 73108 679420
rect 73172 679418 73178 679420
rect 73613 679418 73679 679421
rect 73172 679416 73679 679418
rect 73172 679360 73618 679416
rect 73674 679360 73679 679416
rect 73172 679358 73679 679360
rect 73172 679356 73178 679358
rect 71773 679355 71839 679356
rect 73613 679355 73679 679358
rect 74758 679356 74764 679420
rect 74828 679418 74834 679420
rect 75453 679418 75519 679421
rect 74828 679416 75519 679418
rect 74828 679360 75458 679416
rect 75514 679360 75519 679416
rect 74828 679358 75519 679360
rect 74828 679356 74834 679358
rect 75453 679355 75519 679358
rect 75862 679356 75868 679420
rect 75932 679418 75938 679420
rect 76189 679418 76255 679421
rect 75932 679416 76255 679418
rect 75932 679360 76194 679416
rect 76250 679360 76255 679416
rect 75932 679358 76255 679360
rect 75932 679356 75938 679358
rect 76189 679355 76255 679358
rect 78121 679418 78187 679421
rect 78857 679420 78923 679421
rect 80145 679420 80211 679421
rect 78438 679418 78444 679420
rect 78121 679416 78444 679418
rect 78121 679360 78126 679416
rect 78182 679360 78444 679416
rect 78121 679358 78444 679360
rect 78121 679355 78187 679358
rect 78438 679356 78444 679358
rect 78508 679356 78514 679420
rect 78806 679418 78812 679420
rect 78766 679358 78812 679418
rect 78876 679416 78923 679420
rect 80094 679418 80100 679420
rect 78918 679360 78923 679416
rect 78806 679356 78812 679358
rect 78876 679356 78923 679360
rect 80054 679358 80100 679418
rect 80164 679416 80211 679420
rect 80206 679360 80211 679416
rect 80094 679356 80100 679358
rect 80164 679356 80211 679360
rect 78857 679355 78923 679356
rect 80145 679355 80211 679356
rect 82721 679418 82787 679421
rect 84469 679420 84535 679421
rect 82854 679418 82860 679420
rect 82721 679416 82860 679418
rect 82721 679360 82726 679416
rect 82782 679360 82860 679416
rect 82721 679358 82860 679360
rect 82721 679355 82787 679358
rect 82854 679356 82860 679358
rect 82924 679356 82930 679420
rect 84469 679416 84516 679420
rect 84580 679418 84586 679420
rect 84469 679360 84474 679416
rect 84469 679356 84516 679360
rect 84580 679358 84626 679418
rect 84580 679356 84586 679358
rect 85798 679356 85804 679420
rect 85868 679418 85874 679420
rect 86493 679418 86559 679421
rect 87137 679420 87203 679421
rect 87086 679418 87092 679420
rect 85868 679416 86559 679418
rect 85868 679360 86498 679416
rect 86554 679360 86559 679416
rect 85868 679358 86559 679360
rect 87046 679358 87092 679418
rect 87156 679416 87203 679420
rect 87198 679360 87203 679416
rect 85868 679356 85874 679358
rect 84469 679355 84535 679356
rect 86493 679355 86559 679358
rect 87086 679356 87092 679358
rect 87156 679356 87203 679360
rect 87270 679356 87276 679420
rect 87340 679418 87346 679420
rect 87781 679418 87847 679421
rect 87340 679416 87847 679418
rect 87340 679360 87786 679416
rect 87842 679360 87847 679416
rect 87340 679358 87847 679360
rect 87340 679356 87346 679358
rect 87137 679355 87203 679356
rect 87781 679355 87847 679358
rect 91461 679420 91527 679421
rect 91461 679416 91508 679420
rect 91572 679418 91578 679420
rect 91461 679360 91466 679416
rect 91461 679356 91508 679360
rect 91572 679358 91618 679418
rect 91572 679356 91578 679358
rect 92606 679356 92612 679420
rect 92676 679418 92682 679420
rect 92749 679418 92815 679421
rect 92676 679416 92815 679418
rect 92676 679360 92754 679416
rect 92810 679360 92815 679416
rect 92676 679358 92815 679360
rect 92676 679356 92682 679358
rect 91461 679355 91527 679356
rect 92749 679355 92815 679358
rect 94078 679356 94084 679420
rect 94148 679418 94154 679420
rect 94221 679418 94287 679421
rect 94148 679416 94287 679418
rect 94148 679360 94226 679416
rect 94282 679360 94287 679416
rect 94148 679358 94287 679360
rect 94148 679356 94154 679358
rect 94221 679355 94287 679358
rect 96153 679418 96219 679421
rect 96286 679418 96292 679420
rect 96153 679416 96292 679418
rect 96153 679360 96158 679416
rect 96214 679360 96292 679416
rect 96153 679358 96292 679360
rect 96153 679355 96219 679358
rect 96286 679356 96292 679358
rect 96356 679356 96362 679420
rect 97206 679356 97212 679420
rect 97276 679418 97282 679420
rect 97349 679418 97415 679421
rect 98545 679420 98611 679421
rect 100017 679420 100083 679421
rect 101305 679420 101371 679421
rect 97276 679416 97415 679418
rect 97276 679360 97354 679416
rect 97410 679360 97415 679416
rect 97276 679358 97415 679360
rect 97276 679356 97282 679358
rect 97349 679355 97415 679358
rect 98494 679356 98500 679420
rect 98564 679418 98611 679420
rect 99966 679418 99972 679420
rect 98564 679416 98656 679418
rect 98606 679360 98656 679416
rect 98564 679358 98656 679360
rect 99926 679358 99972 679418
rect 100036 679416 100083 679420
rect 101254 679418 101260 679420
rect 100078 679360 100083 679416
rect 98564 679356 98611 679358
rect 99966 679356 99972 679358
rect 100036 679356 100083 679360
rect 101214 679358 101260 679418
rect 101324 679416 101371 679420
rect 101366 679360 101371 679416
rect 101254 679356 101260 679358
rect 101324 679356 101371 679360
rect 98545 679355 98611 679356
rect 100017 679355 100083 679356
rect 101305 679355 101371 679356
rect 102593 679418 102659 679421
rect 102726 679418 102732 679420
rect 102593 679416 102732 679418
rect 102593 679360 102598 679416
rect 102654 679360 102732 679416
rect 102593 679358 102732 679360
rect 102593 679355 102659 679358
rect 102726 679356 102732 679358
rect 102796 679356 102802 679420
rect 105486 679356 105492 679420
rect 105556 679418 105562 679420
rect 105629 679418 105695 679421
rect 105556 679416 105695 679418
rect 105556 679360 105634 679416
rect 105690 679360 105695 679416
rect 105556 679358 105695 679360
rect 105556 679356 105562 679358
rect 105629 679355 105695 679358
rect 106958 679356 106964 679420
rect 107028 679418 107034 679420
rect 107101 679418 107167 679421
rect 107028 679416 107167 679418
rect 107028 679360 107106 679416
rect 107162 679360 107167 679416
rect 107028 679358 107167 679360
rect 107028 679356 107034 679358
rect 107101 679355 107167 679358
rect 67541 679144 70226 679146
rect 67541 679088 67546 679144
rect 67602 679088 70226 679144
rect 67541 679086 70226 679088
rect 67541 679083 67607 679086
rect 111793 678738 111859 678741
rect 109940 678736 111859 678738
rect 67633 678194 67699 678197
rect 70166 678194 70226 678708
rect 109940 678680 111798 678736
rect 111854 678680 111859 678736
rect 109940 678678 111859 678680
rect 111793 678675 111859 678678
rect 67633 678192 70226 678194
rect 67633 678136 67638 678192
rect 67694 678136 70226 678192
rect 67633 678134 70226 678136
rect 67633 678131 67699 678134
rect 112345 678058 112411 678061
rect 109940 678056 112411 678058
rect 109940 678000 112350 678056
rect 112406 678000 112411 678056
rect 109940 677998 112411 678000
rect 112345 677995 112411 677998
rect 111793 677378 111859 677381
rect 109940 677376 111859 677378
rect 68737 677106 68803 677109
rect 70166 677106 70226 677348
rect 109940 677320 111798 677376
rect 111854 677320 111859 677376
rect 109940 677318 111859 677320
rect 111793 677315 111859 677318
rect 68737 677104 70226 677106
rect 68737 677048 68742 677104
rect 68798 677048 70226 677104
rect 68737 677046 70226 677048
rect 68737 677043 68803 677046
rect 112713 676698 112779 676701
rect 109940 676696 112779 676698
rect 67633 676426 67699 676429
rect 70166 676426 70226 676668
rect 109940 676640 112718 676696
rect 112774 676640 112779 676696
rect 109940 676638 112779 676640
rect 112713 676635 112779 676638
rect 67633 676424 70226 676426
rect 67633 676368 67638 676424
rect 67694 676368 70226 676424
rect 67633 676366 70226 676368
rect 67633 676363 67699 676366
rect 113081 676290 113147 676293
rect 118734 676290 118740 676292
rect 113081 676288 118740 676290
rect 113081 676232 113086 676288
rect 113142 676232 118740 676288
rect 113081 676230 118740 676232
rect 113081 676227 113147 676230
rect 118734 676228 118740 676230
rect 118804 676228 118810 676292
rect 111977 676018 112043 676021
rect 109940 676016 112043 676018
rect 67449 675746 67515 675749
rect 70166 675746 70226 675988
rect 109940 675960 111982 676016
rect 112038 675960 112043 676016
rect 109940 675958 112043 675960
rect 111977 675955 112043 675958
rect 67449 675744 70226 675746
rect 67449 675688 67454 675744
rect 67510 675688 70226 675744
rect 67449 675686 70226 675688
rect 67449 675683 67515 675686
rect 113081 675474 113147 675477
rect 109940 675472 113147 675474
rect 109940 675416 113086 675472
rect 113142 675416 113147 675472
rect 109940 675414 113147 675416
rect 113081 675411 113147 675414
rect 67633 675202 67699 675205
rect 70166 675202 70226 675308
rect 67633 675200 70226 675202
rect 67633 675144 67638 675200
rect 67694 675144 70226 675200
rect 67633 675142 70226 675144
rect 67633 675139 67699 675142
rect 112069 674658 112135 674661
rect 109940 674656 112135 674658
rect 67633 674386 67699 674389
rect 70166 674386 70226 674628
rect 109940 674600 112074 674656
rect 112130 674600 112135 674656
rect 109940 674598 112135 674600
rect 112069 674595 112135 674598
rect 67633 674384 70226 674386
rect 67633 674328 67638 674384
rect 67694 674328 70226 674384
rect 67633 674326 70226 674328
rect 67633 674323 67699 674326
rect 67725 673842 67791 673845
rect 70166 673842 70226 673948
rect 67725 673840 70226 673842
rect 67725 673784 67730 673840
rect 67786 673784 70226 673840
rect 67725 673782 70226 673784
rect 67725 673779 67791 673782
rect 68870 673100 68876 673164
rect 68940 673162 68946 673164
rect 70166 673162 70226 673268
rect 68940 673102 70226 673162
rect 68940 673100 68946 673102
rect 109910 673026 109970 673268
rect 115974 673026 115980 673028
rect 109910 672966 115980 673026
rect 115974 672964 115980 672966
rect 116044 672964 116050 673028
rect 110413 672618 110479 672621
rect 109940 672616 110479 672618
rect 109940 672560 110418 672616
rect 110474 672560 110479 672616
rect 109940 672558 110479 672560
rect 110413 672555 110479 672558
rect 66662 672148 66668 672212
rect 66732 672210 66738 672212
rect 68870 672210 68876 672212
rect 66732 672150 68876 672210
rect 66732 672148 66738 672150
rect 68870 672148 68876 672150
rect 68940 672148 68946 672212
rect 68645 671802 68711 671805
rect 70166 671802 70226 671908
rect 68645 671800 70226 671802
rect 68645 671744 68650 671800
rect 68706 671744 70226 671800
rect 68645 671742 70226 671744
rect 109542 671802 109602 671908
rect 111793 671802 111859 671805
rect 109542 671800 111859 671802
rect 109542 671744 111798 671800
rect 111854 671744 111859 671800
rect 109542 671742 111859 671744
rect 68645 671739 68711 671742
rect 109542 671668 109602 671742
rect 111793 671739 111859 671742
rect 109534 671604 109540 671668
rect 109604 671604 109610 671668
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect 111793 671258 111859 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect 109940 671256 111859 671258
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 67633 670986 67699 670989
rect 70166 670986 70226 671228
rect 109940 671200 111798 671256
rect 111854 671200 111859 671256
rect 109940 671198 111859 671200
rect 111793 671195 111859 671198
rect 67633 670984 70226 670986
rect 67633 670928 67638 670984
rect 67694 670928 70226 670984
rect 67633 670926 70226 670928
rect 67633 670923 67699 670926
rect 580257 670714 580323 670717
rect 582373 670714 582439 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 582378 670712
rect 582434 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 582373 670651 582439 670654
rect 111793 670578 111859 670581
rect 109940 670576 111859 670578
rect 67633 670306 67699 670309
rect 70166 670306 70226 670548
rect 109940 670520 111798 670576
rect 111854 670520 111859 670576
rect 583520 670564 584960 670654
rect 109940 670518 111859 670520
rect 111793 670515 111859 670518
rect 67633 670304 70226 670306
rect 67633 670248 67638 670304
rect 67694 670248 70226 670304
rect 67633 670246 70226 670248
rect 67633 670243 67699 670246
rect 112713 669898 112779 669901
rect 109940 669896 112779 669898
rect 67725 669626 67791 669629
rect 70166 669626 70226 669868
rect 109940 669840 112718 669896
rect 112774 669840 112779 669896
rect 109940 669838 112779 669840
rect 112713 669835 112779 669838
rect 67725 669624 70226 669626
rect 67725 669568 67730 669624
rect 67786 669568 70226 669624
rect 67725 669566 70226 669568
rect 67725 669563 67791 669566
rect 67817 669354 67883 669357
rect 69982 669354 70226 669388
rect 111793 669354 111859 669357
rect 67817 669352 70226 669354
rect 67817 669296 67822 669352
rect 67878 669328 70226 669352
rect 67878 669296 70042 669328
rect 70166 669324 70226 669328
rect 109940 669352 111859 669354
rect 67817 669294 70042 669296
rect 109940 669296 111798 669352
rect 111854 669296 111859 669352
rect 109940 669294 111859 669296
rect 67817 669291 67883 669294
rect 111793 669291 111859 669294
rect 67817 668266 67883 668269
rect 70166 668266 70226 668508
rect 67817 668264 70226 668266
rect 67817 668208 67822 668264
rect 67878 668208 70226 668264
rect 67817 668206 70226 668208
rect 67817 668203 67883 668206
rect 44030 668068 44036 668132
rect 44100 668130 44106 668132
rect 44100 668070 64890 668130
rect 44100 668068 44106 668070
rect 64830 667994 64890 668070
rect 64830 667934 70042 667994
rect 69982 667722 70042 667934
rect 70166 667722 70226 667828
rect 109358 667724 109418 667828
rect 69982 667662 70226 667722
rect 109350 667660 109356 667724
rect 109420 667660 109426 667724
rect 111977 667178 112043 667181
rect 109940 667176 112043 667178
rect 109940 667120 111982 667176
rect 112038 667120 112043 667176
rect 109940 667118 112043 667120
rect 111977 667115 112043 667118
rect 67633 666906 67699 666909
rect 67633 666904 70410 666906
rect 67633 666848 67638 666904
rect 67694 666848 70410 666904
rect 67633 666846 70410 666848
rect 67633 666843 67699 666846
rect 70350 666604 70410 666846
rect 111793 666634 111859 666637
rect 109940 666632 111859 666634
rect 109940 666576 111798 666632
rect 111854 666576 111859 666632
rect 109940 666574 111859 666576
rect 111793 666571 111859 666574
rect 110505 665818 110571 665821
rect 109940 665816 110571 665818
rect 67725 665546 67791 665549
rect 70166 665546 70226 665788
rect 109940 665760 110510 665816
rect 110566 665760 110571 665816
rect 109940 665758 110571 665760
rect 110505 665755 110571 665758
rect 67725 665544 70226 665546
rect 67725 665488 67730 665544
rect 67786 665488 70226 665544
rect 67725 665486 70226 665488
rect 67725 665483 67791 665486
rect 67633 665274 67699 665277
rect 111793 665274 111859 665277
rect 67633 665272 70042 665274
rect 67633 665216 67638 665272
rect 67694 665216 70042 665272
rect 67633 665214 70042 665216
rect 109940 665272 111859 665274
rect 109940 665216 111798 665272
rect 111854 665216 111859 665272
rect 109940 665214 111859 665216
rect 67633 665211 67699 665214
rect 69982 665002 70042 665214
rect 111793 665211 111859 665214
rect 70166 665002 70226 665108
rect 69982 664942 70226 665002
rect 112345 664458 112411 664461
rect 109940 664456 112411 664458
rect 67725 664186 67791 664189
rect 70166 664186 70226 664428
rect 109940 664400 112350 664456
rect 112406 664400 112411 664456
rect 109940 664398 112411 664400
rect 112345 664395 112411 664398
rect 67725 664184 70226 664186
rect 67725 664128 67730 664184
rect 67786 664128 70226 664184
rect 67725 664126 70226 664128
rect 67725 664123 67791 664126
rect 67633 663914 67699 663917
rect 111793 663914 111859 663917
rect 67633 663912 70042 663914
rect 67633 663856 67638 663912
rect 67694 663856 70042 663912
rect 109940 663912 111859 663914
rect 67633 663854 70042 663856
rect 67633 663851 67699 663854
rect 69982 663810 70042 663854
rect 70166 663810 70226 663884
rect 109940 663856 111798 663912
rect 111854 663856 111859 663912
rect 109940 663854 111859 663856
rect 111793 663851 111859 663854
rect 69982 663750 70226 663810
rect 67633 662962 67699 662965
rect 70166 662962 70226 663068
rect 67633 662960 70226 662962
rect 67633 662904 67638 662960
rect 67694 662904 70226 662960
rect 67633 662902 70226 662904
rect 67633 662899 67699 662902
rect 64830 662766 70410 662826
rect 61878 662628 61884 662692
rect 61948 662690 61954 662692
rect 64830 662690 64890 662766
rect 61948 662630 64890 662690
rect 61948 662628 61954 662630
rect 70350 662524 70410 662766
rect 111793 662554 111859 662557
rect 109940 662552 111859 662554
rect 109940 662496 111798 662552
rect 111854 662496 111859 662552
rect 109940 662494 111859 662496
rect 111793 662491 111859 662494
rect 111190 661738 111196 661740
rect 109940 661678 111196 661738
rect 111190 661676 111196 661678
rect 111260 661676 111266 661740
rect 67633 661466 67699 661469
rect 67633 661464 70410 661466
rect 67633 661408 67638 661464
rect 67694 661408 70410 661464
rect 67633 661406 70410 661408
rect 67633 661403 67699 661406
rect 70350 661164 70410 661406
rect 111149 661194 111215 661197
rect 109940 661192 111215 661194
rect 109940 661136 111154 661192
rect 111210 661136 111215 661192
rect 109940 661134 111215 661136
rect 111149 661131 111215 661134
rect 112345 660378 112411 660381
rect 109940 660376 112411 660378
rect 67725 660106 67791 660109
rect 70166 660106 70226 660348
rect 109940 660320 112350 660376
rect 112406 660320 112411 660376
rect 109940 660318 112411 660320
rect 112345 660315 112411 660318
rect 67725 660104 70226 660106
rect 67725 660048 67730 660104
rect 67786 660048 70226 660104
rect 67725 660046 70226 660048
rect 67725 660043 67791 660046
rect 112529 659834 112595 659837
rect 109940 659832 112595 659834
rect 109940 659776 112534 659832
rect 112590 659776 112595 659832
rect 109940 659774 112595 659776
rect 112529 659771 112595 659774
rect 67633 659698 67699 659701
rect 67633 659696 70042 659698
rect 67633 659640 67638 659696
rect 67694 659670 70042 659696
rect 67694 659640 70226 659670
rect 67633 659638 70226 659640
rect 67633 659635 67699 659638
rect 69982 659610 70226 659638
rect 111793 659018 111859 659021
rect 109940 659016 111859 659018
rect 68553 658882 68619 658885
rect 70166 658882 70226 658988
rect 109940 658960 111798 659016
rect 111854 658960 111859 659016
rect 109940 658958 111859 658960
rect 111793 658955 111859 658958
rect 68553 658880 70226 658882
rect 68553 658824 68558 658880
rect 68614 658824 70226 658880
rect 68553 658822 70226 658824
rect 68553 658819 68619 658822
rect 67633 658746 67699 658749
rect 67633 658744 70410 658746
rect 67633 658688 67638 658744
rect 67694 658688 70410 658744
rect 67633 658686 70410 658688
rect 67633 658683 67699 658686
rect 70350 658444 70410 658686
rect 110597 658474 110663 658477
rect 109940 658472 110663 658474
rect 109940 658416 110602 658472
rect 110658 658416 110663 658472
rect 109940 658414 110663 658416
rect 110597 658411 110663 658414
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 67725 657386 67791 657389
rect 70166 657386 70226 657628
rect 67725 657384 70226 657386
rect 67725 657328 67730 657384
rect 67786 657328 70226 657384
rect 67725 657326 70226 657328
rect 67725 657323 67791 657326
rect 583520 657236 584960 657476
rect 112529 656978 112595 656981
rect 109940 656976 112595 656978
rect 68185 656706 68251 656709
rect 70350 656706 70410 656948
rect 109940 656920 112534 656976
rect 112590 656920 112595 656976
rect 109940 656918 112595 656920
rect 112529 656915 112595 656918
rect 68185 656704 70410 656706
rect 68185 656648 68190 656704
rect 68246 656648 70410 656704
rect 68185 656646 70410 656648
rect 68185 656643 68251 656646
rect 112345 656298 112411 656301
rect 109940 656296 112411 656298
rect 109940 656240 112350 656296
rect 112406 656240 112411 656296
rect 109940 656238 112411 656240
rect 112345 656235 112411 656238
rect 67633 656026 67699 656029
rect 67633 656024 70410 656026
rect 67633 655968 67638 656024
rect 67694 655968 70410 656024
rect 67633 655966 70410 655968
rect 67633 655963 67699 655966
rect 70350 655724 70410 655966
rect 112529 655618 112595 655621
rect 109940 655616 112595 655618
rect 109940 655560 112534 655616
rect 112590 655560 112595 655616
rect 109940 655558 112595 655560
rect 112529 655555 112595 655558
rect 111885 654938 111951 654941
rect 109940 654936 111951 654938
rect 67633 654802 67699 654805
rect 68921 654802 68987 654805
rect 70166 654802 70226 654908
rect 109940 654880 111890 654936
rect 111946 654880 111951 654936
rect 109940 654878 111951 654880
rect 111885 654875 111951 654878
rect 67633 654800 70226 654802
rect 67633 654744 67638 654800
rect 67694 654744 68926 654800
rect 68982 654744 70226 654800
rect 67633 654742 70226 654744
rect 67633 654739 67699 654742
rect 68921 654739 68987 654742
rect 110597 654258 110663 654261
rect 109940 654256 110663 654258
rect 68686 653924 68692 653988
rect 68756 653986 68762 653988
rect 70166 653986 70226 654228
rect 109940 654200 110602 654256
rect 110658 654200 110663 654256
rect 109940 654198 110663 654200
rect 110597 654195 110663 654198
rect 68756 653926 70226 653986
rect 68756 653924 68762 653926
rect 111926 653578 111932 653580
rect 67725 653306 67791 653309
rect 70166 653306 70226 653548
rect 109940 653518 111932 653578
rect 111926 653516 111932 653518
rect 111996 653516 112002 653580
rect 67725 653304 70226 653306
rect 67725 653248 67730 653304
rect 67786 653248 70226 653304
rect 67725 653246 70226 653248
rect 67725 653243 67791 653246
rect 113081 652898 113147 652901
rect 109940 652896 113147 652898
rect 67909 652762 67975 652765
rect 70166 652762 70226 652868
rect 109940 652840 113086 652896
rect 113142 652840 113147 652896
rect 109940 652838 113147 652840
rect 113081 652835 113147 652838
rect 67909 652760 70226 652762
rect 67909 652704 67914 652760
rect 67970 652704 70226 652760
rect 67909 652702 70226 652704
rect 67909 652699 67975 652702
rect 67633 651946 67699 651949
rect 70166 651946 70226 652188
rect 67633 651944 70226 651946
rect 67633 651888 67638 651944
rect 67694 651888 70226 651944
rect 67633 651886 70226 651888
rect 67633 651883 67699 651886
rect 112529 651538 112595 651541
rect 109940 651536 112595 651538
rect 68829 651402 68895 651405
rect 70166 651402 70226 651508
rect 109940 651480 112534 651536
rect 112590 651480 112595 651536
rect 109940 651478 112595 651480
rect 112529 651475 112595 651478
rect 68829 651400 70226 651402
rect 68829 651344 68834 651400
rect 68890 651344 70226 651400
rect 68829 651342 70226 651344
rect 68829 651339 68895 651342
rect 112069 650858 112135 650861
rect 109940 650856 112135 650858
rect 109940 650800 112074 650856
rect 112130 650800 112135 650856
rect 109940 650798 112135 650800
rect 112069 650795 112135 650798
rect 111977 650178 112043 650181
rect 109940 650176 112043 650178
rect 67633 650042 67699 650045
rect 70166 650042 70226 650148
rect 109940 650120 111982 650176
rect 112038 650120 112043 650176
rect 109940 650118 112043 650120
rect 111977 650115 112043 650118
rect 67633 650040 70226 650042
rect 67633 649984 67638 650040
rect 67694 649984 70226 650040
rect 67633 649982 70226 649984
rect 67633 649979 67699 649982
rect 113081 649498 113147 649501
rect 109940 649496 113147 649498
rect 67633 649226 67699 649229
rect 70166 649226 70226 649468
rect 109940 649440 113086 649496
rect 113142 649440 113147 649496
rect 109940 649438 113147 649440
rect 113081 649435 113147 649438
rect 67633 649224 70226 649226
rect 67633 649168 67638 649224
rect 67694 649168 70226 649224
rect 67633 649166 70226 649168
rect 67633 649163 67699 649166
rect 112989 648818 113055 648821
rect 109940 648816 113055 648818
rect 68870 648620 68876 648684
rect 68940 648682 68946 648684
rect 70166 648682 70226 648788
rect 109940 648760 112994 648816
rect 113050 648760 113055 648816
rect 109940 648758 113055 648760
rect 112989 648755 113055 648758
rect 68940 648622 70226 648682
rect 68940 648620 68946 648622
rect 111977 648138 112043 648141
rect 109940 648136 112043 648138
rect 67725 647866 67791 647869
rect 70166 647866 70226 648108
rect 109940 648080 111982 648136
rect 112038 648080 112043 648136
rect 109940 648078 112043 648080
rect 111977 648075 112043 648078
rect 67725 647864 70226 647866
rect 67725 647808 67730 647864
rect 67786 647808 70226 647864
rect 67725 647806 70226 647808
rect 67725 647803 67791 647806
rect 113081 647458 113147 647461
rect 109940 647456 113147 647458
rect 67633 647322 67699 647325
rect 70166 647322 70226 647428
rect 109940 647400 113086 647456
rect 113142 647400 113147 647456
rect 109940 647398 113147 647400
rect 113081 647395 113147 647398
rect 67633 647320 70226 647322
rect 67633 647264 67638 647320
rect 67694 647264 70226 647320
rect 67633 647262 70226 647264
rect 67633 647259 67699 647262
rect 67633 646506 67699 646509
rect 70166 646506 70226 646748
rect 67633 646504 70226 646506
rect 67633 646448 67638 646504
rect 67694 646448 70226 646504
rect 67633 646446 70226 646448
rect 67633 646443 67699 646446
rect 66110 645900 66116 645964
rect 66180 645962 66186 645964
rect 70166 645962 70226 646068
rect 109358 645965 109418 646068
rect 66180 645902 70226 645962
rect 109309 645960 109418 645965
rect 109309 645904 109314 645960
rect 109370 645904 109418 645960
rect 109309 645902 109418 645904
rect 66180 645900 66186 645902
rect 109309 645899 109375 645902
rect 112989 645418 113055 645421
rect 109940 645416 113055 645418
rect 109940 645360 112994 645416
rect 113050 645360 113055 645416
rect 109940 645358 113055 645360
rect 112989 645355 113055 645358
rect -960 644996 480 645236
rect 113081 644738 113147 644741
rect 109940 644736 113147 644738
rect 68921 644602 68987 644605
rect 70166 644602 70226 644708
rect 109940 644680 113086 644736
rect 113142 644680 113147 644736
rect 109940 644678 113147 644680
rect 113081 644675 113147 644678
rect 68921 644600 70226 644602
rect 68921 644544 68926 644600
rect 68982 644544 70226 644600
rect 68921 644542 70226 644544
rect 68921 644539 68987 644542
rect 115289 644466 115355 644469
rect 115790 644466 115796 644468
rect 115289 644464 115796 644466
rect 115289 644408 115294 644464
rect 115350 644408 115796 644464
rect 115289 644406 115796 644408
rect 115289 644403 115355 644406
rect 115790 644404 115796 644406
rect 115860 644404 115866 644468
rect 111742 644058 111748 644060
rect 68553 643786 68619 643789
rect 70166 643786 70226 644028
rect 109940 643998 111748 644058
rect 111742 643996 111748 643998
rect 111812 643996 111818 644060
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect 68553 643784 70226 643786
rect 68553 643728 68558 643784
rect 68614 643728 70226 643784
rect 68553 643726 70226 643728
rect 68553 643723 68619 643726
rect 112805 643514 112871 643517
rect 109940 643512 112871 643514
rect 109940 643456 112810 643512
rect 112866 643456 112871 643512
rect 109940 643454 112871 643456
rect 112805 643451 112871 643454
rect 57830 643180 57836 643244
rect 57900 643242 57906 643244
rect 69197 643242 69263 643245
rect 70166 643242 70226 643348
rect 57900 643240 70226 643242
rect 57900 643184 69202 643240
rect 69258 643184 70226 643240
rect 57900 643182 70226 643184
rect 57900 643180 57906 643182
rect 69197 643179 69263 643182
rect 113081 642698 113147 642701
rect 109940 642696 113147 642698
rect 67725 642426 67791 642429
rect 70166 642426 70226 642668
rect 109940 642640 113086 642696
rect 113142 642640 113147 642696
rect 109940 642638 113147 642640
rect 113081 642635 113147 642638
rect 67725 642424 70226 642426
rect 67725 642368 67730 642424
rect 67786 642368 70226 642424
rect 67725 642366 70226 642368
rect 67725 642363 67791 642366
rect 112621 642154 112687 642157
rect 109940 642152 112687 642154
rect 109940 642096 112626 642152
rect 112682 642096 112687 642152
rect 109940 642094 112687 642096
rect 112621 642091 112687 642094
rect 67633 641882 67699 641885
rect 70166 641882 70226 641988
rect 67633 641880 70226 641882
rect 67633 641824 67638 641880
rect 67694 641824 70226 641880
rect 67633 641822 70226 641824
rect 67633 641819 67699 641822
rect 67725 641066 67791 641069
rect 70166 641066 70226 641308
rect 67725 641064 70226 641066
rect 67725 641008 67730 641064
rect 67786 641008 70226 641064
rect 67725 641006 70226 641008
rect 67725 641003 67791 641006
rect 67633 640522 67699 640525
rect 70166 640522 70226 640628
rect 67633 640520 70226 640522
rect 67633 640464 67638 640520
rect 67694 640464 70226 640520
rect 67633 640462 70226 640464
rect 109542 640525 109602 640628
rect 109542 640520 109651 640525
rect 109542 640464 109590 640520
rect 109646 640464 109651 640520
rect 109542 640462 109651 640464
rect 67633 640459 67699 640462
rect 109585 640459 109651 640462
rect 112897 639978 112963 639981
rect 109940 639976 112963 639978
rect 109940 639920 112902 639976
rect 112958 639920 112963 639976
rect 109940 639918 112963 639920
rect 112897 639915 112963 639918
rect 80973 639844 81039 639845
rect 80973 639840 81020 639844
rect 81084 639842 81090 639844
rect 80973 639784 80978 639840
rect 80973 639780 81020 639784
rect 81084 639782 81130 639842
rect 81084 639780 81090 639782
rect 108246 639780 108252 639844
rect 108316 639842 108322 639844
rect 109493 639842 109559 639845
rect 108316 639840 109559 639842
rect 108316 639784 109498 639840
rect 109554 639784 109559 639840
rect 108316 639782 109559 639784
rect 108316 639780 108322 639782
rect 80973 639779 81039 639780
rect 109493 639779 109559 639782
rect 95877 639706 95943 639709
rect 96286 639706 96292 639708
rect 95877 639704 96292 639706
rect 95877 639648 95882 639704
rect 95938 639648 96292 639704
rect 95877 639646 96292 639648
rect 95877 639643 95943 639646
rect 96286 639644 96292 639646
rect 96356 639644 96362 639708
rect 77385 638890 77451 638893
rect 78438 638890 78444 638892
rect 77385 638888 78444 638890
rect 77385 638832 77390 638888
rect 77446 638832 78444 638888
rect 77385 638830 78444 638832
rect 77385 638827 77451 638830
rect 78438 638828 78444 638830
rect 78508 638828 78514 638892
rect 81433 638890 81499 638893
rect 82486 638890 82492 638892
rect 81433 638888 82492 638890
rect 81433 638832 81438 638888
rect 81494 638832 82492 638888
rect 81433 638830 82492 638832
rect 81433 638827 81499 638830
rect 82486 638828 82492 638830
rect 82556 638828 82562 638892
rect 84285 638890 84351 638893
rect 84510 638890 84516 638892
rect 84285 638888 84516 638890
rect 84285 638832 84290 638888
rect 84346 638832 84516 638888
rect 84285 638830 84516 638832
rect 84285 638827 84351 638830
rect 84510 638828 84516 638830
rect 84580 638828 84586 638892
rect 92238 638828 92244 638892
rect 92308 638890 92314 638892
rect 92381 638890 92447 638893
rect 92308 638888 92447 638890
rect 92308 638832 92386 638888
rect 92442 638832 92447 638888
rect 92308 638830 92447 638832
rect 92308 638828 92314 638830
rect 92381 638827 92447 638830
rect 100293 638890 100359 638893
rect 100518 638890 100524 638892
rect 100293 638888 100524 638890
rect 100293 638832 100298 638888
rect 100354 638832 100524 638888
rect 100293 638830 100524 638832
rect 100293 638827 100359 638830
rect 100518 638828 100524 638830
rect 100588 638828 100594 638892
rect 103278 638828 103284 638892
rect 103348 638890 103354 638892
rect 103421 638890 103487 638893
rect 103348 638888 103487 638890
rect 103348 638832 103426 638888
rect 103482 638832 103487 638888
rect 103348 638830 103487 638832
rect 103348 638828 103354 638830
rect 103421 638827 103487 638830
rect 108982 638828 108988 638892
rect 109052 638890 109058 638892
rect 109677 638890 109743 638893
rect 109052 638888 109743 638890
rect 109052 638832 109682 638888
rect 109738 638832 109743 638888
rect 109052 638830 109743 638832
rect 109052 638828 109058 638830
rect 109677 638827 109743 638830
rect 89294 638692 89300 638756
rect 89364 638754 89370 638756
rect 95141 638754 95207 638757
rect 89364 638752 95207 638754
rect 89364 638696 95146 638752
rect 95202 638696 95207 638752
rect 89364 638694 95207 638696
rect 89364 638692 89370 638694
rect 95141 638691 95207 638694
rect 107377 638618 107443 638621
rect 113173 638618 113239 638621
rect 115197 638618 115263 638621
rect 107377 638616 115263 638618
rect 107377 638560 107382 638616
rect 107438 638560 113178 638616
rect 113234 638560 115202 638616
rect 115258 638560 115263 638616
rect 107377 638558 115263 638560
rect 107377 638555 107443 638558
rect 113173 638555 113239 638558
rect 115197 638555 115263 638558
rect 104934 637604 104940 637668
rect 105004 637666 105010 637668
rect 105445 637666 105511 637669
rect 105004 637664 105511 637666
rect 105004 637608 105450 637664
rect 105506 637608 105511 637664
rect 105004 637606 105511 637608
rect 105004 637604 105010 637606
rect 105445 637603 105511 637606
rect 109166 637604 109172 637668
rect 109236 637666 109242 637668
rect 109401 637666 109467 637669
rect 109236 637664 109467 637666
rect 109236 637608 109406 637664
rect 109462 637608 109467 637664
rect 109236 637606 109467 637608
rect 109236 637604 109242 637606
rect 109401 637603 109467 637606
rect -960 632090 480 632180
rect 4061 632090 4127 632093
rect -960 632088 4127 632090
rect -960 632032 4066 632088
rect 4122 632032 4127 632088
rect -960 632030 4127 632032
rect -960 631940 480 632030
rect 4061 632027 4127 632030
rect 579797 630866 579863 630869
rect 583520 630866 584960 630956
rect 579797 630864 584960 630866
rect 579797 630808 579802 630864
rect 579858 630808 584960 630864
rect 579797 630806 584960 630808
rect 579797 630803 579863 630806
rect 583520 630716 584960 630806
rect 55070 629852 55076 629916
rect 55140 629914 55146 629916
rect 85573 629914 85639 629917
rect 55140 629912 85639 629914
rect 55140 629856 85578 629912
rect 85634 629856 85639 629912
rect 55140 629854 85639 629856
rect 55140 629852 55146 629854
rect 85573 629851 85639 629854
rect 86953 629914 87019 629917
rect 121678 629914 121684 629916
rect 86953 629912 121684 629914
rect 86953 629856 86958 629912
rect 87014 629856 121684 629912
rect 86953 629854 121684 629856
rect 86953 629851 87019 629854
rect 121678 629852 121684 629854
rect 121748 629852 121754 629916
rect 89345 627194 89411 627197
rect 122966 627194 122972 627196
rect 89345 627192 122972 627194
rect 89345 627136 89350 627192
rect 89406 627136 122972 627192
rect 89345 627134 122972 627136
rect 89345 627131 89411 627134
rect 122966 627132 122972 627134
rect 123036 627132 123042 627196
rect 50838 624412 50844 624476
rect 50908 624474 50914 624476
rect 77477 624474 77543 624477
rect 50908 624472 77543 624474
rect 50908 624416 77482 624472
rect 77538 624416 77543 624472
rect 50908 624414 77543 624416
rect 50908 624412 50914 624414
rect 77477 624411 77543 624414
rect -960 619170 480 619260
rect 3509 619170 3575 619173
rect -960 619168 3575 619170
rect -960 619112 3514 619168
rect 3570 619112 3575 619168
rect -960 619110 3575 619112
rect -960 619020 480 619110
rect 3509 619107 3575 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3417 606114 3483 606117
rect -960 606112 3483 606114
rect -960 606056 3422 606112
rect 3478 606056 3483 606112
rect -960 606054 3483 606056
rect -960 605964 480 606054
rect 3417 606051 3483 606054
rect 583520 604060 584960 604300
rect 89621 593466 89687 593469
rect 92606 593466 92612 593468
rect 89621 593464 92612 593466
rect 89621 593408 89626 593464
rect 89682 593408 92612 593464
rect 89621 593406 92612 593408
rect 89621 593403 89687 593406
rect 92606 593404 92612 593406
rect 92676 593404 92682 593468
rect 91001 593330 91067 593333
rect 94078 593330 94084 593332
rect 91001 593328 94084 593330
rect 91001 593272 91006 593328
rect 91062 593272 94084 593328
rect 91001 593270 94084 593272
rect 91001 593267 91067 593270
rect 94078 593268 94084 593270
rect 94148 593268 94154 593332
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect 96429 590068 96495 590069
rect 96429 590066 96476 590068
rect 96384 590064 96476 590066
rect 96384 590008 96434 590064
rect 96384 590006 96476 590008
rect 96429 590004 96476 590006
rect 96540 590004 96546 590068
rect 96429 590003 96495 590004
rect 97257 589930 97323 589933
rect 101254 589930 101260 589932
rect 97257 589928 101260 589930
rect 97257 589872 97262 589928
rect 97318 589872 101260 589928
rect 97257 589870 101260 589872
rect 97257 589867 97323 589870
rect 101254 589868 101260 589870
rect 101324 589930 101330 589932
rect 127249 589930 127315 589933
rect 101324 589928 127315 589930
rect 101324 589872 127254 589928
rect 127310 589872 127315 589928
rect 101324 589870 127315 589872
rect 101324 589868 101330 589870
rect 127249 589867 127315 589870
rect 91093 589386 91159 589389
rect 92381 589386 92447 589389
rect 124254 589386 124260 589388
rect 91093 589384 124260 589386
rect 91093 589328 91098 589384
rect 91154 589328 92386 589384
rect 92442 589328 124260 589384
rect 91093 589326 124260 589328
rect 91093 589323 91159 589326
rect 92381 589323 92447 589326
rect 124254 589324 124260 589326
rect 124324 589324 124330 589388
rect 75729 589250 75795 589253
rect 78806 589250 78812 589252
rect 75729 589248 78812 589250
rect 75729 589192 75734 589248
rect 75790 589192 78812 589248
rect 75729 589190 78812 589192
rect 75729 589187 75795 589190
rect 78806 589188 78812 589190
rect 78876 589188 78882 589252
rect 79961 589250 80027 589253
rect 82854 589250 82860 589252
rect 79961 589248 82860 589250
rect 79961 589192 79966 589248
rect 80022 589192 82860 589248
rect 79961 589190 82860 589192
rect 79961 589187 80027 589190
rect 82854 589188 82860 589190
rect 82924 589188 82930 589252
rect 96521 589250 96587 589253
rect 99966 589250 99972 589252
rect 96521 589248 99972 589250
rect 96521 589192 96526 589248
rect 96582 589192 99972 589248
rect 96521 589190 99972 589192
rect 96521 589187 96587 589190
rect 99966 589188 99972 589190
rect 100036 589188 100042 589252
rect 88241 588570 88307 588573
rect 91502 588570 91508 588572
rect 88241 588568 91508 588570
rect 88241 588512 88246 588568
rect 88302 588512 91508 588568
rect 88241 588510 91508 588512
rect 88241 588507 88307 588510
rect 91502 588508 91508 588510
rect 91572 588570 91578 588572
rect 120022 588570 120028 588572
rect 91572 588510 120028 588570
rect 91572 588508 91578 588510
rect 120022 588508 120028 588510
rect 120092 588508 120098 588572
rect 84285 588298 84351 588301
rect 87086 588298 87092 588300
rect 64830 588296 87092 588298
rect 64830 588240 84290 588296
rect 84346 588240 87092 588296
rect 64830 588238 87092 588240
rect 45185 588162 45251 588165
rect 64830 588162 64890 588238
rect 84285 588235 84351 588238
rect 87086 588236 87092 588238
rect 87156 588236 87162 588300
rect 45185 588160 64890 588162
rect 45185 588104 45190 588160
rect 45246 588104 64890 588160
rect 45185 588102 64890 588104
rect 45185 588099 45251 588102
rect 66110 587964 66116 588028
rect 66180 588026 66186 588028
rect 580257 588026 580323 588029
rect 66180 588024 580323 588026
rect 66180 587968 580262 588024
rect 580318 587968 580323 588024
rect 66180 587966 580323 587968
rect 66180 587964 66186 587966
rect 580257 587963 580323 587966
rect 76741 587890 76807 587893
rect 97165 587892 97231 587893
rect 106917 587892 106983 587893
rect 80094 587890 80100 587892
rect 76741 587888 80100 587890
rect 76741 587832 76746 587888
rect 76802 587832 80100 587888
rect 76741 587830 80100 587832
rect 76741 587827 76807 587830
rect 80094 587828 80100 587830
rect 80164 587828 80170 587892
rect 97165 587890 97212 587892
rect 97120 587888 97212 587890
rect 97120 587832 97170 587888
rect 97120 587830 97212 587832
rect 97165 587828 97212 587830
rect 97276 587828 97282 587892
rect 106917 587890 106964 587892
rect 106872 587888 106964 587890
rect 106872 587832 106922 587888
rect 106872 587830 106964 587832
rect 106917 587828 106964 587830
rect 107028 587828 107034 587892
rect 97165 587827 97231 587828
rect 106917 587827 106983 587828
rect 78673 587754 78739 587757
rect 79174 587754 79180 587756
rect 78673 587752 79180 587754
rect 78673 587696 78678 587752
rect 78734 587696 79180 587752
rect 78673 587694 79180 587696
rect 78673 587691 78739 587694
rect 79174 587692 79180 587694
rect 79244 587692 79250 587756
rect 103145 587482 103211 587485
rect 106774 587482 106780 587484
rect 103145 587480 106780 587482
rect 103145 587424 103150 587480
rect 103206 587424 106780 587480
rect 103145 587422 106780 587424
rect 103145 587419 103211 587422
rect 106774 587420 106780 587422
rect 106844 587482 106850 587484
rect 117589 587482 117655 587485
rect 106844 587480 117655 587482
rect 106844 587424 117594 587480
rect 117650 587424 117655 587480
rect 106844 587422 117655 587424
rect 106844 587420 106850 587422
rect 117589 587419 117655 587422
rect 102726 587284 102732 587348
rect 102796 587346 102802 587348
rect 116117 587346 116183 587349
rect 102796 587344 116183 587346
rect 102796 587288 116122 587344
rect 116178 587288 116183 587344
rect 102796 587286 116183 587288
rect 102796 587284 102802 587286
rect 116117 587283 116183 587286
rect 94957 587210 95023 587213
rect 98494 587210 98500 587212
rect 94957 587208 98500 587210
rect 94957 587152 94962 587208
rect 95018 587152 98500 587208
rect 94957 587150 98500 587152
rect 94957 587147 95023 587150
rect 98494 587148 98500 587150
rect 98564 587210 98570 587212
rect 118877 587210 118943 587213
rect 98564 587208 118943 587210
rect 98564 587152 118882 587208
rect 118938 587152 118943 587208
rect 98564 587150 118943 587152
rect 98564 587148 98570 587150
rect 118877 587147 118943 587150
rect 41321 586802 41387 586805
rect 73337 586802 73403 586805
rect 41321 586800 73403 586802
rect 41321 586744 41326 586800
rect 41382 586744 73342 586800
rect 73398 586744 73403 586800
rect 41321 586742 73403 586744
rect 41321 586739 41387 586742
rect 73337 586739 73403 586742
rect 46565 586666 46631 586669
rect 78673 586666 78739 586669
rect 46565 586664 78739 586666
rect 46565 586608 46570 586664
rect 46626 586608 78678 586664
rect 78734 586608 78739 586664
rect 46565 586606 78739 586608
rect 46565 586603 46631 586606
rect 78673 586603 78739 586606
rect 73102 586468 73108 586532
rect 73172 586468 73178 586532
rect 75862 586468 75868 586532
rect 75932 586468 75938 586532
rect 84101 586530 84167 586533
rect 84101 586528 84210 586530
rect 84101 586472 84106 586528
rect 84162 586472 84210 586528
rect 35709 586394 35775 586397
rect 70761 586394 70827 586397
rect 73110 586394 73170 586468
rect 35709 586392 73170 586394
rect 35709 586336 35714 586392
rect 35770 586336 70766 586392
rect 70822 586336 73170 586392
rect 35709 586334 73170 586336
rect 73337 586394 73403 586397
rect 75870 586394 75930 586468
rect 84101 586467 84210 586472
rect 85798 586468 85804 586532
rect 85868 586468 85874 586532
rect 102726 586468 102732 586532
rect 102796 586468 102802 586532
rect 73337 586392 75930 586394
rect 73337 586336 73342 586392
rect 73398 586336 75930 586392
rect 73337 586334 75930 586336
rect 84150 586394 84210 586467
rect 85806 586394 85866 586468
rect 84150 586334 85866 586394
rect 98729 586394 98795 586397
rect 102734 586394 102794 586468
rect 98729 586392 102794 586394
rect 98729 586336 98734 586392
rect 98790 586336 102794 586392
rect 98729 586334 102794 586336
rect 35709 586331 35775 586334
rect 70761 586331 70827 586334
rect 73337 586331 73403 586334
rect 98729 586331 98795 586334
rect 47945 585578 48011 585581
rect 48078 585578 48084 585580
rect 47945 585576 48084 585578
rect 47945 585520 47950 585576
rect 48006 585520 48084 585576
rect 47945 585518 48084 585520
rect 47945 585515 48011 585518
rect 48078 585516 48084 585518
rect 48148 585516 48154 585580
rect 71957 585578 72023 585581
rect 72693 585578 72759 585581
rect 74758 585578 74764 585580
rect 71957 585576 74764 585578
rect 71957 585520 71962 585576
rect 72018 585520 72698 585576
rect 72754 585520 74764 585576
rect 71957 585518 74764 585520
rect 71957 585515 72023 585518
rect 72693 585515 72759 585518
rect 74758 585516 74764 585518
rect 74828 585516 74834 585580
rect 78254 585578 78260 585580
rect 75870 585518 78260 585578
rect 43805 585442 43871 585445
rect 75870 585442 75930 585518
rect 78254 585516 78260 585518
rect 78324 585516 78330 585580
rect 101305 585578 101371 585581
rect 105537 585580 105603 585581
rect 101990 585578 101996 585580
rect 101305 585576 101996 585578
rect 101305 585520 101310 585576
rect 101366 585520 101996 585576
rect 101305 585518 101996 585520
rect 101305 585515 101371 585518
rect 101990 585516 101996 585518
rect 102060 585578 102066 585580
rect 105486 585578 105492 585580
rect 102060 585518 103530 585578
rect 105446 585518 105492 585578
rect 105556 585576 105603 585580
rect 105598 585520 105603 585576
rect 102060 585516 102066 585518
rect 43805 585440 75930 585442
rect 43805 585384 43810 585440
rect 43866 585384 75930 585440
rect 43805 585382 75930 585384
rect 76005 585442 76071 585445
rect 77150 585442 77156 585444
rect 76005 585440 77156 585442
rect 76005 585384 76010 585440
rect 76066 585384 77156 585440
rect 76005 585382 77156 585384
rect 43805 585379 43871 585382
rect 76005 585379 76071 585382
rect 77150 585380 77156 585382
rect 77220 585380 77226 585444
rect 84694 585380 84700 585444
rect 84764 585442 84770 585444
rect 85389 585442 85455 585445
rect 84764 585440 85455 585442
rect 84764 585384 85394 585440
rect 85450 585384 85455 585440
rect 84764 585382 85455 585384
rect 103470 585442 103530 585518
rect 105486 585516 105492 585518
rect 105556 585516 105603 585520
rect 105537 585515 105603 585516
rect 130101 585442 130167 585445
rect 103470 585440 130167 585442
rect 103470 585384 130106 585440
rect 130162 585384 130167 585440
rect 103470 585382 130167 585384
rect 84764 585380 84770 585382
rect 85389 585379 85455 585382
rect 130101 585379 130167 585382
rect 54845 585306 54911 585309
rect 120257 585306 120323 585309
rect 54845 585304 87522 585306
rect 54845 585248 54850 585304
rect 54906 585248 87522 585304
rect 54845 585246 87522 585248
rect 54845 585243 54911 585246
rect 70393 585170 70459 585173
rect 78213 585172 78279 585173
rect 71814 585170 71820 585172
rect 70393 585168 71820 585170
rect 70393 585112 70398 585168
rect 70454 585112 71820 585168
rect 70393 585110 71820 585112
rect 70393 585107 70459 585110
rect 71814 585108 71820 585110
rect 71884 585108 71890 585172
rect 78213 585168 78260 585172
rect 78324 585170 78330 585172
rect 85113 585170 85179 585173
rect 87270 585170 87276 585172
rect 78213 585112 78218 585168
rect 78213 585108 78260 585112
rect 78324 585110 78370 585170
rect 85113 585168 87276 585170
rect 85113 585112 85118 585168
rect 85174 585112 87276 585168
rect 85113 585110 87276 585112
rect 78324 585108 78330 585110
rect 78213 585107 78279 585108
rect 85113 585107 85179 585110
rect 87270 585108 87276 585110
rect 87340 585108 87346 585172
rect 87462 585170 87522 585246
rect 93810 585304 120323 585306
rect 93810 585248 120262 585304
rect 120318 585248 120323 585304
rect 93810 585246 120323 585248
rect 88885 585172 88951 585173
rect 88885 585170 88932 585172
rect 87462 585168 88932 585170
rect 88996 585170 89002 585172
rect 90265 585170 90331 585173
rect 90950 585170 90956 585172
rect 87462 585112 88890 585168
rect 87462 585110 88932 585112
rect 88885 585108 88932 585110
rect 88996 585110 89042 585170
rect 90265 585168 90956 585170
rect 90265 585112 90270 585168
rect 90326 585112 90956 585168
rect 90265 585110 90956 585112
rect 88996 585108 89002 585110
rect 88885 585107 88951 585108
rect 90265 585107 90331 585110
rect 90950 585108 90956 585110
rect 91020 585170 91026 585172
rect 93810 585170 93870 585246
rect 120257 585243 120323 585246
rect 91020 585110 93870 585170
rect 97073 585170 97139 585173
rect 97758 585170 97764 585172
rect 97073 585168 97764 585170
rect 97073 585112 97078 585168
rect 97134 585112 97764 585168
rect 97073 585110 97764 585112
rect 91020 585108 91026 585110
rect 97073 585107 97139 585110
rect 97758 585108 97764 585110
rect 97828 585170 97834 585172
rect 131205 585170 131271 585173
rect 97828 585168 131271 585170
rect 97828 585112 131210 585168
rect 131266 585112 131271 585168
rect 97828 585110 131271 585112
rect 97828 585108 97834 585110
rect 131205 585107 131271 585110
rect 60549 584082 60615 584085
rect 70945 584084 71011 584085
rect 70894 584082 70900 584084
rect 60549 584080 70900 584082
rect 70964 584080 71011 584084
rect 60549 584024 60554 584080
rect 60610 584024 70900 584080
rect 71006 584024 71011 584080
rect 60549 584022 70900 584024
rect 60549 584019 60615 584022
rect 70894 584020 70900 584022
rect 70964 584020 71011 584024
rect 70945 584019 71011 584020
rect 72233 584082 72299 584085
rect 99097 584084 99163 584085
rect 72918 584082 72924 584084
rect 72233 584080 72924 584082
rect 72233 584024 72238 584080
rect 72294 584024 72924 584080
rect 72233 584022 72924 584024
rect 72233 584019 72299 584022
rect 72918 584020 72924 584022
rect 72988 584020 72994 584084
rect 99046 584020 99052 584084
rect 99116 584082 99163 584084
rect 104617 584082 104683 584085
rect 104750 584082 104756 584084
rect 99116 584080 99208 584082
rect 99158 584024 99208 584080
rect 99116 584022 99208 584024
rect 104617 584080 104756 584082
rect 104617 584024 104622 584080
rect 104678 584024 104756 584080
rect 104617 584022 104756 584024
rect 99116 584020 99163 584022
rect 99097 584019 99163 584020
rect 104617 584019 104683 584022
rect 104750 584020 104756 584022
rect 104820 584082 104826 584084
rect 104820 584022 113190 584082
rect 104820 584020 104826 584022
rect 52177 583946 52243 583949
rect 74625 583946 74691 583949
rect 75126 583946 75132 583948
rect 52177 583944 75132 583946
rect 52177 583888 52182 583944
rect 52238 583888 74630 583944
rect 74686 583888 75132 583944
rect 52177 583886 75132 583888
rect 52177 583883 52243 583886
rect 74625 583883 74691 583886
rect 75126 583884 75132 583886
rect 75196 583884 75202 583948
rect 104433 583946 104499 583949
rect 104566 583946 104572 583948
rect 104433 583944 104572 583946
rect 104433 583888 104438 583944
rect 104494 583888 104572 583944
rect 104433 583886 104572 583888
rect 104433 583883 104499 583886
rect 104566 583884 104572 583886
rect 104636 583884 104642 583948
rect 113130 583946 113190 584022
rect 116209 583946 116275 583949
rect 113130 583944 116275 583946
rect 113130 583888 116214 583944
rect 116270 583888 116275 583944
rect 113130 583886 116275 583888
rect 116209 583883 116275 583886
rect 53557 583812 53623 583813
rect 51758 583748 51764 583812
rect 51828 583810 51834 583812
rect 51828 583750 53482 583810
rect 51828 583748 51834 583750
rect 53422 583674 53482 583750
rect 53557 583808 53604 583812
rect 53668 583810 53674 583812
rect 75269 583810 75335 583813
rect 75637 583810 75703 583813
rect 84009 583812 84075 583813
rect 53557 583752 53562 583808
rect 53557 583748 53604 583752
rect 53668 583750 53714 583810
rect 53790 583808 75703 583810
rect 53790 583752 75274 583808
rect 75330 583752 75642 583808
rect 75698 583752 75703 583808
rect 53790 583750 75703 583752
rect 53668 583748 53674 583750
rect 53557 583747 53623 583748
rect 53790 583674 53850 583750
rect 75269 583747 75335 583750
rect 75637 583747 75703 583750
rect 83958 583748 83964 583812
rect 84028 583810 84075 583812
rect 86217 583810 86283 583813
rect 93761 583812 93827 583813
rect 86718 583810 86724 583812
rect 84028 583808 84120 583810
rect 84070 583752 84120 583808
rect 84028 583750 84120 583752
rect 86217 583808 86724 583810
rect 86217 583752 86222 583808
rect 86278 583752 86724 583808
rect 86217 583750 86724 583752
rect 84028 583748 84075 583750
rect 84009 583747 84075 583748
rect 86217 583747 86283 583750
rect 86718 583748 86724 583750
rect 86788 583748 86794 583812
rect 93710 583810 93716 583812
rect 93670 583750 93716 583810
rect 93780 583808 93827 583812
rect 93822 583752 93827 583808
rect 93710 583748 93716 583750
rect 93780 583748 93827 583752
rect 93761 583747 93827 583748
rect 99097 583810 99163 583813
rect 127065 583810 127131 583813
rect 99097 583808 127131 583810
rect 99097 583752 99102 583808
rect 99158 583752 127070 583808
rect 127126 583752 127131 583808
rect 99097 583750 127131 583752
rect 99097 583747 99163 583750
rect 127065 583747 127131 583750
rect 53422 583614 53850 583674
rect 107561 582724 107627 582725
rect 107510 582660 107516 582724
rect 107580 582722 107627 582724
rect 107580 582720 107672 582722
rect 107622 582664 107672 582720
rect 107580 582662 107672 582664
rect 107580 582660 107627 582662
rect 107561 582659 107627 582660
rect 94129 582586 94195 582589
rect 94998 582586 95004 582588
rect 94129 582584 95004 582586
rect 94129 582528 94134 582584
rect 94190 582528 95004 582584
rect 94129 582526 95004 582528
rect 94129 582523 94195 582526
rect 94998 582524 95004 582526
rect 95068 582586 95074 582588
rect 128670 582586 128676 582588
rect 95068 582526 128676 582586
rect 95068 582524 95074 582526
rect 128670 582524 128676 582526
rect 128740 582524 128746 582588
rect 83273 582450 83339 582453
rect 84009 582450 84075 582453
rect 117998 582450 118004 582452
rect 83273 582448 118004 582450
rect 83273 582392 83278 582448
rect 83334 582392 84014 582448
rect 84070 582392 118004 582448
rect 83273 582390 118004 582392
rect 83273 582387 83339 582390
rect 84009 582387 84075 582390
rect 117998 582388 118004 582390
rect 118068 582388 118074 582452
rect 58934 581980 58940 582044
rect 59004 582042 59010 582044
rect 81893 582042 81959 582045
rect 82670 582042 82676 582044
rect 59004 582040 82676 582042
rect 59004 581984 81898 582040
rect 81954 581984 82676 582040
rect 59004 581982 82676 581984
rect 59004 581980 59010 581982
rect 81893 581979 81959 581982
rect 82670 581980 82676 581982
rect 82740 581980 82746 582044
rect 100569 581906 100635 581909
rect 125726 581906 125732 581908
rect 100569 581904 125732 581906
rect 100569 581848 100574 581904
rect 100630 581848 125732 581904
rect 100569 581846 125732 581848
rect 100569 581843 100635 581846
rect 125726 581844 125732 581846
rect 125796 581844 125802 581908
rect 121729 581634 121795 581637
rect 122046 581634 122052 581636
rect 121729 581632 122052 581634
rect 121729 581576 121734 581632
rect 121790 581576 122052 581632
rect 121729 581574 122052 581576
rect 121729 581571 121795 581574
rect 122046 581572 122052 581574
rect 122116 581572 122122 581636
rect 70350 581229 70410 581468
rect 70209 581228 70275 581229
rect 70158 581226 70164 581228
rect 70118 581166 70164 581226
rect 70228 581224 70275 581228
rect 70270 581168 70275 581224
rect 70158 581164 70164 581166
rect 70228 581164 70275 581168
rect 70350 581224 70459 581229
rect 70350 581168 70398 581224
rect 70454 581168 70459 581224
rect 70350 581166 70459 581168
rect 70209 581163 70275 581164
rect 70393 581163 70459 581166
rect 108941 580954 109007 580957
rect 105892 580952 109007 580954
rect 105892 580896 108946 580952
rect 109002 580896 109007 580952
rect 105892 580894 109007 580896
rect 108941 580891 109007 580894
rect 69289 580682 69355 580685
rect 69657 580682 69723 580685
rect 70166 580682 70226 580788
rect 69289 580680 70226 580682
rect 69289 580624 69294 580680
rect 69350 580624 69662 580680
rect 69718 580624 70226 580680
rect 69289 580622 70226 580624
rect 69289 580619 69355 580622
rect 69657 580619 69723 580622
rect 108021 580274 108087 580277
rect 105892 580272 108087 580274
rect 105892 580216 108026 580272
rect 108082 580216 108087 580272
rect 105892 580214 108087 580216
rect 108021 580211 108087 580214
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 118693 579730 118759 579733
rect 122598 579730 122604 579732
rect 118693 579728 122604 579730
rect 118693 579672 118698 579728
rect 118754 579672 122604 579728
rect 118693 579670 122604 579672
rect 118693 579667 118759 579670
rect 122598 579668 122604 579670
rect 122668 579668 122674 579732
rect 108941 579594 109007 579597
rect 105892 579592 109007 579594
rect 105892 579536 108946 579592
rect 109002 579536 109007 579592
rect 105892 579534 109007 579536
rect 108941 579531 109007 579534
rect 67633 579322 67699 579325
rect 70350 579324 70410 579428
rect 67633 579320 70226 579322
rect 67633 579264 67638 579320
rect 67694 579264 70226 579320
rect 67633 579262 70226 579264
rect 67633 579259 67699 579262
rect 70166 578884 70226 579262
rect 70342 579260 70348 579324
rect 70412 579260 70418 579324
rect 107510 578778 107516 578780
rect 105892 578718 107516 578778
rect 107510 578716 107516 578718
rect 107580 578778 107586 578780
rect 108665 578778 108731 578781
rect 107580 578776 108731 578778
rect 107580 578720 108670 578776
rect 108726 578720 108731 578776
rect 107580 578718 108731 578720
rect 107580 578716 107586 578718
rect 108665 578715 108731 578718
rect 64638 578444 64644 578508
rect 64708 578506 64714 578508
rect 70342 578506 70348 578508
rect 64708 578446 70348 578506
rect 64708 578444 64714 578446
rect 70342 578444 70348 578446
rect 70412 578444 70418 578508
rect 62982 578172 62988 578236
rect 63052 578234 63058 578236
rect 64689 578234 64755 578237
rect 67725 578234 67791 578237
rect 106089 578234 106155 578237
rect 108113 578234 108179 578237
rect 63052 578232 67791 578234
rect 63052 578176 64694 578232
rect 64750 578176 67730 578232
rect 67786 578176 67791 578232
rect 63052 578174 67791 578176
rect 105892 578232 108179 578234
rect 105892 578176 106094 578232
rect 106150 578176 108118 578232
rect 108174 578176 108179 578232
rect 105892 578174 108179 578176
rect 63052 578172 63058 578174
rect 64689 578171 64755 578174
rect 67725 578171 67791 578174
rect 106089 578171 106155 578174
rect 108113 578171 108179 578174
rect 116393 578234 116459 578237
rect 117078 578234 117084 578236
rect 116393 578232 117084 578234
rect 116393 578176 116398 578232
rect 116454 578176 117084 578232
rect 116393 578174 117084 578176
rect 116393 578171 116459 578174
rect 117078 578172 117084 578174
rect 117148 578234 117154 578236
rect 118734 578234 118740 578236
rect 117148 578174 118740 578234
rect 117148 578172 117154 578174
rect 118734 578172 118740 578174
rect 118804 578172 118810 578236
rect 67633 577826 67699 577829
rect 70350 577826 70410 578068
rect 67633 577824 70410 577826
rect 67633 577768 67638 577824
rect 67694 577768 70410 577824
rect 67633 577766 70410 577768
rect 67633 577763 67699 577766
rect 107009 577690 107075 577693
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 107009 577688 113190 577690
rect 107009 577632 107014 577688
rect 107070 577632 113190 577688
rect 107009 577630 113190 577632
rect 107009 577627 107075 577630
rect 108941 577554 109007 577557
rect 105892 577552 109007 577554
rect 105892 577496 108946 577552
rect 109002 577496 109007 577552
rect 105892 577494 109007 577496
rect 113130 577554 113190 577630
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 118734 577554 118740 577556
rect 113130 577494 118740 577554
rect 108941 577491 109007 577494
rect 118734 577492 118740 577494
rect 118804 577492 118810 577556
rect 583520 577540 584960 577630
rect 67725 577282 67791 577285
rect 70166 577282 70226 577388
rect 67725 577280 70226 577282
rect 67725 577224 67730 577280
rect 67786 577224 70226 577280
rect 67725 577222 70226 577224
rect 67725 577219 67791 577222
rect 108757 576738 108823 576741
rect 105892 576736 108823 576738
rect 68645 576602 68711 576605
rect 70166 576602 70226 576708
rect 105892 576680 108762 576736
rect 108818 576680 108823 576736
rect 105892 576678 108823 576680
rect 108757 576675 108823 576678
rect 68645 576600 70226 576602
rect 68645 576544 68650 576600
rect 68706 576544 70226 576600
rect 68645 576542 70226 576544
rect 68645 576539 68711 576542
rect 107510 576194 107516 576196
rect 105892 576134 107516 576194
rect 107510 576132 107516 576134
rect 107580 576194 107586 576196
rect 108665 576194 108731 576197
rect 107580 576192 108731 576194
rect 107580 576136 108670 576192
rect 108726 576136 108731 576192
rect 107580 576134 108731 576136
rect 107580 576132 107586 576134
rect 108665 576131 108731 576134
rect 115974 576132 115980 576196
rect 116044 576194 116050 576196
rect 116301 576194 116367 576197
rect 117129 576194 117195 576197
rect 116044 576192 117195 576194
rect 116044 576136 116306 576192
rect 116362 576136 117134 576192
rect 117190 576136 117195 576192
rect 116044 576134 117195 576136
rect 116044 576132 116050 576134
rect 116301 576131 116367 576134
rect 117129 576131 117195 576134
rect 67633 575786 67699 575789
rect 70166 575786 70226 576028
rect 67633 575784 70226 575786
rect 67633 575728 67638 575784
rect 67694 575728 70226 575784
rect 67633 575726 70226 575728
rect 67633 575723 67699 575726
rect 61694 575316 61700 575380
rect 61764 575378 61770 575380
rect 61764 575318 64890 575378
rect 61764 575316 61770 575318
rect 64830 575242 64890 575318
rect 67449 575242 67515 575245
rect 70166 575242 70226 575348
rect 64830 575240 70226 575242
rect 64830 575184 67454 575240
rect 67510 575184 70226 575240
rect 64830 575182 70226 575184
rect 67449 575179 67515 575182
rect 106917 575106 106983 575109
rect 114502 575106 114508 575108
rect 106917 575104 114508 575106
rect 106917 575048 106922 575104
rect 106978 575048 114508 575104
rect 106917 575046 114508 575048
rect 106917 575043 106983 575046
rect 114502 575044 114508 575046
rect 114572 575044 114578 575108
rect 107101 574698 107167 574701
rect 115974 574698 115980 574700
rect 107101 574696 115980 574698
rect 67633 574562 67699 574565
rect 70166 574562 70226 574668
rect 67633 574560 70226 574562
rect 67633 574504 67638 574560
rect 67694 574504 70226 574560
rect 67633 574502 70226 574504
rect 67633 574499 67699 574502
rect 105678 574429 105738 574668
rect 107101 574640 107106 574696
rect 107162 574640 115980 574696
rect 107101 574638 115980 574640
rect 107101 574635 107167 574638
rect 115974 574636 115980 574638
rect 116044 574636 116050 574700
rect 105629 574424 105738 574429
rect 105629 574368 105634 574424
rect 105690 574368 105738 574424
rect 105629 574366 105738 574368
rect 105629 574363 105695 574366
rect 60590 573956 60596 574020
rect 60660 574018 60666 574020
rect 66069 574018 66135 574021
rect 67725 574018 67791 574021
rect 108941 574018 109007 574021
rect 60660 574016 67791 574018
rect 60660 573960 66074 574016
rect 66130 573960 67730 574016
rect 67786 573960 67791 574016
rect 105892 574016 109007 574018
rect 60660 573958 67791 573960
rect 60660 573956 60666 573958
rect 66069 573955 66135 573958
rect 67725 573955 67791 573958
rect 67633 573882 67699 573885
rect 70166 573882 70226 573988
rect 105892 573960 108946 574016
rect 109002 573960 109007 574016
rect 105892 573958 109007 573960
rect 108941 573955 109007 573958
rect 67633 573880 70226 573882
rect 67633 573824 67638 573880
rect 67694 573824 70226 573880
rect 67633 573822 70226 573824
rect 67633 573819 67699 573822
rect 67725 573338 67791 573341
rect 108941 573338 109007 573341
rect 67725 573336 70226 573338
rect 67725 573280 67730 573336
rect 67786 573280 70226 573336
rect 67725 573278 70226 573280
rect 105892 573336 109007 573338
rect 105892 573280 108946 573336
rect 109002 573280 109007 573336
rect 105892 573278 109007 573280
rect 67725 573275 67791 573278
rect 70166 572764 70226 573278
rect 108941 573275 109007 573278
rect 107377 572794 107443 572797
rect 108573 572794 108639 572797
rect 122925 572796 122991 572797
rect 122925 572794 122972 572796
rect 105892 572792 108639 572794
rect 105892 572736 107382 572792
rect 107438 572736 108578 572792
rect 108634 572736 108639 572792
rect 105892 572734 108639 572736
rect 122880 572792 122972 572794
rect 122880 572736 122930 572792
rect 122880 572734 122972 572736
rect 107377 572731 107443 572734
rect 108573 572731 108639 572734
rect 122925 572732 122972 572734
rect 123036 572732 123042 572796
rect 122925 572731 122991 572732
rect 66662 572324 66668 572388
rect 66732 572386 66738 572388
rect 66732 572326 70410 572386
rect 66732 572324 66738 572326
rect 70350 572084 70410 572326
rect 108297 571978 108363 571981
rect 105892 571976 108363 571978
rect 105892 571920 108302 571976
rect 108358 571920 108363 571976
rect 105892 571918 108363 571920
rect 108297 571915 108363 571918
rect 67633 571706 67699 571709
rect 67633 571704 70226 571706
rect 67633 571648 67638 571704
rect 67694 571648 70226 571704
rect 67633 571646 70226 571648
rect 67633 571643 67699 571646
rect 70166 571404 70226 571646
rect 108021 571434 108087 571437
rect 105892 571432 108087 571434
rect 105892 571376 108026 571432
rect 108082 571376 108087 571432
rect 105892 571374 108087 571376
rect 108021 571371 108087 571374
rect 66110 570964 66116 571028
rect 66180 571026 66186 571028
rect 67633 571026 67699 571029
rect 66180 571024 70410 571026
rect 66180 570968 67638 571024
rect 67694 570968 70410 571024
rect 66180 570966 70410 570968
rect 66180 570964 66186 570966
rect 67633 570963 67699 570966
rect 70350 570724 70410 570966
rect 108798 570754 108804 570756
rect 105892 570694 108804 570754
rect 108798 570692 108804 570694
rect 108868 570754 108874 570756
rect 136909 570754 136975 570757
rect 108868 570752 136975 570754
rect 108868 570696 136914 570752
rect 136970 570696 136975 570752
rect 108868 570694 136975 570696
rect 108868 570692 108874 570694
rect 136909 570691 136975 570694
rect 139485 570618 139551 570621
rect 113130 570616 139551 570618
rect 113130 570560 139490 570616
rect 139546 570560 139551 570616
rect 113130 570558 139551 570560
rect 108246 570482 108252 570484
rect 105862 570422 108252 570482
rect 67725 570346 67791 570349
rect 67725 570344 70226 570346
rect 67725 570288 67730 570344
rect 67786 570288 70226 570344
rect 67725 570286 70226 570288
rect 67725 570283 67791 570286
rect 70166 570044 70226 570286
rect 105862 570044 105922 570422
rect 108246 570420 108252 570422
rect 108316 570482 108322 570484
rect 113130 570482 113190 570558
rect 139485 570555 139551 570558
rect 108316 570422 113190 570482
rect 108316 570420 108322 570422
rect 108941 569258 109007 569261
rect 105892 569256 109007 569258
rect 67633 569122 67699 569125
rect 70166 569122 70226 569228
rect 105892 569200 108946 569256
rect 109002 569200 109007 569256
rect 105892 569198 109007 569200
rect 108941 569195 109007 569198
rect 67633 569120 70226 569122
rect 67633 569064 67638 569120
rect 67694 569064 70226 569120
rect 67633 569062 70226 569064
rect 67633 569059 67699 569062
rect 67817 568986 67883 568989
rect 67817 568984 70410 568986
rect 67817 568928 67822 568984
rect 67878 568928 70410 568984
rect 67817 568926 70410 568928
rect 67817 568923 67883 568926
rect 70350 568684 70410 568926
rect 43713 568578 43779 568581
rect 44030 568578 44036 568580
rect 43713 568576 44036 568578
rect 43713 568520 43718 568576
rect 43774 568520 44036 568576
rect 43713 568518 44036 568520
rect 43713 568515 43779 568518
rect 44030 568516 44036 568518
rect 44100 568516 44106 568580
rect 113214 568516 113220 568580
rect 113284 568578 113290 568580
rect 113449 568578 113515 568581
rect 113284 568576 113515 568578
rect 113284 568520 113454 568576
rect 113510 568520 113515 568576
rect 113284 568518 113515 568520
rect 113284 568516 113290 568518
rect 113449 568515 113515 568518
rect 67633 568306 67699 568309
rect 67633 568304 70410 568306
rect 67633 568248 67638 568304
rect 67694 568248 70410 568304
rect 67633 568246 70410 568248
rect 67633 568243 67699 568246
rect 70350 568004 70410 568246
rect 108941 567898 109007 567901
rect 105892 567896 109007 567898
rect 105892 567840 108946 567896
rect 109002 567840 109007 567896
rect 105892 567838 109007 567840
rect 108941 567835 109007 567838
rect 67633 567762 67699 567765
rect 67633 567760 70226 567762
rect 67633 567704 67638 567760
rect 67694 567704 70226 567760
rect 67633 567702 70226 567704
rect 67633 567699 67699 567702
rect 70166 567324 70226 567702
rect 108849 567354 108915 567357
rect 105892 567352 108915 567354
rect 105892 567296 108854 567352
rect 108910 567296 108915 567352
rect 105892 567294 108915 567296
rect 108849 567291 108915 567294
rect -960 566946 480 567036
rect 3233 566946 3299 566949
rect -960 566944 3299 566946
rect -960 566888 3238 566944
rect 3294 566888 3299 566944
rect -960 566886 3299 566888
rect -960 566796 480 566886
rect 3233 566883 3299 566886
rect 108941 566538 109007 566541
rect 105892 566536 109007 566538
rect 105892 566480 108946 566536
rect 109002 566480 109007 566536
rect 105892 566478 109007 566480
rect 108941 566475 109007 566478
rect 67633 566402 67699 566405
rect 67633 566400 70226 566402
rect 67633 566344 67638 566400
rect 67694 566344 70226 566400
rect 67633 566342 70226 566344
rect 67633 566339 67699 566342
rect 70166 565964 70226 566342
rect 108941 565858 109007 565861
rect 105892 565856 109007 565858
rect 105892 565800 108946 565856
rect 109002 565800 109007 565856
rect 105892 565798 109007 565800
rect 108941 565795 109007 565798
rect 108849 565314 108915 565317
rect 105892 565312 108915 565314
rect 105892 565256 108854 565312
rect 108910 565256 108915 565312
rect 105892 565254 108915 565256
rect 108849 565251 108915 565254
rect 67633 565042 67699 565045
rect 70166 565042 70226 565148
rect 111190 565042 111196 565044
rect 67633 565040 70226 565042
rect 67633 564984 67638 565040
rect 67694 564984 70226 565040
rect 67633 564982 70226 564984
rect 105862 564982 111196 565042
rect 67633 564979 67699 564982
rect 67633 564906 67699 564909
rect 67633 564904 70410 564906
rect 67633 564848 67638 564904
rect 67694 564848 70410 564904
rect 67633 564846 70410 564848
rect 67633 564843 67699 564846
rect 70350 564604 70410 564846
rect 105862 564604 105922 564982
rect 111190 564980 111196 564982
rect 111260 565042 111266 565044
rect 138105 565042 138171 565045
rect 111260 565040 138171 565042
rect 111260 564984 138110 565040
rect 138166 564984 138171 565040
rect 111260 564982 138171 564984
rect 111260 564980 111266 564982
rect 138105 564979 138171 564982
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 67633 564226 67699 564229
rect 67633 564224 70226 564226
rect 67633 564168 67638 564224
rect 67694 564168 70226 564224
rect 583520 564212 584960 564302
rect 67633 564166 70226 564168
rect 67633 564163 67699 564166
rect 70166 563924 70226 564166
rect 108941 563818 109007 563821
rect 105892 563816 109007 563818
rect 105892 563760 108946 563816
rect 109002 563760 109007 563816
rect 105892 563758 109007 563760
rect 108941 563755 109007 563758
rect 67725 563682 67791 563685
rect 67725 563680 70226 563682
rect 67725 563624 67730 563680
rect 67786 563624 70226 563680
rect 67725 563622 70226 563624
rect 67725 563619 67791 563622
rect 70166 563244 70226 563622
rect 108941 563138 109007 563141
rect 105892 563136 109007 563138
rect 105892 563080 108946 563136
rect 109002 563080 109007 563136
rect 105892 563078 109007 563080
rect 108941 563075 109007 563078
rect 108849 562458 108915 562461
rect 105892 562456 108915 562458
rect 67633 562322 67699 562325
rect 70166 562322 70226 562428
rect 105892 562400 108854 562456
rect 108910 562400 108915 562456
rect 105892 562398 108915 562400
rect 108849 562395 108915 562398
rect 67633 562320 70226 562322
rect 67633 562264 67638 562320
rect 67694 562264 70226 562320
rect 67633 562262 70226 562264
rect 67633 562259 67699 562262
rect 64830 562126 70410 562186
rect 58750 561852 58756 561916
rect 58820 561914 58826 561916
rect 61878 561914 61884 561916
rect 58820 561854 61884 561914
rect 58820 561852 58826 561854
rect 61878 561852 61884 561854
rect 61948 561914 61954 561916
rect 64830 561914 64890 562126
rect 61948 561854 64890 561914
rect 70350 561884 70410 562126
rect 61948 561852 61954 561854
rect 67633 561506 67699 561509
rect 67633 561504 70226 561506
rect 67633 561448 67638 561504
rect 67694 561448 70226 561504
rect 67633 561446 70226 561448
rect 67633 561443 67699 561446
rect 70166 561204 70226 561446
rect 108941 561098 109007 561101
rect 105892 561096 109007 561098
rect 105892 561040 108946 561096
rect 109002 561040 109007 561096
rect 105892 561038 109007 561040
rect 108941 561035 109007 561038
rect 67725 560962 67791 560965
rect 67725 560960 70226 560962
rect 67725 560904 67730 560960
rect 67786 560904 70226 560960
rect 67725 560902 70226 560904
rect 67725 560899 67791 560902
rect 70166 560524 70226 560902
rect 107469 560554 107535 560557
rect 108941 560554 109007 560557
rect 105892 560552 109007 560554
rect 105892 560496 107474 560552
rect 107530 560496 108946 560552
rect 109002 560496 109007 560552
rect 105892 560494 109007 560496
rect 107469 560491 107535 560494
rect 108941 560491 109007 560494
rect 108941 559738 109007 559741
rect 105892 559736 109007 559738
rect 105892 559680 108946 559736
rect 109002 559680 109007 559736
rect 105892 559678 109007 559680
rect 108941 559675 109007 559678
rect 67633 559602 67699 559605
rect 67633 559600 70226 559602
rect 67633 559544 67638 559600
rect 67694 559544 70226 559600
rect 67633 559542 70226 559544
rect 67633 559539 67699 559542
rect 70166 559164 70226 559542
rect 108021 559058 108087 559061
rect 105892 559056 108087 559058
rect 105892 559000 108026 559056
rect 108082 559000 108087 559056
rect 105892 558998 108087 559000
rect 108021 558995 108087 558998
rect 107878 558452 107884 558516
rect 107948 558514 107954 558516
rect 108021 558514 108087 558517
rect 107948 558512 108087 558514
rect 107948 558456 108026 558512
rect 108082 558456 108087 558512
rect 107948 558454 108087 558456
rect 107948 558452 107954 558454
rect 108021 558451 108087 558454
rect 108941 558378 109007 558381
rect 105892 558376 109007 558378
rect 67725 558106 67791 558109
rect 70166 558106 70226 558348
rect 105892 558320 108946 558376
rect 109002 558320 109007 558376
rect 105892 558318 109007 558320
rect 108941 558315 109007 558318
rect 111558 558180 111564 558244
rect 111628 558242 111634 558244
rect 121678 558242 121684 558244
rect 111628 558182 121684 558242
rect 111628 558180 111634 558182
rect 121678 558180 121684 558182
rect 121748 558180 121754 558244
rect 67725 558104 70226 558106
rect 67725 558048 67730 558104
rect 67786 558048 70226 558104
rect 67725 558046 70226 558048
rect 67725 558043 67791 558046
rect 107745 557834 107811 557837
rect 105892 557832 107811 557834
rect 105892 557776 107750 557832
rect 107806 557776 107811 557832
rect 105892 557774 107811 557776
rect 107745 557771 107811 557774
rect 67633 557562 67699 557565
rect 70166 557562 70226 557668
rect 67633 557560 70226 557562
rect 67633 557504 67638 557560
rect 67694 557504 70226 557560
rect 67633 557502 70226 557504
rect 67633 557499 67699 557502
rect 67817 557426 67883 557429
rect 67817 557424 70226 557426
rect 67817 557368 67822 557424
rect 67878 557368 70226 557424
rect 67817 557366 70226 557368
rect 67817 557363 67883 557366
rect 70166 557124 70226 557366
rect 108941 557154 109007 557157
rect 105892 557152 109007 557154
rect 105892 557096 108946 557152
rect 109002 557096 109007 557152
rect 105892 557094 109007 557096
rect 108941 557091 109007 557094
rect 67633 556882 67699 556885
rect 67633 556880 70226 556882
rect 67633 556824 67638 556880
rect 67694 556824 70226 556880
rect 67633 556822 70226 556824
rect 67633 556819 67699 556822
rect 70166 556444 70226 556822
rect 105486 556684 105492 556748
rect 105556 556746 105562 556748
rect 108297 556746 108363 556749
rect 105556 556744 108363 556746
rect 105556 556688 108302 556744
rect 108358 556688 108363 556744
rect 105556 556686 108363 556688
rect 105556 556684 105562 556686
rect 108297 556683 108363 556686
rect 107694 556474 107700 556476
rect 105892 556414 107700 556474
rect 107694 556412 107700 556414
rect 107764 556474 107770 556476
rect 111926 556474 111932 556476
rect 107764 556414 111932 556474
rect 107764 556412 107770 556414
rect 111926 556412 111932 556414
rect 111996 556412 112002 556476
rect 108849 555658 108915 555661
rect 105892 555656 108915 555658
rect 67633 555386 67699 555389
rect 70166 555386 70226 555628
rect 105892 555600 108854 555656
rect 108910 555600 108915 555656
rect 105892 555598 108915 555600
rect 108849 555595 108915 555598
rect 67633 555384 70226 555386
rect 67633 555328 67638 555384
rect 67694 555328 70226 555384
rect 67633 555326 70226 555328
rect 67633 555323 67699 555326
rect 67725 554842 67791 554845
rect 70166 554842 70226 554948
rect 67725 554840 70226 554842
rect 67725 554784 67730 554840
rect 67786 554784 70226 554840
rect 67725 554782 70226 554784
rect 67725 554779 67791 554782
rect 67909 554706 67975 554709
rect 68686 554706 68692 554708
rect 67909 554704 68692 554706
rect 67909 554648 67914 554704
rect 67970 554648 68692 554704
rect 67909 554646 68692 554648
rect 67909 554643 67975 554646
rect 68686 554644 68692 554646
rect 68756 554706 68762 554708
rect 68756 554646 70410 554706
rect 68756 554644 68762 554646
rect 70350 554404 70410 554646
rect 108941 554434 109007 554437
rect 105892 554432 109007 554434
rect 105892 554376 108946 554432
rect 109002 554376 109007 554432
rect 105892 554374 109007 554376
rect 108941 554371 109007 554374
rect 67633 554162 67699 554165
rect 67633 554160 70226 554162
rect 67633 554104 67638 554160
rect 67694 554104 70226 554160
rect 67633 554102 70226 554104
rect 67633 554099 67699 554102
rect -960 553890 480 553980
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 70166 553724 70226 554102
rect 108941 553754 109007 553757
rect 105892 553752 109007 553754
rect 105892 553696 108946 553752
rect 109002 553696 109007 553752
rect 105892 553694 109007 553696
rect 108941 553691 109007 553694
rect 56542 553420 56548 553484
rect 56612 553482 56618 553484
rect 57605 553482 57671 553485
rect 56612 553480 57671 553482
rect 56612 553424 57610 553480
rect 57666 553424 57671 553480
rect 56612 553422 57671 553424
rect 56612 553420 56618 553422
rect 57605 553419 57671 553422
rect 108297 552938 108363 552941
rect 105892 552936 108363 552938
rect 105892 552880 108302 552936
rect 108358 552880 108363 552936
rect 105892 552878 108363 552880
rect 108297 552875 108363 552878
rect 67633 552666 67699 552669
rect 67633 552664 70226 552666
rect 67633 552608 67638 552664
rect 67694 552608 70226 552664
rect 67633 552606 70226 552608
rect 67633 552603 67699 552606
rect 70166 552364 70226 552606
rect 108941 552258 109007 552261
rect 105892 552256 109007 552258
rect 105892 552200 108946 552256
rect 109002 552200 109007 552256
rect 105892 552198 109007 552200
rect 108941 552195 109007 552198
rect 67633 551986 67699 551989
rect 67633 551984 70226 551986
rect 67633 551928 67638 551984
rect 67694 551928 70226 551984
rect 67633 551926 70226 551928
rect 67633 551923 67699 551926
rect 70166 551684 70226 551926
rect 108941 551578 109007 551581
rect 105892 551576 109007 551578
rect 105892 551520 108946 551576
rect 109002 551520 109007 551576
rect 105892 551518 109007 551520
rect 108941 551515 109007 551518
rect 68829 551442 68895 551445
rect 68829 551440 70226 551442
rect 68829 551384 68834 551440
rect 68890 551384 70226 551440
rect 68829 551382 70226 551384
rect 68829 551379 68895 551382
rect 70166 551004 70226 551382
rect 106365 551034 106431 551037
rect 106733 551034 106799 551037
rect 105892 551032 106799 551034
rect 105892 550976 106370 551032
rect 106426 550976 106738 551032
rect 106794 550976 106799 551032
rect 583520 551020 584960 551260
rect 105892 550974 106799 550976
rect 106365 550971 106431 550974
rect 106733 550971 106799 550974
rect 108849 550218 108915 550221
rect 105892 550216 108915 550218
rect 70166 549946 70226 550188
rect 105892 550160 108854 550216
rect 108910 550160 108915 550216
rect 105892 550158 108915 550160
rect 108849 550155 108915 550158
rect 109125 549946 109191 549949
rect 122230 549946 122236 549948
rect 64830 549886 70226 549946
rect 105862 549944 122236 549946
rect 105862 549888 109130 549944
rect 109186 549888 122236 549944
rect 105862 549886 122236 549888
rect 64830 549402 64890 549886
rect 105862 549644 105922 549886
rect 109125 549883 109191 549886
rect 122230 549884 122236 549886
rect 122300 549884 122306 549948
rect 60782 549342 64890 549402
rect 67633 549402 67699 549405
rect 70166 549402 70226 549508
rect 67633 549400 70226 549402
rect 67633 549344 67638 549400
rect 67694 549344 70226 549400
rect 67633 549342 70226 549344
rect 33777 549266 33843 549269
rect 34421 549266 34487 549269
rect 60782 549266 60842 549342
rect 67633 549339 67699 549342
rect 33777 549264 60842 549266
rect 33777 549208 33782 549264
rect 33838 549208 34426 549264
rect 34482 549208 60842 549264
rect 33777 549206 60842 549208
rect 67725 549266 67791 549269
rect 68870 549266 68876 549268
rect 67725 549264 68876 549266
rect 67725 549208 67730 549264
rect 67786 549208 68876 549264
rect 67725 549206 68876 549208
rect 33777 549203 33843 549206
rect 34421 549203 34487 549206
rect 67725 549203 67791 549206
rect 68870 549204 68876 549206
rect 68940 549266 68946 549268
rect 68940 549206 70226 549266
rect 68940 549204 68946 549206
rect 70166 548964 70226 549206
rect 108941 548994 109007 548997
rect 105892 548992 109007 548994
rect 105892 548936 108946 548992
rect 109002 548936 109007 548992
rect 105892 548934 109007 548936
rect 108941 548931 109007 548934
rect 67633 548586 67699 548589
rect 67633 548584 70226 548586
rect 67633 548528 67638 548584
rect 67694 548528 70226 548584
rect 67633 548526 70226 548528
rect 67633 548523 67699 548526
rect 70166 548284 70226 548526
rect 108941 547498 109007 547501
rect 105892 547496 109007 547498
rect 67633 547226 67699 547229
rect 70166 547226 70226 547468
rect 105892 547440 108946 547496
rect 109002 547440 109007 547496
rect 105892 547438 109007 547440
rect 108941 547435 109007 547438
rect 67633 547224 70226 547226
rect 67633 547168 67638 547224
rect 67694 547168 70226 547224
rect 67633 547166 70226 547168
rect 67633 547163 67699 547166
rect 108757 546954 108823 546957
rect 111742 546954 111748 546956
rect 105892 546952 111748 546954
rect 105892 546896 108762 546952
rect 108818 546896 111748 546952
rect 105892 546894 111748 546896
rect 108757 546891 108823 546894
rect 111742 546892 111748 546894
rect 111812 546892 111818 546956
rect 67633 546546 67699 546549
rect 70166 546546 70226 546788
rect 67633 546544 70226 546546
rect 67633 546488 67638 546544
rect 67694 546488 70226 546544
rect 67633 546486 70226 546488
rect 67633 546483 67699 546486
rect 37089 546410 37155 546413
rect 60733 546410 60799 546413
rect 61326 546410 61332 546412
rect 37089 546408 61332 546410
rect 37089 546352 37094 546408
rect 37150 546352 60738 546408
rect 60794 546352 61332 546408
rect 37089 546350 61332 546352
rect 37089 546347 37155 546350
rect 60733 546347 60799 546350
rect 61326 546348 61332 546350
rect 61396 546348 61402 546412
rect 65977 546140 66043 546141
rect 65926 546138 65932 546140
rect 65886 546078 65932 546138
rect 65996 546136 66043 546140
rect 108941 546138 109007 546141
rect 66038 546080 66043 546136
rect 65926 546076 65932 546078
rect 65996 546076 66043 546080
rect 105892 546136 109007 546138
rect 105892 546080 108946 546136
rect 109002 546080 109007 546136
rect 105892 546078 109007 546080
rect 65977 546075 66043 546076
rect 108941 546075 109007 546078
rect 108849 545458 108915 545461
rect 105892 545456 108915 545458
rect 67633 545186 67699 545189
rect 70166 545186 70226 545428
rect 105892 545400 108854 545456
rect 108910 545400 108915 545456
rect 105892 545398 108915 545400
rect 108849 545395 108915 545398
rect 67633 545184 70226 545186
rect 67633 545128 67638 545184
rect 67694 545128 70226 545184
rect 67633 545126 70226 545128
rect 115197 545186 115263 545189
rect 115790 545186 115796 545188
rect 115197 545184 115796 545186
rect 115197 545128 115202 545184
rect 115258 545128 115796 545184
rect 115197 545126 115796 545128
rect 67633 545123 67699 545126
rect 115197 545123 115263 545126
rect 115790 545124 115796 545126
rect 115860 545186 115866 545188
rect 118785 545186 118851 545189
rect 115860 545184 118851 545186
rect 115860 545128 118790 545184
rect 118846 545128 118851 545184
rect 115860 545126 118851 545128
rect 115860 545124 115866 545126
rect 118785 545123 118851 545126
rect 108941 544778 109007 544781
rect 105892 544776 109007 544778
rect 68829 544506 68895 544509
rect 70166 544506 70226 544748
rect 105892 544720 108946 544776
rect 109002 544720 109007 544776
rect 105892 544718 109007 544720
rect 108941 544715 109007 544718
rect 68829 544504 70226 544506
rect 68829 544448 68834 544504
rect 68890 544448 70226 544504
rect 68829 544446 70226 544448
rect 68829 544443 68895 544446
rect 55070 544308 55076 544372
rect 55140 544370 55146 544372
rect 69841 544370 69907 544373
rect 55140 544368 69907 544370
rect 55140 544312 69846 544368
rect 69902 544312 69907 544368
rect 55140 544310 69907 544312
rect 55140 544308 55146 544310
rect 69841 544307 69907 544310
rect 108849 544098 108915 544101
rect 105892 544096 108915 544098
rect 68185 543826 68251 543829
rect 68553 543826 68619 543829
rect 70166 543826 70226 544068
rect 105892 544040 108854 544096
rect 108910 544040 108915 544096
rect 105892 544038 108915 544040
rect 108849 544035 108915 544038
rect 68185 543824 70226 543826
rect 68185 543768 68190 543824
rect 68246 543768 68558 543824
rect 68614 543768 70226 543824
rect 68185 543766 70226 543768
rect 68185 543763 68251 543766
rect 68553 543763 68619 543766
rect 108941 543554 109007 543557
rect 105892 543552 109007 543554
rect 105892 543496 108946 543552
rect 109002 543496 109007 543552
rect 105892 543494 109007 543496
rect 108941 543491 109007 543494
rect 67633 543282 67699 543285
rect 70166 543282 70226 543388
rect 67633 543280 70226 543282
rect 67633 543224 67638 543280
rect 67694 543224 70226 543280
rect 67633 543222 70226 543224
rect 67633 543219 67699 543222
rect 67725 543146 67791 543149
rect 67725 543144 70226 543146
rect 67725 543088 67730 543144
rect 67786 543088 70226 543144
rect 67725 543086 70226 543088
rect 67725 543083 67791 543086
rect 56409 543010 56475 543013
rect 57830 543010 57836 543012
rect 56409 543008 57836 543010
rect 56409 542952 56414 543008
rect 56470 542952 57836 543008
rect 56409 542950 57836 542952
rect 56409 542947 56475 542950
rect 57830 542948 57836 542950
rect 57900 543010 57906 543012
rect 60733 543010 60799 543013
rect 57900 543008 60799 543010
rect 57900 542952 60738 543008
rect 60794 542952 60799 543008
rect 57900 542950 60799 542952
rect 57900 542948 57906 542950
rect 60733 542947 60799 542950
rect 70166 542844 70226 543086
rect 107653 542874 107719 542877
rect 109166 542874 109172 542876
rect 105892 542872 109172 542874
rect 105892 542816 107658 542872
rect 107714 542816 109172 542872
rect 105892 542814 109172 542816
rect 107653 542811 107719 542814
rect 109166 542812 109172 542814
rect 109236 542812 109242 542876
rect 108849 542058 108915 542061
rect 105892 542056 108915 542058
rect 65926 541724 65932 541788
rect 65996 541786 66002 541788
rect 70166 541786 70226 542028
rect 105892 542000 108854 542056
rect 108910 542000 108915 542056
rect 105892 541998 108915 542000
rect 108849 541995 108915 541998
rect 65996 541726 70226 541786
rect 65996 541724 66002 541726
rect 67633 541242 67699 541245
rect 70166 541242 70226 541348
rect 67633 541240 70226 541242
rect 67633 541184 67638 541240
rect 67694 541184 70226 541240
rect 67633 541182 70226 541184
rect 67633 541179 67699 541182
rect -960 540684 480 540924
rect 108941 540834 109007 540837
rect 105892 540832 109007 540834
rect 105892 540776 108946 540832
rect 109002 540776 109007 540832
rect 105892 540774 109007 540776
rect 108941 540771 109007 540774
rect 67633 540562 67699 540565
rect 70166 540562 70226 540668
rect 67633 540560 70226 540562
rect 67633 540504 67638 540560
rect 67694 540504 70226 540560
rect 67633 540502 70226 540504
rect 67633 540499 67699 540502
rect 108021 540018 108087 540021
rect 105892 540016 108087 540018
rect 105892 539988 108026 540016
rect 105862 539960 108026 539988
rect 108082 539960 108087 540016
rect 105862 539958 108087 539960
rect 104801 539882 104867 539885
rect 104934 539882 104940 539884
rect 104801 539880 104940 539882
rect 104801 539824 104806 539880
rect 104862 539824 104940 539880
rect 104801 539822 104940 539824
rect 104801 539819 104867 539822
rect 104934 539820 104940 539822
rect 105004 539820 105010 539884
rect 105862 539613 105922 539958
rect 108021 539955 108087 539958
rect 105813 539608 105922 539613
rect 105813 539552 105818 539608
rect 105874 539552 105922 539608
rect 105813 539550 105922 539552
rect 105813 539547 105879 539550
rect 50838 539412 50844 539476
rect 50908 539474 50914 539476
rect 52361 539474 52427 539477
rect 50908 539472 52427 539474
rect 50908 539416 52366 539472
rect 52422 539416 52427 539472
rect 50908 539414 52427 539416
rect 50908 539412 50914 539414
rect 52361 539411 52427 539414
rect 61377 538794 61443 538797
rect 70342 538794 70348 538796
rect 61377 538792 70348 538794
rect 61377 538736 61382 538792
rect 61438 538736 70348 538792
rect 61377 538734 70348 538736
rect 61377 538731 61443 538734
rect 70342 538732 70348 538734
rect 70412 538732 70418 538796
rect 94037 538794 94103 538797
rect 125726 538794 125732 538796
rect 94037 538792 125732 538794
rect 94037 538736 94042 538792
rect 94098 538736 125732 538792
rect 94037 538734 125732 538736
rect 94037 538731 94103 538734
rect 125726 538732 125732 538734
rect 125796 538732 125802 538796
rect 57789 538114 57855 538117
rect 81617 538114 81683 538117
rect 57789 538112 81683 538114
rect 57789 538056 57794 538112
rect 57850 538056 81622 538112
rect 81678 538056 81683 538112
rect 57789 538054 81683 538056
rect 57789 538051 57855 538054
rect 81617 538051 81683 538054
rect 99649 538114 99715 538117
rect 105445 538114 105511 538117
rect 106273 538114 106339 538117
rect 99649 538112 106339 538114
rect 99649 538056 99654 538112
rect 99710 538056 105450 538112
rect 105506 538056 106278 538112
rect 106334 538056 106339 538112
rect 99649 538054 106339 538056
rect 99649 538051 99715 538054
rect 105445 538051 105511 538054
rect 106273 538051 106339 538054
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect 58934 537372 58940 537436
rect 59004 537434 59010 537436
rect 74533 537434 74599 537437
rect 59004 537432 74599 537434
rect 59004 537376 74538 537432
rect 74594 537376 74599 537432
rect 59004 537374 74599 537376
rect 59004 537372 59010 537374
rect 74533 537371 74599 537374
rect 104157 536890 104223 536893
rect 104801 536890 104867 536893
rect 104157 536888 104867 536890
rect 104157 536832 104162 536888
rect 104218 536832 104806 536888
rect 104862 536832 104867 536888
rect 104157 536830 104867 536832
rect 104157 536827 104223 536830
rect 104801 536827 104867 536830
rect 70158 536692 70164 536756
rect 70228 536754 70234 536756
rect 91921 536754 91987 536757
rect 70228 536752 91987 536754
rect 70228 536696 91926 536752
rect 91982 536696 91987 536752
rect 70228 536694 91987 536696
rect 70228 536692 70234 536694
rect 91921 536691 91987 536694
rect 99373 536754 99439 536757
rect 111558 536754 111564 536756
rect 99373 536752 111564 536754
rect 99373 536696 99378 536752
rect 99434 536696 111564 536752
rect 99373 536694 111564 536696
rect 99373 536691 99439 536694
rect 111558 536692 111564 536694
rect 111628 536754 111634 536756
rect 111628 536694 113190 536754
rect 111628 536692 111634 536694
rect 113130 536346 113190 536694
rect 114686 536346 114692 536348
rect 113130 536286 114692 536346
rect 114686 536284 114692 536286
rect 114756 536284 114762 536348
rect 125542 535468 125548 535532
rect 125612 535530 125618 535532
rect 125961 535530 126027 535533
rect 125612 535528 126027 535530
rect 125612 535472 125966 535528
rect 126022 535472 126027 535528
rect 125612 535470 126027 535472
rect 125612 535468 125618 535470
rect 125961 535467 126027 535470
rect 49325 534170 49391 534173
rect 50838 534170 50844 534172
rect 49325 534168 50844 534170
rect 49325 534112 49330 534168
rect 49386 534112 50844 534168
rect 49325 534110 50844 534112
rect 49325 534107 49391 534110
rect 50838 534108 50844 534110
rect 50908 534108 50914 534172
rect 54886 533836 54892 533900
rect 54956 533898 54962 533900
rect 56542 533898 56548 533900
rect 54956 533838 56548 533898
rect 54956 533836 54962 533838
rect 56542 533836 56548 533838
rect 56612 533898 56618 533900
rect 57881 533898 57947 533901
rect 56612 533896 57947 533898
rect 56612 533840 57886 533896
rect 57942 533840 57947 533896
rect 56612 533838 57947 533840
rect 56612 533836 56618 533838
rect 57881 533835 57947 533838
rect 55029 533628 55095 533629
rect 55029 533624 55076 533628
rect 55140 533626 55146 533628
rect 55029 533568 55034 533624
rect 55029 533564 55076 533568
rect 55140 533566 55186 533626
rect 55140 533564 55146 533566
rect 55029 533563 55095 533564
rect 97809 533354 97875 533357
rect 114502 533354 114508 533356
rect 97809 533352 114508 533354
rect 97809 533296 97814 533352
rect 97870 533296 114508 533352
rect 97809 533294 114508 533296
rect 97809 533291 97875 533294
rect 114502 533292 114508 533294
rect 114572 533292 114578 533356
rect 99189 532266 99255 532269
rect 125542 532266 125548 532268
rect 99189 532264 125548 532266
rect 99189 532208 99194 532264
rect 99250 532208 125548 532264
rect 99189 532206 125548 532208
rect 99189 532203 99255 532206
rect 125542 532204 125548 532206
rect 125612 532204 125618 532268
rect 93669 532130 93735 532133
rect 120022 532130 120028 532132
rect 93669 532128 120028 532130
rect 93669 532072 93674 532128
rect 93730 532072 120028 532128
rect 93669 532070 120028 532072
rect 93669 532067 93735 532070
rect 120022 532068 120028 532070
rect 120092 532068 120098 532132
rect 86953 531994 87019 531997
rect 128670 531994 128676 531996
rect 86953 531992 128676 531994
rect 86953 531936 86958 531992
rect 87014 531936 128676 531992
rect 86953 531934 128676 531936
rect 86953 531931 87019 531934
rect 128670 531932 128676 531934
rect 128740 531932 128746 531996
rect -960 527914 480 528004
rect 3141 527914 3207 527917
rect -960 527912 3207 527914
rect -960 527856 3146 527912
rect 3202 527856 3207 527912
rect -960 527854 3207 527856
rect -960 527764 480 527854
rect 3141 527851 3207 527854
rect 37181 525738 37247 525741
rect 65926 525738 65932 525740
rect 37181 525736 65932 525738
rect 37181 525680 37186 525736
rect 37242 525680 65932 525736
rect 37181 525678 65932 525680
rect 37181 525675 37247 525678
rect 65926 525676 65932 525678
rect 65996 525676 66002 525740
rect 65926 524452 65932 524516
rect 65996 524514 66002 524516
rect 583520 524514 584960 524604
rect 65996 524454 584960 524514
rect 65996 524452 66002 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3141 501802 3207 501805
rect -960 501800 3207 501802
rect -960 501744 3146 501800
rect 3202 501744 3207 501800
rect -960 501742 3207 501744
rect -960 501652 480 501742
rect 3141 501739 3207 501742
rect 86217 498810 86283 498813
rect 118918 498810 118924 498812
rect 86217 498808 118924 498810
rect 86217 498752 86222 498808
rect 86278 498752 118924 498808
rect 86217 498750 118924 498752
rect 86217 498747 86283 498750
rect 118918 498748 118924 498750
rect 118988 498748 118994 498812
rect 121453 498266 121519 498269
rect 122046 498266 122052 498268
rect 121453 498264 122052 498266
rect 121453 498208 121458 498264
rect 121514 498208 122052 498264
rect 121453 498206 122052 498208
rect 121453 498203 121519 498206
rect 122046 498204 122052 498206
rect 122116 498204 122122 498268
rect 583520 497844 584960 498084
rect 84837 497450 84903 497453
rect 115974 497450 115980 497452
rect 84837 497448 115980 497450
rect 84837 497392 84842 497448
rect 84898 497392 115980 497448
rect 84837 497390 115980 497392
rect 84837 497387 84903 497390
rect 115974 497388 115980 497390
rect 116044 497450 116050 497452
rect 117589 497450 117655 497453
rect 116044 497448 117655 497450
rect 116044 497392 117594 497448
rect 117650 497392 117655 497448
rect 116044 497390 117655 497392
rect 116044 497388 116050 497390
rect 117589 497387 117655 497390
rect 83457 496090 83523 496093
rect 110638 496090 110644 496092
rect 83457 496088 110644 496090
rect 83457 496032 83462 496088
rect 83518 496032 110644 496088
rect 83457 496030 110644 496032
rect 83457 496027 83523 496030
rect 110638 496028 110644 496030
rect 110708 496028 110714 496092
rect 124305 495548 124371 495549
rect 124254 495546 124260 495548
rect 124214 495486 124260 495546
rect 124324 495544 124371 495548
rect 124366 495488 124371 495544
rect 124254 495484 124260 495486
rect 124324 495484 124371 495488
rect 124305 495483 124371 495484
rect 76465 494730 76531 494733
rect 117998 494730 118004 494732
rect 76465 494728 118004 494730
rect 76465 494672 76470 494728
rect 76526 494672 118004 494728
rect 76465 494670 118004 494672
rect 76465 494667 76531 494670
rect 117998 494668 118004 494670
rect 118068 494730 118074 494732
rect 122833 494730 122899 494733
rect 118068 494728 122899 494730
rect 118068 494672 122838 494728
rect 122894 494672 122899 494728
rect 118068 494670 122899 494672
rect 118068 494668 118074 494670
rect 122833 494667 122899 494670
rect 95785 493370 95851 493373
rect 113214 493370 113220 493372
rect 95785 493368 113220 493370
rect 95785 493312 95790 493368
rect 95846 493312 113220 493368
rect 95785 493310 113220 493312
rect 95785 493307 95851 493310
rect 113214 493308 113220 493310
rect 113284 493370 113290 493372
rect 114461 493370 114527 493373
rect 113284 493368 114527 493370
rect 113284 493312 114466 493368
rect 114522 493312 114527 493368
rect 113284 493310 114527 493312
rect 113284 493308 113290 493310
rect 114461 493307 114527 493310
rect 57830 492764 57836 492828
rect 57900 492826 57906 492828
rect 70853 492826 70919 492829
rect 74993 492826 75059 492829
rect 57900 492824 70919 492826
rect 57900 492768 70858 492824
rect 70914 492768 70919 492824
rect 57900 492766 70919 492768
rect 57900 492764 57906 492766
rect 70853 492763 70919 492766
rect 74490 492824 75059 492826
rect 74490 492768 74998 492824
rect 75054 492768 75059 492824
rect 74490 492766 75059 492768
rect 53598 492628 53604 492692
rect 53668 492690 53674 492692
rect 74490 492690 74550 492766
rect 74993 492763 75059 492766
rect 79685 492826 79751 492829
rect 112294 492826 112300 492828
rect 79685 492824 112300 492826
rect 79685 492768 79690 492824
rect 79746 492768 112300 492824
rect 79685 492766 112300 492768
rect 79685 492763 79751 492766
rect 112294 492764 112300 492766
rect 112364 492826 112370 492828
rect 112364 492766 113190 492826
rect 112364 492764 112370 492766
rect 53668 492630 74550 492690
rect 53668 492628 53674 492630
rect 113130 492554 113190 492766
rect 118734 492554 118740 492556
rect 113130 492494 118740 492554
rect 118734 492492 118740 492494
rect 118804 492492 118810 492556
rect 95049 491466 95115 491469
rect 99230 491466 99236 491468
rect 95049 491464 99236 491466
rect 95049 491408 95054 491464
rect 95110 491408 99236 491464
rect 95049 491406 99236 491408
rect 95049 491403 95115 491406
rect 99230 491404 99236 491406
rect 99300 491404 99306 491468
rect 97073 491330 97139 491333
rect 109125 491330 109191 491333
rect 97073 491328 109191 491330
rect 97073 491272 97078 491328
rect 97134 491272 109130 491328
rect 109186 491272 109191 491328
rect 97073 491270 109191 491272
rect 97073 491267 97139 491270
rect 109125 491267 109191 491270
rect 110505 491194 110571 491197
rect 111558 491194 111564 491196
rect 110505 491192 111564 491194
rect 110505 491136 110510 491192
rect 110566 491136 111564 491192
rect 110505 491134 111564 491136
rect 110505 491131 110571 491134
rect 111558 491132 111564 491134
rect 111628 491194 111634 491196
rect 136817 491194 136883 491197
rect 111628 491192 136883 491194
rect 111628 491136 136822 491192
rect 136878 491136 136883 491192
rect 111628 491134 136883 491136
rect 111628 491132 111634 491134
rect 136817 491131 136883 491134
rect 87367 490106 87433 490109
rect 101254 490106 101260 490108
rect 87367 490104 101260 490106
rect 87367 490048 87372 490104
rect 87428 490048 101260 490104
rect 87367 490046 101260 490048
rect 87367 490043 87433 490046
rect 101254 490044 101260 490046
rect 101324 490044 101330 490108
rect 94129 489970 94195 489973
rect 109677 489970 109743 489973
rect 94129 489968 109743 489970
rect 94129 489912 94134 489968
rect 94190 489912 109682 489968
rect 109738 489912 109743 489968
rect 94129 489910 109743 489912
rect 94129 489907 94195 489910
rect 109677 489907 109743 489910
rect 48078 489772 48084 489836
rect 48148 489834 48154 489836
rect 48957 489834 49023 489837
rect 48148 489832 49023 489834
rect 48148 489776 48962 489832
rect 49018 489776 49023 489832
rect 48148 489774 49023 489776
rect 48148 489772 48154 489774
rect 48957 489771 49023 489774
rect 67725 489154 67791 489157
rect 70166 489154 70226 489668
rect 67725 489152 70226 489154
rect 67725 489096 67730 489152
rect 67786 489096 70226 489152
rect 67725 489094 70226 489096
rect 67725 489091 67791 489094
rect -960 488596 480 488836
rect 50286 488548 50292 488612
rect 50356 488610 50362 488612
rect 51758 488610 51764 488612
rect 50356 488550 51764 488610
rect 50356 488548 50362 488550
rect 51758 488548 51764 488550
rect 51828 488610 51834 488612
rect 52177 488610 52243 488613
rect 51828 488608 52243 488610
rect 51828 488552 52182 488608
rect 52238 488552 52243 488608
rect 51828 488550 52243 488552
rect 99790 488610 99850 488988
rect 103421 488610 103487 488613
rect 99790 488608 103487 488610
rect 99790 488552 103426 488608
rect 103482 488552 103487 488608
rect 99790 488550 103487 488552
rect 51828 488548 51834 488550
rect 52177 488547 52243 488550
rect 103421 488547 103487 488550
rect 117221 488474 117287 488477
rect 122598 488474 122604 488476
rect 117221 488472 122604 488474
rect 117221 488416 117226 488472
rect 117282 488416 122604 488472
rect 117221 488414 122604 488416
rect 117221 488411 117287 488414
rect 122598 488412 122604 488414
rect 122668 488412 122674 488476
rect 67633 488066 67699 488069
rect 70350 488066 70410 488308
rect 67633 488064 70410 488066
rect 67633 488008 67638 488064
rect 67694 488008 70410 488064
rect 67633 488006 70410 488008
rect 67633 488003 67699 488006
rect 67633 487930 67699 487933
rect 99606 487930 99666 488308
rect 103421 487930 103487 487933
rect 67633 487928 70226 487930
rect 67633 487872 67638 487928
rect 67694 487872 70226 487928
rect 67633 487870 70226 487872
rect 99606 487928 103487 487930
rect 99606 487872 103426 487928
rect 103482 487872 103487 487928
rect 99606 487870 103487 487872
rect 67633 487867 67699 487870
rect 70166 487764 70226 487870
rect 103421 487867 103487 487870
rect 99606 487386 99666 487628
rect 103329 487386 103395 487389
rect 99606 487384 103395 487386
rect 99606 487328 103334 487384
rect 103390 487328 103395 487384
rect 99606 487326 103395 487328
rect 103329 487323 103395 487326
rect 102777 487250 102843 487253
rect 99790 487248 102843 487250
rect 99790 487192 102782 487248
rect 102838 487192 102843 487248
rect 99790 487190 102843 487192
rect 99790 487084 99850 487190
rect 102777 487187 102843 487190
rect 67725 486570 67791 486573
rect 70166 486570 70226 486948
rect 103329 486570 103395 486573
rect 67725 486568 70226 486570
rect 67725 486512 67730 486568
rect 67786 486512 70226 486568
rect 67725 486510 70226 486512
rect 99790 486568 103395 486570
rect 99790 486512 103334 486568
rect 103390 486512 103395 486568
rect 99790 486510 103395 486512
rect 67725 486507 67791 486510
rect 99790 486404 99850 486510
rect 103329 486507 103395 486510
rect 67633 485890 67699 485893
rect 70166 485890 70226 486268
rect 99322 485964 99328 486028
rect 99392 486026 99398 486028
rect 106917 486026 106983 486029
rect 99392 486024 106983 486026
rect 99392 485968 106922 486024
rect 106978 485968 106983 486024
rect 99392 485966 106983 485968
rect 99392 485964 99398 485966
rect 106917 485963 106983 485966
rect 67633 485888 70226 485890
rect 67633 485832 67638 485888
rect 67694 485832 70226 485888
rect 67633 485830 70226 485832
rect 67633 485827 67699 485830
rect 117078 485692 117084 485756
rect 117148 485754 117154 485756
rect 117221 485754 117287 485757
rect 117148 485752 117287 485754
rect 117148 485696 117226 485752
rect 117282 485696 117287 485752
rect 117148 485694 117287 485696
rect 117148 485692 117154 485694
rect 117221 485691 117287 485694
rect 67633 485210 67699 485213
rect 70166 485210 70226 485588
rect 99790 485346 99850 485588
rect 102409 485346 102475 485349
rect 99790 485344 102475 485346
rect 99790 485288 102414 485344
rect 102470 485288 102475 485344
rect 99790 485286 102475 485288
rect 102409 485283 102475 485286
rect 102133 485210 102199 485213
rect 67633 485208 70226 485210
rect 67633 485152 67638 485208
rect 67694 485152 70226 485208
rect 67633 485150 70226 485152
rect 99790 485208 102199 485210
rect 99790 485152 102138 485208
rect 102194 485152 102199 485208
rect 99790 485150 102199 485152
rect 67633 485147 67699 485150
rect 99790 485044 99850 485150
rect 102133 485147 102199 485150
rect 114461 485074 114527 485077
rect 117405 485074 117471 485077
rect 142245 485074 142311 485077
rect 114461 485072 142311 485074
rect 114461 485016 114466 485072
rect 114522 485016 117410 485072
rect 117466 485016 142250 485072
rect 142306 485016 142311 485072
rect 114461 485014 142311 485016
rect 114461 485011 114527 485014
rect 117405 485011 117471 485014
rect 142245 485011 142311 485014
rect 68461 484666 68527 484669
rect 70166 484666 70226 484908
rect 70342 484666 70348 484668
rect 68461 484664 70348 484666
rect 68461 484608 68466 484664
rect 68522 484608 70348 484664
rect 68461 484606 70348 484608
rect 68461 484603 68527 484606
rect 70342 484604 70348 484606
rect 70412 484604 70418 484668
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 107510 484468 107516 484532
rect 107580 484530 107586 484532
rect 123334 484530 123340 484532
rect 107580 484470 123340 484530
rect 107580 484468 107586 484470
rect 123334 484468 123340 484470
rect 123404 484468 123410 484532
rect 583520 484516 584960 484606
rect 67633 483986 67699 483989
rect 70166 483986 70226 484228
rect 67633 483984 70226 483986
rect 67633 483928 67638 483984
rect 67694 483928 70226 483984
rect 67633 483926 70226 483928
rect 67633 483923 67699 483926
rect 99790 483170 99850 483548
rect 107510 483170 107516 483172
rect 99790 483110 107516 483170
rect 107510 483108 107516 483110
rect 107580 483108 107586 483172
rect 107510 482972 107516 483036
rect 107580 483034 107586 483036
rect 140957 483034 141023 483037
rect 107580 483032 141023 483034
rect 107580 482976 140962 483032
rect 141018 482976 141023 483032
rect 107580 482974 141023 482976
rect 107580 482972 107586 482974
rect 140957 482971 141023 482974
rect 68921 482626 68987 482629
rect 69105 482626 69171 482629
rect 70350 482626 70410 482868
rect 68921 482624 70410 482626
rect 68921 482568 68926 482624
rect 68982 482568 69110 482624
rect 69166 482568 70410 482624
rect 68921 482566 70410 482568
rect 99606 482626 99666 482868
rect 102133 482626 102199 482629
rect 99606 482624 102199 482626
rect 99606 482568 102138 482624
rect 102194 482568 102199 482624
rect 99606 482566 102199 482568
rect 68921 482563 68987 482566
rect 69105 482563 69171 482566
rect 102133 482563 102199 482566
rect 68001 482490 68067 482493
rect 69013 482490 69079 482493
rect 68001 482488 70226 482490
rect 68001 482432 68006 482488
rect 68062 482432 69018 482488
rect 69074 482432 70226 482488
rect 68001 482430 70226 482432
rect 68001 482427 68067 482430
rect 69013 482427 69079 482430
rect 70166 482324 70226 482430
rect 99790 481810 99850 482188
rect 107510 481810 107516 481812
rect 99790 481750 107516 481810
rect 107510 481748 107516 481750
rect 107580 481748 107586 481812
rect 64638 481476 64644 481540
rect 64708 481538 64714 481540
rect 68093 481538 68159 481541
rect 64708 481536 68159 481538
rect 64708 481480 68098 481536
rect 68154 481480 68159 481536
rect 64708 481478 68159 481480
rect 64708 481476 64714 481478
rect 68093 481475 68159 481478
rect 67633 481130 67699 481133
rect 70166 481130 70226 481508
rect 67633 481128 70226 481130
rect 67633 481072 67638 481128
rect 67694 481072 70226 481128
rect 67633 481070 70226 481072
rect 99606 481130 99666 481508
rect 106774 481476 106780 481540
rect 106844 481538 106850 481540
rect 109033 481538 109099 481541
rect 106844 481536 109099 481538
rect 106844 481480 109038 481536
rect 109094 481480 109099 481536
rect 106844 481478 109099 481480
rect 106844 481476 106850 481478
rect 109033 481475 109099 481478
rect 102133 481130 102199 481133
rect 99606 481128 102199 481130
rect 99606 481072 102138 481128
rect 102194 481072 102199 481128
rect 99606 481070 102199 481072
rect 67633 481067 67699 481070
rect 102133 481067 102199 481070
rect 68093 480586 68159 480589
rect 69197 480586 69263 480589
rect 70350 480586 70410 480828
rect 68093 480584 70410 480586
rect 68093 480528 68098 480584
rect 68154 480528 69202 480584
rect 69258 480528 70410 480584
rect 68093 480526 70410 480528
rect 99606 480586 99666 480828
rect 102225 480586 102291 480589
rect 99606 480584 102291 480586
rect 99606 480528 102230 480584
rect 102286 480528 102291 480584
rect 99606 480526 102291 480528
rect 68093 480523 68159 480526
rect 69197 480523 69263 480526
rect 102225 480523 102291 480526
rect 99790 480210 100034 480270
rect 99790 480148 99850 480210
rect 99974 480178 100034 480210
rect 105486 480178 105492 480180
rect 67633 479770 67699 479773
rect 70166 479770 70226 480148
rect 99974 480118 105492 480178
rect 105486 480116 105492 480118
rect 105556 480116 105562 480180
rect 102133 479906 102199 479909
rect 67633 479768 70226 479770
rect 67633 479712 67638 479768
rect 67694 479712 70226 479768
rect 67633 479710 70226 479712
rect 99790 479904 102199 479906
rect 99790 479848 102138 479904
rect 102194 479848 102199 479904
rect 99790 479846 102199 479848
rect 67633 479707 67699 479710
rect 99790 479604 99850 479846
rect 102133 479843 102199 479846
rect 67541 479226 67607 479229
rect 70350 479226 70410 479468
rect 67541 479224 70410 479226
rect 67541 479168 67546 479224
rect 67602 479168 70410 479224
rect 67541 479166 70410 479168
rect 67541 479163 67607 479166
rect 105537 479092 105603 479093
rect 105486 479090 105492 479092
rect 105446 479030 105492 479090
rect 105556 479088 105603 479092
rect 105598 479032 105603 479088
rect 105486 479028 105492 479030
rect 105556 479028 105603 479032
rect 105537 479027 105603 479028
rect 106181 478954 106247 478957
rect 107878 478954 107884 478956
rect 106181 478952 107884 478954
rect 106181 478896 106186 478952
rect 106242 478896 107884 478952
rect 106181 478894 107884 478896
rect 106181 478891 106247 478894
rect 107878 478892 107884 478894
rect 107948 478892 107954 478956
rect 67633 478274 67699 478277
rect 70166 478274 70226 478788
rect 67633 478272 70226 478274
rect 67633 478216 67638 478272
rect 67694 478216 70226 478272
rect 67633 478214 70226 478216
rect 67633 478211 67699 478214
rect 99790 477730 99850 478108
rect 103421 477730 103487 477733
rect 99790 477728 103487 477730
rect 99790 477672 103426 477728
rect 103482 477672 103487 477728
rect 99790 477670 103487 477672
rect 103421 477667 103487 477670
rect 63033 477596 63099 477597
rect 62982 477594 62988 477596
rect 62942 477534 62988 477594
rect 63052 477592 63099 477596
rect 63094 477536 63099 477592
rect 62982 477532 62988 477534
rect 63052 477532 63099 477536
rect 63033 477531 63099 477532
rect 68645 477050 68711 477053
rect 70166 477050 70226 477428
rect 99790 477186 99850 477428
rect 102317 477186 102383 477189
rect 99790 477184 102383 477186
rect 99790 477128 102322 477184
rect 102378 477128 102383 477184
rect 99790 477126 102383 477128
rect 102317 477123 102383 477126
rect 102133 477050 102199 477053
rect 68645 477048 70226 477050
rect 68645 476992 68650 477048
rect 68706 476992 70226 477048
rect 68645 476990 70226 476992
rect 99790 477048 102199 477050
rect 99790 476992 102138 477048
rect 102194 476992 102199 477048
rect 99790 476990 102199 476992
rect 68645 476987 68711 476990
rect 99790 476884 99850 476990
rect 102133 476987 102199 476990
rect 67633 476506 67699 476509
rect 70166 476506 70226 476748
rect 102225 476506 102291 476509
rect 67633 476504 70226 476506
rect 67633 476448 67638 476504
rect 67694 476448 70226 476504
rect 67633 476446 70226 476448
rect 99790 476504 102291 476506
rect 99790 476448 102230 476504
rect 102286 476448 102291 476504
rect 99790 476446 102291 476448
rect 67633 476443 67699 476446
rect 61694 476308 61700 476372
rect 61764 476370 61770 476372
rect 62982 476370 62988 476372
rect 61764 476310 62988 476370
rect 61764 476308 61770 476310
rect 62982 476308 62988 476310
rect 63052 476370 63058 476372
rect 63052 476310 70226 476370
rect 63052 476308 63058 476310
rect 70166 476204 70226 476310
rect 99790 476204 99850 476446
rect 102225 476443 102291 476446
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 67633 475690 67699 475693
rect 102133 475690 102199 475693
rect 67633 475688 70226 475690
rect 67633 475632 67638 475688
rect 67694 475632 70226 475688
rect 67633 475630 70226 475632
rect 67633 475627 67699 475630
rect 70166 475524 70226 475630
rect 99790 475688 102199 475690
rect 99790 475632 102138 475688
rect 102194 475632 102199 475688
rect 99790 475630 102199 475632
rect 99790 475524 99850 475630
rect 102133 475627 102199 475630
rect 67725 475010 67791 475013
rect 102133 475010 102199 475013
rect 67725 475008 70226 475010
rect 67725 474952 67730 475008
rect 67786 474952 70226 475008
rect 67725 474950 70226 474952
rect 67725 474947 67791 474950
rect 70166 474844 70226 474950
rect 99790 475008 102199 475010
rect 99790 474952 102138 475008
rect 102194 474952 102199 475008
rect 99790 474950 102199 474952
rect 99790 474844 99850 474950
rect 102133 474947 102199 474950
rect 102225 474330 102291 474333
rect 99790 474328 102291 474330
rect 99790 474272 102230 474328
rect 102286 474272 102291 474328
rect 99790 474270 102291 474272
rect 99790 474164 99850 474270
rect 102225 474267 102291 474270
rect 66662 473786 66668 473788
rect 60690 473726 66668 473786
rect 59118 473452 59124 473516
rect 59188 473514 59194 473516
rect 60690 473514 60750 473726
rect 66662 473724 66668 473726
rect 66732 473786 66738 473788
rect 68921 473786 68987 473789
rect 66732 473784 68987 473786
rect 66732 473728 68926 473784
rect 68982 473728 68987 473784
rect 66732 473726 68987 473728
rect 66732 473724 66738 473726
rect 68921 473723 68987 473726
rect 70166 473650 70226 474028
rect 59188 473454 60750 473514
rect 65566 473590 70226 473650
rect 59188 473452 59194 473454
rect 60590 473316 60596 473380
rect 60660 473378 60666 473380
rect 65566 473378 65626 473590
rect 60660 473318 65626 473378
rect 68921 473378 68987 473381
rect 68921 473376 70042 473378
rect 68921 473320 68926 473376
rect 68982 473370 70042 473376
rect 68982 473320 70226 473370
rect 68921 473318 70226 473320
rect 60660 473316 60666 473318
rect 68921 473315 68987 473318
rect 69982 473310 70226 473318
rect 102133 472970 102199 472973
rect 99790 472968 102199 472970
rect 99790 472912 102138 472968
rect 102194 472912 102199 472968
rect 99790 472910 102199 472912
rect 99790 472804 99850 472910
rect 102133 472907 102199 472910
rect 67633 472698 67699 472701
rect 67633 472696 70226 472698
rect 67633 472640 67638 472696
rect 67694 472640 70226 472696
rect 67633 472638 70226 472640
rect 67633 472635 67699 472638
rect 70166 472124 70226 472638
rect 102133 472290 102199 472293
rect 99790 472288 102199 472290
rect 99790 472232 102138 472288
rect 102194 472232 102199 472288
rect 99790 472230 102199 472232
rect 99790 472124 99850 472230
rect 102133 472227 102199 472230
rect 66110 471548 66116 471612
rect 66180 471610 66186 471612
rect 102133 471610 102199 471613
rect 66180 471550 70226 471610
rect 66180 471548 66186 471550
rect 70166 471444 70226 471550
rect 99790 471608 102199 471610
rect 99790 471552 102138 471608
rect 102194 471552 102199 471608
rect 99790 471550 102199 471552
rect 99790 471444 99850 471550
rect 102133 471547 102199 471550
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 67725 471066 67791 471069
rect 67725 471064 70226 471066
rect 67725 471008 67730 471064
rect 67786 471008 70226 471064
rect 67725 471006 70226 471008
rect 67725 471003 67791 471006
rect 70166 470764 70226 471006
rect 102133 470930 102199 470933
rect 99790 470928 102199 470930
rect 99790 470872 102138 470928
rect 102194 470872 102199 470928
rect 99790 470870 102199 470872
rect 99790 470764 99850 470870
rect 102133 470867 102199 470870
rect 67633 470250 67699 470253
rect 101949 470250 102015 470253
rect 67633 470248 70226 470250
rect 67633 470192 67638 470248
rect 67694 470192 70226 470248
rect 67633 470190 70226 470192
rect 67633 470187 67699 470190
rect 70166 470084 70226 470190
rect 99790 470248 102015 470250
rect 99790 470192 101954 470248
rect 102010 470192 102015 470248
rect 99790 470190 102015 470192
rect 99790 470084 99850 470190
rect 101949 470187 102015 470190
rect 67725 469706 67791 469709
rect 67725 469704 70226 469706
rect 67725 469648 67730 469704
rect 67786 469648 70226 469704
rect 67725 469646 70226 469648
rect 67725 469643 67791 469646
rect 70166 469404 70226 469646
rect 102133 469570 102199 469573
rect 99790 469568 102199 469570
rect 99790 469512 102138 469568
rect 102194 469512 102199 469568
rect 99790 469510 102199 469512
rect 99790 469404 99850 469510
rect 102133 469507 102199 469510
rect 108389 469298 108455 469301
rect 114686 469298 114692 469300
rect 108389 469296 114692 469298
rect 108389 469240 108394 469296
rect 108450 469240 114692 469296
rect 108389 469238 114692 469240
rect 108389 469235 108455 469238
rect 114686 469236 114692 469238
rect 114756 469236 114762 469300
rect 67633 468890 67699 468893
rect 102133 468890 102199 468893
rect 67633 468888 70226 468890
rect 67633 468832 67638 468888
rect 67694 468832 70226 468888
rect 67633 468830 70226 468832
rect 67633 468827 67699 468830
rect 70166 468724 70226 468830
rect 99790 468888 102199 468890
rect 99790 468832 102138 468888
rect 102194 468832 102199 468888
rect 99790 468830 102199 468832
rect 99790 468724 99850 468830
rect 102133 468827 102199 468830
rect 30281 468482 30347 468485
rect 64229 468482 64295 468485
rect 30281 468480 64295 468482
rect 30281 468424 30286 468480
rect 30342 468424 64234 468480
rect 64290 468424 64295 468480
rect 30281 468422 64295 468424
rect 30281 468419 30347 468422
rect 64229 468419 64295 468422
rect 67633 468210 67699 468213
rect 67633 468208 70226 468210
rect 67633 468152 67638 468208
rect 67694 468152 70226 468208
rect 67633 468150 70226 468152
rect 67633 468147 67699 468150
rect 70166 468044 70226 468150
rect 64086 467876 64092 467940
rect 64156 467938 64162 467940
rect 64229 467938 64295 467941
rect 64156 467936 64295 467938
rect 64156 467880 64234 467936
rect 64290 467880 64295 467936
rect 64156 467878 64295 467880
rect 64156 467876 64162 467878
rect 64229 467875 64295 467878
rect 107561 467938 107627 467941
rect 107694 467938 107700 467940
rect 107561 467936 107700 467938
rect 107561 467880 107566 467936
rect 107622 467880 107700 467936
rect 107561 467878 107700 467880
rect 107561 467875 107627 467878
rect 107694 467876 107700 467878
rect 107764 467876 107770 467940
rect 102133 467530 102199 467533
rect 99790 467528 102199 467530
rect 99790 467472 102138 467528
rect 102194 467472 102199 467528
rect 99790 467470 102199 467472
rect 99790 467364 99850 467470
rect 102133 467467 102199 467470
rect 102225 466986 102291 466989
rect 99790 466984 102291 466986
rect 99790 466928 102230 466984
rect 102286 466928 102291 466984
rect 99790 466926 102291 466928
rect 67449 466850 67515 466853
rect 67449 466848 70226 466850
rect 67449 466792 67454 466848
rect 67510 466792 70226 466848
rect 67449 466790 70226 466792
rect 67449 466787 67515 466790
rect 70166 466684 70226 466790
rect 99790 466684 99850 466926
rect 102225 466923 102291 466926
rect 67725 466170 67791 466173
rect 102225 466170 102291 466173
rect 67725 466168 70226 466170
rect 67725 466112 67730 466168
rect 67786 466112 70226 466168
rect 67725 466110 70226 466112
rect 67725 466107 67791 466110
rect 70166 466004 70226 466110
rect 99790 466168 102291 466170
rect 99790 466112 102230 466168
rect 102286 466112 102291 466168
rect 99790 466110 102291 466112
rect 99790 466004 99850 466110
rect 102225 466107 102291 466110
rect 67633 465626 67699 465629
rect 104065 465628 104131 465629
rect 104014 465626 104020 465628
rect 67633 465624 70226 465626
rect 67633 465568 67638 465624
rect 67694 465568 70226 465624
rect 67633 465566 70226 465568
rect 67633 465563 67699 465566
rect 70166 465324 70226 465566
rect 99606 465566 104020 465626
rect 104084 465624 104131 465628
rect 104126 465568 104131 465624
rect 99606 465324 99666 465566
rect 104014 465564 104020 465566
rect 104084 465564 104131 465568
rect 104065 465563 104131 465564
rect 102317 464946 102383 464949
rect 99790 464944 102383 464946
rect 99790 464888 102322 464944
rect 102378 464888 102383 464944
rect 99790 464886 102383 464888
rect 67633 464810 67699 464813
rect 67633 464808 70226 464810
rect 67633 464752 67638 464808
rect 67694 464752 70226 464808
rect 67633 464750 70226 464752
rect 67633 464747 67699 464750
rect 70166 464644 70226 464750
rect 99790 464644 99850 464886
rect 102317 464883 102383 464886
rect 67725 464266 67791 464269
rect 102133 464266 102199 464269
rect 67725 464264 70226 464266
rect 67725 464208 67730 464264
rect 67786 464208 70226 464264
rect 67725 464206 70226 464208
rect 67725 464203 67791 464206
rect 70166 463964 70226 464206
rect 99790 464264 102199 464266
rect 99790 464208 102138 464264
rect 102194 464208 102199 464264
rect 99790 464206 102199 464208
rect 99790 463964 99850 464206
rect 102133 464203 102199 464206
rect 58750 463524 58756 463588
rect 58820 463586 58826 463588
rect 61377 463586 61443 463589
rect 58820 463584 61443 463586
rect 58820 463528 61382 463584
rect 61438 463528 61443 463584
rect 58820 463526 61443 463528
rect 58820 463524 58826 463526
rect 61377 463523 61443 463526
rect 102133 463450 102199 463453
rect 99790 463448 102199 463450
rect 99790 463392 102138 463448
rect 102194 463392 102199 463448
rect 99790 463390 102199 463392
rect 99790 463284 99850 463390
rect 102133 463387 102199 463390
rect 67633 462770 67699 462773
rect 70166 462770 70226 463148
rect 67633 462768 70226 462770
rect -960 462634 480 462724
rect 67633 462712 67638 462768
rect 67694 462712 70226 462768
rect 67633 462710 70226 462712
rect 67633 462707 67699 462710
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 61377 462362 61443 462365
rect 61377 462360 69858 462362
rect 61377 462304 61382 462360
rect 61438 462304 69858 462360
rect 61377 462302 69858 462304
rect 61377 462299 61443 462302
rect 58985 462228 59051 462229
rect 58934 462226 58940 462228
rect 58894 462166 58940 462226
rect 59004 462224 59051 462228
rect 59046 462168 59051 462224
rect 58934 462164 58940 462166
rect 59004 462164 59051 462168
rect 69798 462226 69858 462302
rect 70350 462226 70410 462468
rect 69798 462166 70410 462226
rect 58985 462163 59051 462164
rect 102133 462090 102199 462093
rect 99790 462088 102199 462090
rect 99790 462032 102138 462088
rect 102194 462032 102199 462088
rect 99790 462030 102199 462032
rect 99790 461924 99850 462030
rect 102133 462027 102199 462030
rect 58934 461484 58940 461548
rect 59004 461546 59010 461548
rect 102225 461546 102291 461549
rect 59004 461486 70226 461546
rect 59004 461484 59010 461486
rect 70166 461244 70226 461486
rect 99790 461544 102291 461546
rect 99790 461488 102230 461544
rect 102286 461488 102291 461544
rect 99790 461486 102291 461488
rect 99790 461244 99850 461486
rect 102225 461483 102291 461486
rect 102133 460730 102199 460733
rect 99790 460728 102199 460730
rect 99790 460672 102138 460728
rect 102194 460672 102199 460728
rect 99790 460670 102199 460672
rect 99790 460564 99850 460670
rect 102133 460667 102199 460670
rect 67633 460186 67699 460189
rect 70350 460186 70410 460428
rect 67633 460184 70410 460186
rect 67633 460128 67638 460184
rect 67694 460128 70410 460184
rect 67633 460126 70410 460128
rect 67633 460123 67699 460126
rect 102133 460050 102199 460053
rect 67774 459990 70226 460050
rect 42609 459506 42675 459509
rect 67774 459506 67834 459990
rect 70166 459884 70226 459990
rect 99790 460048 102199 460050
rect 99790 459992 102138 460048
rect 102194 459992 102199 460048
rect 99790 459990 102199 459992
rect 99790 459884 99850 459990
rect 102133 459987 102199 459990
rect 118785 459644 118851 459645
rect 118734 459580 118740 459644
rect 118804 459642 118851 459644
rect 118804 459640 118896 459642
rect 118846 459584 118896 459640
rect 118804 459582 118896 459584
rect 118804 459580 118851 459582
rect 118785 459579 118851 459580
rect 42609 459504 67834 459506
rect 42609 459448 42614 459504
rect 42670 459448 67834 459504
rect 42609 459446 67834 459448
rect 42609 459443 42675 459446
rect 67725 459370 67791 459373
rect 102133 459370 102199 459373
rect 67725 459368 70226 459370
rect 67725 459312 67730 459368
rect 67786 459312 70226 459368
rect 67725 459310 70226 459312
rect 67725 459307 67791 459310
rect 70166 459204 70226 459310
rect 99790 459368 102199 459370
rect 99790 459312 102138 459368
rect 102194 459312 102199 459368
rect 99790 459310 102199 459312
rect 99790 459204 99850 459310
rect 102133 459307 102199 459310
rect 67633 458826 67699 458829
rect 102225 458826 102291 458829
rect 67633 458824 70410 458826
rect 67633 458768 67638 458824
rect 67694 458768 70410 458824
rect 67633 458766 70410 458768
rect 67633 458763 67699 458766
rect 70350 458524 70410 458766
rect 99790 458824 102291 458826
rect 99790 458768 102230 458824
rect 102286 458768 102291 458824
rect 99790 458766 102291 458768
rect 99790 458524 99850 458766
rect 102225 458763 102291 458766
rect 101305 458146 101371 458149
rect 99790 458144 101371 458146
rect 99790 458088 101310 458144
rect 101366 458088 101371 458144
rect 99790 458086 101371 458088
rect 99790 457844 99850 458086
rect 101305 458083 101371 458086
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 67633 457466 67699 457469
rect 70350 457466 70410 457708
rect 67633 457464 70410 457466
rect 67633 457408 67638 457464
rect 67694 457408 70410 457464
rect 67633 457406 70410 457408
rect 67633 457403 67699 457406
rect 67633 457330 67699 457333
rect 67633 457328 70226 457330
rect 67633 457272 67638 457328
rect 67694 457272 70226 457328
rect 67633 457270 70226 457272
rect 67633 457267 67699 457270
rect 70166 457164 70226 457270
rect 67725 456242 67791 456245
rect 67725 456240 70226 456242
rect 67725 456184 67730 456240
rect 67786 456184 70226 456240
rect 67725 456182 70226 456184
rect 67725 456179 67791 456182
rect 70166 455804 70226 456182
rect 99790 456106 99850 456348
rect 102869 456106 102935 456109
rect 99790 456104 102935 456106
rect 99790 456048 102874 456104
rect 102930 456048 102935 456104
rect 99790 456046 102935 456048
rect 102869 456043 102935 456046
rect 121545 456106 121611 456109
rect 122230 456106 122236 456108
rect 121545 456104 122236 456106
rect 121545 456048 121550 456104
rect 121606 456048 122236 456104
rect 121545 456046 122236 456048
rect 121545 456043 121611 456046
rect 122230 456044 122236 456046
rect 122300 456106 122306 456108
rect 132534 456106 132540 456108
rect 122300 456046 132540 456106
rect 122300 456044 122306 456046
rect 132534 456044 132540 456046
rect 132604 456044 132610 456108
rect 103605 455970 103671 455973
rect 99790 455968 103671 455970
rect 99790 455912 103610 455968
rect 103666 455912 103671 455968
rect 99790 455910 103671 455912
rect 99790 455804 99850 455910
rect 103605 455907 103671 455910
rect 102225 455426 102291 455429
rect 99790 455424 102291 455426
rect 99790 455368 102230 455424
rect 102286 455368 102291 455424
rect 99790 455366 102291 455368
rect 99790 455124 99850 455366
rect 102225 455363 102291 455366
rect 67633 454610 67699 454613
rect 70166 454610 70226 454988
rect 102133 454746 102199 454749
rect 67633 454608 70226 454610
rect 67633 454552 67638 454608
rect 67694 454552 70226 454608
rect 67633 454550 70226 454552
rect 99790 454744 102199 454746
rect 99790 454688 102138 454744
rect 102194 454688 102199 454744
rect 99790 454686 102199 454688
rect 67633 454547 67699 454550
rect 99790 454444 99850 454686
rect 102133 454683 102199 454686
rect 68001 454066 68067 454069
rect 70166 454066 70226 454308
rect 68001 454064 70226 454066
rect 68001 454008 68006 454064
rect 68062 454008 70226 454064
rect 68001 454006 70226 454008
rect 68001 454003 68067 454006
rect 68878 453932 68938 454006
rect 68870 453868 68876 453932
rect 68940 453868 68946 453932
rect 67357 453386 67423 453389
rect 70166 453386 70226 453628
rect 67357 453384 70226 453386
rect 67357 453328 67362 453384
rect 67418 453328 70226 453384
rect 67357 453326 70226 453328
rect 99790 453386 99850 453628
rect 102869 453386 102935 453389
rect 99790 453384 102935 453386
rect 99790 453328 102874 453384
rect 102930 453328 102935 453384
rect 99790 453326 102935 453328
rect 67357 453323 67423 453326
rect 102869 453323 102935 453326
rect 67633 453250 67699 453253
rect 102133 453250 102199 453253
rect 118785 453252 118851 453253
rect 118734 453250 118740 453252
rect 67633 453248 70226 453250
rect 67633 453192 67638 453248
rect 67694 453192 70226 453248
rect 67633 453190 70226 453192
rect 67633 453187 67699 453190
rect 70166 453084 70226 453190
rect 99790 453248 102199 453250
rect 99790 453192 102138 453248
rect 102194 453192 102199 453248
rect 99790 453190 102199 453192
rect 118658 453190 118740 453250
rect 118804 453250 118851 453252
rect 128854 453250 128860 453252
rect 118804 453248 128860 453250
rect 118846 453192 128860 453248
rect 99790 453084 99850 453190
rect 102133 453187 102199 453190
rect 118734 453188 118740 453190
rect 118804 453190 128860 453192
rect 118804 453188 118851 453190
rect 128854 453188 128860 453190
rect 128924 453188 128930 453252
rect 118785 453187 118851 453188
rect 67633 452570 67699 452573
rect 108849 452570 108915 452573
rect 112294 452570 112300 452572
rect 67633 452568 70226 452570
rect 67633 452512 67638 452568
rect 67694 452512 70226 452568
rect 67633 452510 70226 452512
rect 67633 452507 67699 452510
rect 70166 452404 70226 452510
rect 108849 452568 112300 452570
rect 108849 452512 108854 452568
rect 108910 452512 112300 452568
rect 108849 452510 112300 452512
rect 108849 452507 108915 452510
rect 112294 452508 112300 452510
rect 112364 452508 112370 452572
rect 99606 452026 99666 452268
rect 102317 452026 102383 452029
rect 99606 452024 102383 452026
rect 99606 451968 102322 452024
rect 102378 451968 102383 452024
rect 99606 451966 102383 451968
rect 102317 451963 102383 451966
rect 68737 451890 68803 451893
rect 68737 451888 70226 451890
rect 68737 451832 68742 451888
rect 68798 451832 70226 451888
rect 68737 451830 70226 451832
rect 68737 451827 68803 451830
rect 70166 451724 70226 451830
rect 101581 451210 101647 451213
rect 99790 451208 101647 451210
rect 99790 451152 101586 451208
rect 101642 451152 101647 451208
rect 99790 451150 101647 451152
rect 99790 451044 99850 451150
rect 101581 451147 101647 451150
rect 67633 450802 67699 450805
rect 67633 450800 70226 450802
rect 67633 450744 67638 450800
rect 67694 450744 70226 450800
rect 67633 450742 70226 450744
rect 67633 450739 67699 450742
rect 70166 450364 70226 450742
rect 102133 450666 102199 450669
rect 99790 450664 102199 450666
rect 99790 450608 102138 450664
rect 102194 450608 102199 450664
rect 99790 450606 102199 450608
rect 99790 450364 99850 450606
rect 102133 450603 102199 450606
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 67725 449170 67791 449173
rect 70166 449170 70226 449548
rect 99790 449306 99850 449548
rect 102869 449306 102935 449309
rect 99790 449304 102935 449306
rect 99790 449248 102874 449304
rect 102930 449248 102935 449304
rect 99790 449246 102935 449248
rect 102869 449243 102935 449246
rect 102133 449170 102199 449173
rect 67725 449168 70226 449170
rect 67725 449112 67730 449168
rect 67786 449112 70226 449168
rect 67725 449110 70226 449112
rect 99790 449168 102199 449170
rect 99790 449112 102138 449168
rect 102194 449112 102199 449168
rect 99790 449110 102199 449112
rect 67725 449107 67791 449110
rect 99790 449004 99850 449110
rect 102133 449107 102199 449110
rect 70166 448626 70226 448868
rect 67406 448566 70226 448626
rect 41137 448490 41203 448493
rect 67406 448490 67466 448566
rect 41137 448488 67466 448490
rect 41137 448432 41142 448488
rect 41198 448432 67466 448488
rect 41137 448430 67466 448432
rect 67633 448490 67699 448493
rect 102225 448490 102291 448493
rect 67633 448488 70226 448490
rect 67633 448432 67638 448488
rect 67694 448432 70226 448488
rect 67633 448430 70226 448432
rect 41137 448427 41203 448430
rect 67633 448427 67699 448430
rect 70166 448324 70226 448430
rect 99790 448488 102291 448490
rect 99790 448432 102230 448488
rect 102286 448432 102291 448488
rect 99790 448430 102291 448432
rect 99790 448324 99850 448430
rect 102225 448427 102291 448430
rect 102133 447946 102199 447949
rect 99790 447944 102199 447946
rect 99790 447888 102138 447944
rect 102194 447888 102199 447944
rect 99790 447886 102199 447888
rect 35617 447810 35683 447813
rect 41137 447810 41203 447813
rect 35617 447808 41203 447810
rect 35617 447752 35622 447808
rect 35678 447752 41142 447808
rect 41198 447752 41203 447808
rect 35617 447750 41203 447752
rect 35617 447747 35683 447750
rect 41137 447747 41203 447750
rect 99790 447644 99850 447886
rect 102133 447883 102199 447886
rect 61837 447268 61903 447269
rect 61837 447266 61884 447268
rect 61792 447264 61884 447266
rect 61792 447208 61842 447264
rect 61792 447206 61884 447208
rect 61837 447204 61884 447206
rect 61948 447204 61954 447268
rect 67633 447266 67699 447269
rect 70166 447266 70226 447508
rect 67633 447264 70226 447266
rect 67633 447208 67638 447264
rect 67694 447208 70226 447264
rect 67633 447206 70226 447208
rect 61837 447203 61903 447204
rect 67633 447203 67699 447206
rect 67633 446450 67699 446453
rect 70166 446450 70226 446828
rect 99465 446586 99531 446589
rect 99790 446586 99850 446828
rect 102593 446586 102659 446589
rect 99465 446584 102659 446586
rect 99465 446528 99470 446584
rect 99526 446528 102598 446584
rect 102654 446528 102659 446584
rect 99465 446526 102659 446528
rect 99465 446523 99531 446526
rect 102593 446523 102659 446526
rect 67633 446448 70226 446450
rect 67633 446392 67638 446448
rect 67694 446392 70226 446448
rect 67633 446390 70226 446392
rect 67633 446387 67699 446390
rect 61326 445980 61332 446044
rect 61396 446042 61402 446044
rect 63125 446042 63191 446045
rect 61396 446040 63191 446042
rect 61396 445984 63130 446040
rect 63186 445984 63191 446040
rect 61396 445982 63191 445984
rect 61396 445980 61402 445982
rect 63125 445979 63191 445982
rect 65374 445770 65380 445772
rect 64830 445710 65380 445770
rect 38377 445634 38443 445637
rect 64830 445634 64890 445710
rect 65374 445708 65380 445710
rect 65444 445770 65450 445772
rect 70166 445770 70226 446148
rect 102501 445770 102567 445773
rect 65444 445710 70226 445770
rect 99790 445768 102567 445770
rect 99790 445712 102506 445768
rect 102562 445712 102567 445768
rect 99790 445710 102567 445712
rect 65444 445708 65450 445710
rect 38377 445632 64890 445634
rect 38377 445576 38382 445632
rect 38438 445576 64890 445632
rect 99790 445604 99850 445710
rect 102501 445707 102567 445710
rect 38377 445574 64890 445576
rect 38377 445571 38443 445574
rect 68921 445498 68987 445501
rect 68921 445496 70226 445498
rect 68921 445440 68926 445496
rect 68982 445440 70226 445496
rect 68921 445438 70226 445440
rect 68921 445435 68987 445438
rect 70166 444924 70226 445438
rect 103237 445226 103303 445229
rect 99790 445224 103303 445226
rect 99790 445168 103242 445224
rect 103298 445168 103303 445224
rect 99790 445166 103303 445168
rect 99790 444924 99850 445166
rect 103237 445163 103303 445166
rect 583520 444668 584960 444908
rect 69982 444350 70226 444410
rect 68185 444274 68251 444277
rect 69982 444274 70042 444350
rect 68185 444272 70042 444274
rect 68185 444216 68190 444272
rect 68246 444216 70042 444272
rect 70166 444244 70226 444350
rect 68185 444214 70042 444216
rect 68185 444211 68251 444214
rect 99606 443869 99666 444108
rect 67633 443866 67699 443869
rect 67633 443864 70226 443866
rect 67633 443808 67638 443864
rect 67694 443808 70226 443864
rect 67633 443806 70226 443808
rect 99606 443864 99715 443869
rect 99606 443808 99654 443864
rect 99710 443808 99715 443864
rect 99606 443806 99715 443808
rect 67633 443803 67699 443806
rect 70166 443564 70226 443806
rect 99649 443803 99715 443806
rect 99741 443730 99807 443733
rect 102225 443730 102291 443733
rect 99660 443728 102291 443730
rect 99660 443672 99746 443728
rect 99802 443672 102230 443728
rect 102286 443672 102291 443728
rect 99660 443670 102291 443672
rect 99741 443667 99850 443670
rect 102225 443667 102291 443670
rect 99790 443564 99850 443667
rect 102869 443050 102935 443053
rect 99790 443048 102935 443050
rect 99790 442992 102874 443048
rect 102930 442992 102935 443048
rect 99790 442990 102935 442992
rect 99790 442884 99850 442990
rect 102869 442987 102935 442990
rect 69790 442642 69796 442644
rect 64830 442582 69796 442642
rect 51574 442444 51580 442508
rect 51644 442506 51650 442508
rect 64830 442506 64890 442582
rect 69790 442580 69796 442582
rect 69860 442580 69866 442644
rect 51644 442446 64890 442506
rect 67725 442506 67791 442509
rect 70166 442506 70226 442748
rect 67725 442504 70226 442506
rect 67725 442448 67730 442504
rect 67786 442448 70226 442504
rect 67725 442446 70226 442448
rect 51644 442444 51650 442446
rect 67725 442443 67791 442446
rect 99414 442444 99420 442508
rect 99484 442506 99490 442508
rect 113173 442506 113239 442509
rect 99484 442504 113239 442506
rect 99484 442448 113178 442504
rect 113234 442448 113239 442504
rect 99484 442446 113239 442448
rect 99484 442444 99490 442446
rect 113173 442443 113239 442446
rect 67633 442370 67699 442373
rect 99373 442370 99439 442373
rect 132861 442370 132927 442373
rect 67633 442368 70226 442370
rect 67633 442312 67638 442368
rect 67694 442312 70226 442368
rect 67633 442310 70226 442312
rect 67633 442307 67699 442310
rect 70166 442204 70226 442310
rect 99373 442368 132927 442370
rect 99373 442312 99378 442368
rect 99434 442312 132866 442368
rect 132922 442312 132927 442368
rect 99373 442310 132927 442312
rect 99373 442307 99439 442310
rect 132861 442307 132927 442310
rect 99790 441690 99850 442068
rect 102041 441690 102107 441693
rect 121678 441690 121684 441692
rect 99790 441688 121684 441690
rect 99790 441632 102046 441688
rect 102102 441632 121684 441688
rect 99790 441630 121684 441632
rect 102041 441627 102107 441630
rect 121678 441628 121684 441630
rect 121748 441628 121754 441692
rect 67633 441146 67699 441149
rect 70350 441146 70410 441388
rect 67633 441144 70410 441146
rect 67633 441088 67638 441144
rect 67694 441088 70410 441144
rect 67633 441086 70410 441088
rect 99465 441146 99531 441149
rect 99606 441146 99666 441388
rect 102593 441146 102659 441149
rect 99465 441144 102659 441146
rect 99465 441088 99470 441144
rect 99526 441088 102598 441144
rect 102654 441088 102659 441144
rect 99465 441086 102659 441088
rect 67633 441083 67699 441086
rect 99465 441083 99531 441086
rect 102593 441083 102659 441086
rect 67633 441010 67699 441013
rect 67633 441008 70226 441010
rect 67633 440952 67638 441008
rect 67694 440952 70226 441008
rect 67633 440950 70226 440952
rect 67633 440947 67699 440950
rect 70166 440844 70226 440950
rect 97717 439922 97783 439925
rect 99046 439922 99052 439924
rect 97717 439920 99052 439922
rect 97717 439864 97722 439920
rect 97778 439864 99052 439920
rect 97717 439862 99052 439864
rect 97717 439859 97783 439862
rect 99046 439860 99052 439862
rect 99116 439860 99122 439924
rect 99606 439786 99666 440028
rect 102041 439786 102107 439789
rect 99606 439784 102107 439786
rect 99606 439728 102046 439784
rect 102102 439728 102107 439784
rect 99606 439726 102107 439728
rect 102041 439723 102107 439726
rect 121545 439378 121611 439381
rect 121729 439378 121795 439381
rect 124254 439378 124260 439380
rect 121545 439376 124260 439378
rect 121545 439320 121550 439376
rect 121606 439320 121734 439376
rect 121790 439320 124260 439376
rect 121545 439318 124260 439320
rect 121545 439315 121611 439318
rect 121729 439315 121795 439318
rect 124254 439316 124260 439318
rect 124324 439316 124330 439380
rect 69197 439106 69263 439109
rect 71037 439106 71103 439109
rect 69197 439104 71103 439106
rect 69197 439048 69202 439104
rect 69258 439048 71042 439104
rect 71098 439048 71103 439104
rect 69197 439046 71103 439048
rect 69197 439043 69263 439046
rect 71037 439043 71103 439046
rect 54886 438908 54892 438972
rect 54956 438970 54962 438972
rect 84193 438970 84259 438973
rect 85481 438970 85547 438973
rect 54956 438968 85547 438970
rect 54956 438912 84198 438968
rect 84254 438912 85486 438968
rect 85542 438912 85547 438968
rect 54956 438910 85547 438912
rect 54956 438908 54962 438910
rect 84193 438907 84259 438910
rect 85481 438907 85547 438910
rect 50797 438834 50863 438837
rect 50981 438834 51047 438837
rect 71957 438834 72023 438837
rect 50797 438832 72023 438834
rect 50797 438776 50802 438832
rect 50858 438776 50986 438832
rect 51042 438776 71962 438832
rect 72018 438776 72023 438832
rect 50797 438774 72023 438776
rect 50797 438771 50863 438774
rect 50981 438771 51047 438774
rect 71957 438771 72023 438774
rect 92565 438698 92631 438701
rect 106774 438698 106780 438700
rect 92565 438696 106780 438698
rect 92565 438640 92570 438696
rect 92626 438640 106780 438696
rect 92565 438638 106780 438640
rect 92565 438635 92631 438638
rect 106774 438636 106780 438638
rect 106844 438636 106850 438700
rect 59118 438092 59124 438156
rect 59188 438154 59194 438156
rect 69054 438154 69060 438156
rect 59188 438094 69060 438154
rect 59188 438092 59194 438094
rect 69054 438092 69060 438094
rect 69124 438092 69130 438156
rect 98361 437882 98427 437885
rect 99281 437882 99347 437885
rect 98361 437880 99347 437882
rect 98361 437824 98366 437880
rect 98422 437824 99286 437880
rect 99342 437824 99347 437880
rect 98361 437822 99347 437824
rect 98361 437819 98427 437822
rect 99281 437819 99347 437822
rect 50838 437412 50844 437476
rect 50908 437474 50914 437476
rect 78857 437474 78923 437477
rect 79685 437474 79751 437477
rect 50908 437472 79751 437474
rect 50908 437416 78862 437472
rect 78918 437416 79690 437472
rect 79746 437416 79751 437472
rect 50908 437414 79751 437416
rect 50908 437412 50914 437414
rect 78857 437411 78923 437414
rect 79685 437411 79751 437414
rect 87597 437474 87663 437477
rect 118918 437474 118924 437476
rect 87597 437472 118924 437474
rect 87597 437416 87602 437472
rect 87658 437416 118924 437472
rect 87597 437414 118924 437416
rect 87597 437411 87663 437414
rect 118918 437412 118924 437414
rect 118988 437412 118994 437476
rect 70342 437276 70348 437340
rect 70412 437338 70418 437340
rect 77293 437338 77359 437341
rect 77753 437338 77819 437341
rect 70412 437336 77819 437338
rect 70412 437280 77298 437336
rect 77354 437280 77758 437336
rect 77814 437280 77819 437336
rect 70412 437278 77819 437280
rect 70412 437276 70418 437278
rect 77293 437275 77359 437278
rect 77753 437275 77819 437278
rect 86217 437338 86283 437341
rect 110638 437338 110644 437340
rect 86217 437336 110644 437338
rect 86217 437280 86222 437336
rect 86278 437280 110644 437336
rect 86217 437278 110644 437280
rect 86217 437275 86283 437278
rect 110638 437276 110644 437278
rect 110708 437276 110714 437340
rect -960 436508 480 436748
rect 55070 435916 55076 435980
rect 55140 435978 55146 435980
rect 84285 435978 84351 435981
rect 84837 435978 84903 435981
rect 55140 435976 84903 435978
rect 55140 435920 84290 435976
rect 84346 435920 84842 435976
rect 84898 435920 84903 435976
rect 55140 435918 84903 435920
rect 55140 435916 55146 435918
rect 84285 435915 84351 435918
rect 84837 435915 84903 435918
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3509 423602 3575 423605
rect -960 423600 3575 423602
rect -960 423544 3514 423600
rect 3570 423544 3575 423600
rect -960 423542 3575 423544
rect -960 423452 480 423542
rect 3509 423539 3575 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 99281 407826 99347 407829
rect 129774 407826 129780 407828
rect 99281 407824 129780 407826
rect 99281 407768 99286 407824
rect 99342 407768 129780 407824
rect 99281 407766 129780 407768
rect 99281 407763 99347 407766
rect 129774 407764 129780 407766
rect 129844 407764 129850 407828
rect 74625 407554 74691 407557
rect 75177 407554 75243 407557
rect 74625 407552 75243 407554
rect 74625 407496 74630 407552
rect 74686 407496 75182 407552
rect 75238 407496 75243 407552
rect 74625 407494 75243 407496
rect 74625 407491 74691 407494
rect 75177 407491 75243 407494
rect 75177 407146 75243 407149
rect 338246 407146 338252 407148
rect 75177 407144 338252 407146
rect 75177 407088 75182 407144
rect 75238 407088 338252 407144
rect 75177 407086 338252 407088
rect 75177 407083 75243 407086
rect 338246 407084 338252 407086
rect 338316 407084 338322 407148
rect 115841 406330 115907 406333
rect 331254 406330 331260 406332
rect 115841 406328 331260 406330
rect 115841 406272 115846 406328
rect 115902 406272 331260 406328
rect 115841 406270 331260 406272
rect 115841 406267 115907 406270
rect 331254 406268 331260 406270
rect 331324 406268 331330 406332
rect 71681 405786 71747 405789
rect 180006 405786 180012 405788
rect 71681 405784 180012 405786
rect 71681 405728 71686 405784
rect 71742 405728 180012 405784
rect 71681 405726 180012 405728
rect 71681 405723 71747 405726
rect 180006 405724 180012 405726
rect 180076 405724 180082 405788
rect 92381 404970 92447 404973
rect 127014 404970 127020 404972
rect 92381 404968 127020 404970
rect 92381 404912 92386 404968
rect 92442 404912 127020 404968
rect 92381 404910 127020 404912
rect 92381 404907 92447 404910
rect 127014 404908 127020 404910
rect 127084 404908 127090 404972
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 66161 404426 66227 404429
rect 342294 404426 342300 404428
rect 66161 404424 342300 404426
rect 66161 404368 66166 404424
rect 66222 404368 342300 404424
rect 66161 404366 342300 404368
rect 66161 404363 66227 404366
rect 342294 404364 342300 404366
rect 342364 404364 342370 404428
rect 48957 402250 49023 402253
rect 88241 402250 88307 402253
rect 120022 402250 120028 402252
rect 48957 402248 84210 402250
rect 48957 402192 48962 402248
rect 49018 402192 84210 402248
rect 48957 402190 84210 402192
rect 48957 402187 49023 402190
rect 64086 401644 64092 401708
rect 64156 401706 64162 401708
rect 64781 401706 64847 401709
rect 64156 401704 64847 401706
rect 64156 401648 64786 401704
rect 64842 401648 64847 401704
rect 64156 401646 64847 401648
rect 84150 401706 84210 402190
rect 88241 402248 120028 402250
rect 88241 402192 88246 402248
rect 88302 402192 120028 402248
rect 88241 402190 120028 402192
rect 88241 402187 88307 402190
rect 120022 402188 120028 402190
rect 120092 402188 120098 402252
rect 85665 401706 85731 401709
rect 339534 401706 339540 401708
rect 84150 401704 339540 401706
rect 84150 401648 85670 401704
rect 85726 401648 339540 401704
rect 84150 401646 339540 401648
rect 64156 401644 64162 401646
rect 64781 401643 64847 401646
rect 85665 401643 85731 401646
rect 339534 401644 339540 401646
rect 339604 401644 339610 401708
rect 98637 400890 98703 400893
rect 125726 400890 125732 400892
rect 98637 400888 125732 400890
rect 98637 400832 98642 400888
rect 98698 400832 125732 400888
rect 98637 400830 125732 400832
rect 98637 400827 98703 400830
rect 125726 400828 125732 400830
rect 125796 400828 125802 400892
rect 101121 400346 101187 400349
rect 101254 400346 101260 400348
rect 101121 400344 101260 400346
rect 101121 400288 101126 400344
rect 101182 400288 101260 400344
rect 101121 400286 101260 400288
rect 101121 400283 101187 400286
rect 101254 400284 101260 400286
rect 101324 400346 101330 400348
rect 155217 400346 155283 400349
rect 101324 400344 155283 400346
rect 101324 400288 155222 400344
rect 155278 400288 155283 400344
rect 101324 400286 155283 400288
rect 101324 400284 101330 400286
rect 155217 400283 155283 400286
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 97993 397490 98059 397493
rect 345054 397490 345060 397492
rect 97993 397488 345060 397490
rect 97993 397432 97998 397488
rect 98054 397432 345060 397488
rect 97993 397430 345060 397432
rect 97993 397427 98059 397430
rect 345054 397428 345060 397430
rect 345124 397428 345130 397492
rect 104014 396612 104020 396676
rect 104084 396674 104090 396676
rect 117589 396674 117655 396677
rect 104084 396672 117655 396674
rect 104084 396616 117594 396672
rect 117650 396616 117655 396672
rect 104084 396614 117655 396616
rect 104084 396612 104090 396614
rect 117589 396611 117655 396614
rect 105537 395450 105603 395453
rect 118734 395450 118740 395452
rect 105537 395448 118740 395450
rect 105537 395392 105542 395448
rect 105598 395392 118740 395448
rect 105537 395390 118740 395392
rect 105537 395387 105603 395390
rect 118734 395388 118740 395390
rect 118804 395388 118810 395452
rect 102225 395314 102291 395317
rect 108941 395314 109007 395317
rect 170254 395314 170260 395316
rect 102225 395312 170260 395314
rect 102225 395256 102230 395312
rect 102286 395256 108946 395312
rect 109002 395256 170260 395312
rect 102225 395254 170260 395256
rect 102225 395251 102291 395254
rect 108941 395251 109007 395254
rect 170254 395252 170260 395254
rect 170324 395252 170330 395316
rect 68686 394708 68692 394772
rect 68756 394770 68762 394772
rect 231853 394770 231919 394773
rect 68756 394768 231919 394770
rect 68756 394712 231858 394768
rect 231914 394712 231919 394768
rect 68756 394710 231919 394712
rect 68756 394708 68762 394710
rect 231853 394707 231919 394710
rect 57830 393892 57836 393956
rect 57900 393954 57906 393956
rect 82997 393954 83063 393957
rect 57900 393952 83063 393954
rect 57900 393896 83002 393952
rect 83058 393896 83063 393952
rect 57900 393894 83063 393896
rect 57900 393892 57906 393894
rect 82997 393891 83063 393894
rect 95141 393954 95207 393957
rect 118918 393954 118924 393956
rect 95141 393952 118924 393954
rect 95141 393896 95146 393952
rect 95202 393896 118924 393952
rect 95141 393894 118924 393896
rect 95141 393891 95207 393894
rect 118918 393892 118924 393894
rect 118988 393892 118994 393956
rect 112621 392594 112687 392597
rect 124397 392594 124463 392597
rect 112621 392592 124463 392594
rect 112621 392536 112626 392592
rect 112682 392536 124402 392592
rect 124458 392536 124463 392592
rect 112621 392534 124463 392536
rect 112621 392531 112687 392534
rect 124397 392531 124463 392534
rect 583520 391628 584960 391868
rect 103421 391234 103487 391237
rect 114502 391234 114508 391236
rect 103421 391232 114508 391234
rect 103421 391176 103426 391232
rect 103482 391176 114508 391232
rect 103421 391174 114508 391176
rect 103421 391171 103487 391174
rect 114502 391172 114508 391174
rect 114572 391172 114578 391236
rect 50286 390764 50292 390828
rect 50356 390826 50362 390828
rect 50981 390826 51047 390829
rect 50356 390824 51047 390826
rect 50356 390768 50986 390824
rect 51042 390768 51047 390824
rect 50356 390766 51047 390768
rect 50356 390764 50362 390766
rect 50981 390763 51047 390766
rect 111558 390764 111564 390828
rect 111628 390826 111634 390828
rect 113909 390826 113975 390829
rect 169017 390826 169083 390829
rect 111628 390824 169083 390826
rect 111628 390768 113914 390824
rect 113970 390768 169022 390824
rect 169078 390768 169083 390824
rect 111628 390766 169083 390768
rect 111628 390764 111634 390766
rect 113909 390763 113975 390766
rect 169017 390763 169083 390766
rect 84929 390690 84995 390693
rect 166206 390690 166212 390692
rect 84929 390688 166212 390690
rect 84929 390632 84934 390688
rect 84990 390632 166212 390688
rect 84929 390630 166212 390632
rect 84929 390627 84995 390630
rect 166206 390628 166212 390630
rect 166276 390628 166282 390692
rect 69606 389812 69612 389876
rect 69676 389874 69682 389876
rect 78857 389874 78923 389877
rect 69676 389872 78923 389874
rect 69676 389816 78862 389872
rect 78918 389816 78923 389872
rect 69676 389814 78923 389816
rect 69676 389812 69682 389814
rect 78857 389811 78923 389814
rect 61694 389268 61700 389332
rect 61764 389330 61770 389332
rect 253197 389330 253263 389333
rect 61764 389328 253263 389330
rect 61764 389272 253202 389328
rect 253258 389272 253263 389328
rect 61764 389270 253263 389272
rect 61764 389268 61770 389270
rect 253197 389267 253263 389270
rect 68870 389132 68876 389196
rect 68940 389194 68946 389196
rect 335537 389194 335603 389197
rect 68940 389192 335603 389194
rect 68940 389136 335542 389192
rect 335598 389136 335603 389192
rect 68940 389134 335603 389136
rect 68940 389132 68946 389134
rect 335537 389131 335603 389134
rect 100017 388378 100083 388381
rect 122046 388378 122052 388380
rect 100017 388376 122052 388378
rect 100017 388320 100022 388376
rect 100078 388320 122052 388376
rect 100017 388318 122052 388320
rect 100017 388315 100083 388318
rect 122046 388316 122052 388318
rect 122116 388378 122122 388380
rect 191230 388378 191236 388380
rect 122116 388318 191236 388378
rect 122116 388316 122122 388318
rect 191230 388316 191236 388318
rect 191300 388316 191306 388380
rect 53598 387908 53604 387972
rect 53668 387970 53674 387972
rect 53741 387970 53807 387973
rect 53668 387968 53807 387970
rect 53668 387912 53746 387968
rect 53802 387912 53807 387968
rect 53668 387910 53807 387912
rect 53668 387908 53674 387910
rect 53741 387907 53807 387910
rect 109677 387970 109743 387973
rect 177297 387970 177363 387973
rect 109677 387968 177363 387970
rect 109677 387912 109682 387968
rect 109738 387912 177302 387968
rect 177358 387912 177363 387968
rect 109677 387910 177363 387912
rect 109677 387907 109743 387910
rect 177297 387907 177363 387910
rect 121545 387834 121611 387837
rect 121862 387834 121868 387836
rect 121545 387832 121868 387834
rect 121545 387776 121550 387832
rect 121606 387776 121868 387832
rect 121545 387774 121868 387776
rect 121545 387771 121611 387774
rect 121862 387772 121868 387774
rect 121932 387772 121938 387836
rect 104157 387018 104223 387021
rect 122598 387018 122604 387020
rect 104157 387016 122604 387018
rect 104157 386960 104162 387016
rect 104218 386960 122604 387016
rect 104157 386958 122604 386960
rect 104157 386955 104223 386958
rect 122598 386956 122604 386958
rect 122668 386956 122674 387020
rect 70945 385658 71011 385661
rect 340822 385658 340828 385660
rect 70945 385656 340828 385658
rect 70166 385250 70226 385628
rect 70945 385600 70950 385656
rect 71006 385600 340828 385656
rect 70945 385598 340828 385600
rect 70945 385595 71011 385598
rect 340822 385596 340828 385598
rect 340892 385596 340898 385660
rect 177246 385250 177252 385252
rect 64830 385190 177252 385250
rect 61878 385052 61884 385116
rect 61948 385114 61954 385116
rect 64830 385114 64890 385190
rect 177246 385188 177252 385190
rect 177316 385188 177322 385252
rect 61948 385054 64890 385114
rect 61948 385052 61954 385054
rect 117497 384978 117563 384981
rect 118509 384978 118575 384981
rect 115828 384976 118575 384978
rect 67633 384842 67699 384845
rect 70166 384842 70226 384948
rect 115828 384920 117502 384976
rect 117558 384920 118514 384976
rect 118570 384920 118575 384976
rect 115828 384918 118575 384920
rect 117497 384915 117563 384918
rect 118509 384915 118575 384918
rect 67633 384840 70226 384842
rect 67633 384784 67638 384840
rect 67694 384784 70226 384840
rect 67633 384782 70226 384784
rect 67633 384779 67699 384782
rect -960 384284 480 384524
rect 118601 384298 118667 384301
rect 115828 384296 118667 384298
rect 115828 384240 118606 384296
rect 118662 384240 118667 384296
rect 115828 384238 118667 384240
rect 118601 384235 118667 384238
rect 118601 383618 118667 383621
rect 115828 383616 118667 383618
rect 68737 383482 68803 383485
rect 70166 383482 70226 383588
rect 115828 383560 118606 383616
rect 118662 383560 118667 383616
rect 115828 383558 118667 383560
rect 118601 383555 118667 383558
rect 68737 383480 70226 383482
rect 68737 383424 68742 383480
rect 68798 383424 70226 383480
rect 68737 383422 70226 383424
rect 68737 383419 68803 383422
rect 67633 382530 67699 382533
rect 70166 382530 70226 382908
rect 67633 382528 70226 382530
rect 67633 382472 67638 382528
rect 67694 382472 70226 382528
rect 67633 382470 70226 382472
rect 67633 382467 67699 382470
rect 118601 382258 118667 382261
rect 115828 382256 118667 382258
rect 70166 381578 70226 382228
rect 115828 382200 118606 382256
rect 118662 382200 118667 382256
rect 115828 382198 118667 382200
rect 118601 382195 118667 382198
rect 118601 381578 118667 381581
rect 64830 381518 70226 381578
rect 115828 381576 118667 381578
rect 115828 381520 118606 381576
rect 118662 381520 118667 381576
rect 115828 381518 118667 381520
rect 62982 380972 62988 381036
rect 63052 381034 63058 381036
rect 64830 381034 64890 381518
rect 118601 381515 118667 381518
rect 63052 380974 64890 381034
rect 63052 380972 63058 380974
rect 60590 380836 60596 380900
rect 60660 380898 60666 380900
rect 67633 380898 67699 380901
rect 116393 380898 116459 380901
rect 60660 380896 67699 380898
rect 60660 380840 67638 380896
rect 67694 380840 67699 380896
rect 115828 380896 116459 380898
rect 60660 380838 67699 380840
rect 60660 380836 60666 380838
rect 67633 380835 67699 380838
rect 67909 380762 67975 380765
rect 68686 380762 68692 380764
rect 67909 380760 68692 380762
rect 67909 380704 67914 380760
rect 67970 380704 68692 380760
rect 67909 380702 68692 380704
rect 67909 380699 67975 380702
rect 68686 380700 68692 380702
rect 68756 380762 68762 380764
rect 70166 380762 70226 380868
rect 115828 380840 116398 380896
rect 116454 380840 116459 380896
rect 115828 380838 116459 380840
rect 116393 380835 116459 380838
rect 68756 380702 70226 380762
rect 68756 380700 68762 380702
rect 67541 380354 67607 380357
rect 69105 380354 69171 380357
rect 67541 380352 70226 380354
rect 67541 380296 67546 380352
rect 67602 380296 69110 380352
rect 69166 380296 70226 380352
rect 67541 380294 70226 380296
rect 67541 380291 67607 380294
rect 69105 380291 69171 380294
rect 70166 380188 70226 380294
rect 67633 379946 67699 379949
rect 67633 379944 70226 379946
rect 67633 379888 67638 379944
rect 67694 379888 70226 379944
rect 67633 379886 70226 379888
rect 67633 379883 67699 379886
rect 59353 379538 59419 379541
rect 60590 379538 60596 379540
rect 59353 379536 60596 379538
rect 59353 379480 59358 379536
rect 59414 379480 60596 379536
rect 59353 379478 60596 379480
rect 59353 379475 59419 379478
rect 60590 379476 60596 379478
rect 60660 379476 60666 379540
rect 70166 379508 70226 379886
rect 117405 379538 117471 379541
rect 118325 379538 118391 379541
rect 115828 379536 118391 379538
rect 115828 379480 117410 379536
rect 117466 379480 118330 379536
rect 118386 379480 118391 379536
rect 115828 379478 118391 379480
rect 117405 379475 117471 379478
rect 118325 379475 118391 379478
rect 209037 379538 209103 379541
rect 349102 379538 349108 379540
rect 209037 379536 349108 379538
rect 209037 379480 209042 379536
rect 209098 379480 349108 379536
rect 209037 379478 349108 379480
rect 209037 379475 209103 379478
rect 349102 379476 349108 379478
rect 349172 379476 349178 379540
rect 118601 378858 118667 378861
rect 115828 378856 118667 378858
rect 115828 378800 118606 378856
rect 118662 378800 118667 378856
rect 115828 378798 118667 378800
rect 118601 378795 118667 378798
rect 123334 378660 123340 378724
rect 123404 378722 123410 378724
rect 124121 378722 124187 378725
rect 129917 378722 129983 378725
rect 123404 378720 129983 378722
rect 123404 378664 124126 378720
rect 124182 378664 129922 378720
rect 129978 378664 129983 378720
rect 123404 378662 129983 378664
rect 123404 378660 123410 378662
rect 124121 378659 124187 378662
rect 129917 378659 129983 378662
rect 69054 378524 69060 378588
rect 69124 378586 69130 378588
rect 115933 378586 115999 378589
rect 69124 378526 70226 378586
rect 69124 378524 69130 378526
rect 70166 378148 70226 378526
rect 115798 378584 115999 378586
rect 115798 378528 115938 378584
rect 115994 378528 115999 378584
rect 115798 378526 115999 378528
rect 115798 378178 115858 378526
rect 115933 378523 115999 378526
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 118049 378178 118115 378181
rect 115798 378176 118115 378178
rect 115798 378148 118054 378176
rect 115828 378120 118054 378148
rect 118110 378120 118115 378176
rect 115828 378118 118115 378120
rect 118049 378115 118115 378118
rect 115473 377500 115539 377501
rect 115422 377498 115428 377500
rect 67633 377090 67699 377093
rect 70166 377090 70226 377468
rect 115382 377438 115428 377498
rect 115492 377496 115539 377500
rect 115534 377440 115539 377496
rect 115422 377436 115428 377438
rect 115492 377436 115539 377440
rect 115473 377435 115539 377436
rect 67633 377088 70226 377090
rect 67633 377032 67638 377088
rect 67694 377032 70226 377088
rect 67633 377030 70226 377032
rect 67633 377027 67699 377030
rect 59118 376892 59124 376956
rect 59188 376954 59194 376956
rect 66110 376954 66116 376956
rect 59188 376894 66116 376954
rect 59188 376892 59194 376894
rect 66110 376892 66116 376894
rect 66180 376954 66186 376956
rect 66180 376894 70226 376954
rect 66180 376892 66186 376894
rect 70166 376788 70226 376894
rect 118233 376818 118299 376821
rect 115828 376816 118299 376818
rect 115828 376760 118238 376816
rect 118294 376760 118299 376816
rect 115828 376758 118299 376760
rect 118233 376755 118299 376758
rect 118601 376138 118667 376141
rect 115828 376136 118667 376138
rect 115828 376080 118606 376136
rect 118662 376080 118667 376136
rect 115828 376078 118667 376080
rect 118601 376075 118667 376078
rect 67633 375594 67699 375597
rect 67633 375592 70226 375594
rect 67633 375536 67638 375592
rect 67694 375536 70226 375592
rect 67633 375534 70226 375536
rect 67633 375531 67699 375534
rect 70166 375428 70226 375534
rect 118141 375458 118207 375461
rect 115828 375456 118207 375458
rect 115828 375400 118146 375456
rect 118202 375400 118207 375456
rect 115828 375398 118207 375400
rect 118141 375395 118207 375398
rect 67633 374642 67699 374645
rect 70166 374642 70226 374748
rect 67633 374640 70226 374642
rect 67633 374584 67638 374640
rect 67694 374584 70226 374640
rect 67633 374582 70226 374584
rect 115289 374642 115355 374645
rect 188286 374642 188292 374644
rect 115289 374640 188292 374642
rect 115289 374584 115294 374640
rect 115350 374584 188292 374640
rect 115289 374582 188292 374584
rect 67633 374579 67699 374582
rect 115289 374579 115355 374582
rect 67725 374506 67791 374509
rect 67725 374504 70226 374506
rect 67725 374448 67730 374504
rect 67786 374448 70226 374504
rect 67725 374446 70226 374448
rect 67725 374443 67791 374446
rect 70166 374068 70226 374446
rect 115430 374068 115490 374582
rect 188286 374580 188292 374582
rect 188356 374580 188362 374644
rect 118601 373418 118667 373421
rect 115828 373416 118667 373418
rect 115828 373360 118606 373416
rect 118662 373360 118667 373416
rect 115828 373358 118667 373360
rect 118601 373355 118667 373358
rect 67725 373282 67791 373285
rect 67725 373280 70226 373282
rect 67725 373224 67730 373280
rect 67786 373224 70226 373280
rect 67725 373222 70226 373224
rect 67725 373219 67791 373222
rect 70166 372708 70226 373222
rect 115473 373146 115539 373149
rect 115473 373144 115858 373146
rect 115473 373088 115478 373144
rect 115534 373088 115858 373144
rect 115473 373086 115858 373088
rect 115473 373083 115539 373086
rect 115798 372738 115858 373086
rect 117865 372738 117931 372741
rect 115798 372736 117931 372738
rect 115798 372708 117870 372736
rect 115828 372680 117870 372708
rect 117926 372680 117931 372736
rect 115828 372678 117931 372680
rect 117865 372675 117931 372678
rect 67633 372466 67699 372469
rect 67633 372464 70226 372466
rect 67633 372408 67638 372464
rect 67694 372408 70226 372464
rect 67633 372406 70226 372408
rect 67633 372403 67699 372406
rect 70166 372028 70226 372406
rect 115289 371922 115355 371925
rect 115289 371920 115858 371922
rect 115289 371864 115294 371920
rect 115350 371864 115858 371920
rect 115289 371862 115858 371864
rect 115289 371859 115355 371862
rect 67449 371786 67515 371789
rect 67449 371784 70226 371786
rect 67449 371728 67454 371784
rect 67510 371728 70226 371784
rect 67449 371726 70226 371728
rect 67449 371723 67515 371726
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect 70166 371348 70226 371726
rect 115798 371378 115858 371862
rect 117773 371378 117839 371381
rect 115798 371376 117839 371378
rect 115798 371348 117778 371376
rect -960 371318 3575 371320
rect 115828 371320 117778 371348
rect 117834 371320 117839 371376
rect 115828 371318 117839 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 117773 371315 117839 371318
rect 141049 371378 141115 371381
rect 143533 371378 143599 371381
rect 324262 371378 324268 371380
rect 141049 371376 324268 371378
rect 141049 371320 141054 371376
rect 141110 371320 143538 371376
rect 143594 371320 324268 371376
rect 141049 371318 324268 371320
rect 141049 371315 141115 371318
rect 143533 371315 143599 371318
rect 324262 371316 324268 371318
rect 324332 371316 324338 371380
rect 118601 370698 118667 370701
rect 115828 370696 118667 370698
rect 115828 370640 118606 370696
rect 118662 370640 118667 370696
rect 115828 370638 118667 370640
rect 118601 370635 118667 370638
rect 67633 370426 67699 370429
rect 67633 370424 70226 370426
rect 67633 370368 67638 370424
rect 67694 370368 70226 370424
rect 67633 370366 70226 370368
rect 67633 370363 67699 370366
rect 70166 369988 70226 370366
rect 116669 370018 116735 370021
rect 118601 370018 118667 370021
rect 115828 370016 118667 370018
rect 115828 369960 116674 370016
rect 116730 369960 118606 370016
rect 118662 369960 118667 370016
rect 115828 369958 118667 369960
rect 116669 369955 116735 369958
rect 118601 369955 118667 369958
rect 67633 369746 67699 369749
rect 67633 369744 70226 369746
rect 67633 369688 67638 369744
rect 67694 369688 70226 369744
rect 67633 369686 70226 369688
rect 67633 369683 67699 369686
rect 70166 369308 70226 369686
rect 118417 368658 118483 368661
rect 115828 368656 118483 368658
rect 67633 368522 67699 368525
rect 70166 368522 70226 368628
rect 115828 368600 118422 368656
rect 118478 368600 118483 368656
rect 115828 368598 118483 368600
rect 118417 368595 118483 368598
rect 67633 368520 70226 368522
rect 67633 368464 67638 368520
rect 67694 368464 70226 368520
rect 67633 368462 70226 368464
rect 67633 368459 67699 368462
rect 118601 367978 118667 367981
rect 115828 367976 118667 367978
rect 115828 367920 118606 367976
rect 118662 367920 118667 367976
rect 115828 367918 118667 367920
rect 118601 367915 118667 367918
rect 117773 367298 117839 367301
rect 115828 367296 117839 367298
rect 115828 367268 117778 367296
rect 60549 367162 60615 367165
rect 61878 367162 61884 367164
rect 60549 367160 61884 367162
rect 60549 367104 60554 367160
rect 60610 367104 61884 367160
rect 60549 367102 61884 367104
rect 60549 367099 60615 367102
rect 61878 367100 61884 367102
rect 61948 367162 61954 367164
rect 70166 367162 70226 367268
rect 115798 367240 117778 367268
rect 117834 367240 117839 367296
rect 115798 367238 117839 367240
rect 115798 367162 115858 367238
rect 117773 367235 117839 367238
rect 61948 367102 70226 367162
rect 115430 367102 115858 367162
rect 61948 367100 61954 367102
rect 60590 366964 60596 367028
rect 60660 367026 60666 367028
rect 61377 367026 61443 367029
rect 67633 367026 67699 367029
rect 115289 367026 115355 367029
rect 115430 367026 115490 367102
rect 60660 367024 64890 367026
rect 60660 366968 61382 367024
rect 61438 366968 64890 367024
rect 60660 366966 64890 366968
rect 60660 366964 60666 366966
rect 61377 366963 61443 366966
rect 64830 366346 64890 366966
rect 67633 367024 70226 367026
rect 67633 366968 67638 367024
rect 67694 366968 70226 367024
rect 67633 366966 70226 366968
rect 67633 366963 67699 366966
rect 70166 366588 70226 366966
rect 115289 367024 115490 367026
rect 115289 366968 115294 367024
rect 115350 366968 115490 367024
rect 115289 366966 115490 366968
rect 115289 366963 115355 366966
rect 64830 366286 70226 366346
rect 70166 365908 70226 366286
rect 118141 365938 118207 365941
rect 115828 365936 118207 365938
rect 115828 365880 118146 365936
rect 118202 365880 118207 365936
rect 115828 365878 118207 365880
rect 118141 365875 118207 365878
rect 206461 365802 206527 365805
rect 326654 365802 326660 365804
rect 206461 365800 326660 365802
rect 206461 365744 206466 365800
rect 206522 365744 326660 365800
rect 206461 365742 326660 365744
rect 206461 365739 206527 365742
rect 326654 365740 326660 365742
rect 326724 365740 326730 365804
rect 117313 365258 117379 365261
rect 115828 365256 117379 365258
rect 115828 365200 117318 365256
rect 117374 365200 117379 365256
rect 115828 365198 117379 365200
rect 117313 365195 117379 365198
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect 118049 364578 118115 364581
rect 115828 364576 118115 364578
rect 115828 364548 118054 364576
rect 58934 364380 58940 364444
rect 59004 364442 59010 364444
rect 64505 364442 64571 364445
rect 70166 364442 70226 364548
rect 59004 364440 70226 364442
rect 59004 364384 64510 364440
rect 64566 364384 70226 364440
rect 59004 364382 70226 364384
rect 115798 364520 118054 364548
rect 118110 364520 118115 364576
rect 115798 364518 118115 364520
rect 115798 364442 115858 364518
rect 118049 364515 118115 364518
rect 198590 364516 198596 364580
rect 198660 364578 198666 364580
rect 261845 364578 261911 364581
rect 198660 364576 261911 364578
rect 198660 364520 261850 364576
rect 261906 364520 261911 364576
rect 198660 364518 261911 364520
rect 198660 364516 198666 364518
rect 261845 364515 261911 364518
rect 247033 364442 247099 364445
rect 332542 364442 332548 364444
rect 115798 364382 115990 364442
rect 59004 364380 59010 364382
rect 64505 364379 64571 364382
rect 115930 364309 115990 364382
rect 247033 364440 332548 364442
rect 247033 364384 247038 364440
rect 247094 364384 332548 364440
rect 247033 364382 332548 364384
rect 247033 364379 247099 364382
rect 332542 364380 332548 364382
rect 332612 364380 332618 364444
rect 67633 364306 67699 364309
rect 67633 364304 70226 364306
rect 67633 364248 67638 364304
rect 67694 364248 70226 364304
rect 67633 364246 70226 364248
rect 115930 364304 115999 364309
rect 115930 364248 115938 364304
rect 115994 364248 115999 364304
rect 115930 364246 115999 364248
rect 67633 364243 67699 364246
rect 70166 363868 70226 364246
rect 115933 364243 115999 364246
rect 139301 363626 139367 363629
rect 184054 363626 184060 363628
rect 139301 363624 184060 363626
rect 139301 363568 139306 363624
rect 139362 363568 184060 363624
rect 139301 363566 184060 363568
rect 139301 363563 139367 363566
rect 184054 363564 184060 363566
rect 184124 363564 184130 363628
rect 69197 363354 69263 363357
rect 69197 363352 70226 363354
rect 69197 363296 69202 363352
rect 69258 363296 70226 363352
rect 69197 363294 70226 363296
rect 69197 363291 69263 363294
rect 70166 363188 70226 363294
rect 118141 363218 118207 363221
rect 115828 363216 118207 363218
rect 115828 363160 118146 363216
rect 118202 363160 118207 363216
rect 115828 363158 118207 363160
rect 118141 363155 118207 363158
rect 196566 363156 196572 363220
rect 196636 363218 196642 363220
rect 285029 363218 285095 363221
rect 334014 363218 334020 363220
rect 196636 363216 334020 363218
rect 196636 363160 285034 363216
rect 285090 363160 334020 363216
rect 196636 363158 334020 363160
rect 196636 363156 196642 363158
rect 285029 363155 285095 363158
rect 334014 363156 334020 363158
rect 334084 363156 334090 363220
rect 227713 363082 227779 363085
rect 328494 363082 328500 363084
rect 227713 363080 328500 363082
rect 227713 363024 227718 363080
rect 227774 363024 328500 363080
rect 227713 363022 328500 363024
rect 227713 363019 227779 363022
rect 328494 363020 328500 363022
rect 328564 363020 328570 363084
rect 67633 362674 67699 362677
rect 67633 362672 70226 362674
rect 67633 362616 67638 362672
rect 67694 362616 70226 362672
rect 67633 362614 70226 362616
rect 67633 362611 67699 362614
rect 70166 362508 70226 362614
rect 117957 362538 118023 362541
rect 115828 362536 118023 362538
rect 115828 362480 117962 362536
rect 118018 362480 118023 362536
rect 115828 362478 118023 362480
rect 117957 362475 118023 362478
rect 195094 362340 195100 362404
rect 195164 362402 195170 362404
rect 217961 362402 218027 362405
rect 195164 362400 218027 362402
rect 195164 362344 217966 362400
rect 218022 362344 218027 362400
rect 195164 362342 218027 362344
rect 195164 362340 195170 362342
rect 217961 362339 218027 362342
rect 199326 362204 199332 362268
rect 199396 362266 199402 362268
rect 223481 362266 223547 362269
rect 199396 362264 223547 362266
rect 199396 362208 223486 362264
rect 223542 362208 223547 362264
rect 199396 362206 223547 362208
rect 199396 362204 199402 362206
rect 223481 362203 223547 362206
rect 274725 361994 274791 361997
rect 359457 361994 359523 361997
rect 274725 361992 359523 361994
rect 274725 361936 274730 361992
rect 274786 361936 359462 361992
rect 359518 361936 359523 361992
rect 274725 361934 359523 361936
rect 274725 361931 274791 361934
rect 359457 361931 359523 361934
rect 117681 361858 117747 361861
rect 115828 361856 117747 361858
rect 115828 361800 117686 361856
rect 117742 361800 117747 361856
rect 115828 361798 117747 361800
rect 117681 361795 117747 361798
rect 300117 361858 300183 361861
rect 319897 361858 319963 361861
rect 300117 361856 319963 361858
rect 300117 361800 300122 361856
rect 300178 361800 319902 361856
rect 319958 361800 319963 361856
rect 300117 361798 319963 361800
rect 300117 361795 300183 361798
rect 319897 361795 319963 361798
rect 200614 361660 200620 361724
rect 200684 361722 200690 361724
rect 248965 361722 249031 361725
rect 249701 361722 249767 361725
rect 200684 361720 249767 361722
rect 200684 361664 248970 361720
rect 249026 361664 249706 361720
rect 249762 361664 249767 361720
rect 200684 361662 249767 361664
rect 200684 361660 200690 361662
rect 248965 361659 249031 361662
rect 249701 361659 249767 361662
rect 119705 361586 119771 361589
rect 121678 361586 121684 361588
rect 119705 361584 121684 361586
rect 119705 361528 119710 361584
rect 119766 361528 121684 361584
rect 119705 361526 121684 361528
rect 119705 361523 119771 361526
rect 121678 361524 121684 361526
rect 121748 361586 121754 361588
rect 274725 361586 274791 361589
rect 121748 361584 274791 361586
rect 121748 361528 274730 361584
rect 274786 361528 274791 361584
rect 121748 361526 274791 361528
rect 121748 361524 121754 361526
rect 274725 361523 274791 361526
rect 118601 361178 118667 361181
rect 115828 361176 118667 361178
rect 67633 360770 67699 360773
rect 70166 360770 70226 361148
rect 115828 361120 118606 361176
rect 118662 361120 118667 361176
rect 115828 361118 118667 361120
rect 118601 361115 118667 361118
rect 67633 360768 70226 360770
rect 67633 360712 67638 360768
rect 67694 360712 70226 360768
rect 67633 360710 70226 360712
rect 67633 360707 67699 360710
rect 293217 360498 293283 360501
rect 320214 360498 320220 360500
rect 293217 360496 320220 360498
rect 67725 360226 67791 360229
rect 70166 360226 70226 360468
rect 293217 360440 293222 360496
rect 293278 360440 320220 360496
rect 293217 360438 320220 360440
rect 293217 360435 293283 360438
rect 320214 360436 320220 360438
rect 320284 360436 320290 360500
rect 195237 360362 195303 360365
rect 353385 360362 353451 360365
rect 353937 360362 354003 360365
rect 195237 360360 354003 360362
rect 195237 360304 195242 360360
rect 195298 360304 353390 360360
rect 353446 360304 353942 360360
rect 353998 360304 354003 360360
rect 195237 360302 354003 360304
rect 195237 360299 195303 360302
rect 353385 360299 353451 360302
rect 353937 360299 354003 360302
rect 67725 360224 70226 360226
rect 67725 360168 67730 360224
rect 67786 360168 70226 360224
rect 67725 360166 70226 360168
rect 117957 360226 118023 360229
rect 118918 360226 118924 360228
rect 117957 360224 118924 360226
rect 117957 360168 117962 360224
rect 118018 360168 118924 360224
rect 117957 360166 118924 360168
rect 67725 360163 67791 360166
rect 117957 360163 118023 360166
rect 118918 360164 118924 360166
rect 118988 360164 118994 360228
rect 198181 360226 198247 360229
rect 291469 360226 291535 360229
rect 198181 360224 291535 360226
rect 198181 360168 198186 360224
rect 198242 360168 291474 360224
rect 291530 360168 291535 360224
rect 198181 360166 291535 360168
rect 198181 360163 198247 360166
rect 291469 360163 291535 360166
rect 304349 360226 304415 360229
rect 499573 360226 499639 360229
rect 304349 360224 499639 360226
rect 304349 360168 304354 360224
rect 304410 360168 499578 360224
rect 499634 360168 499639 360224
rect 304349 360166 499639 360168
rect 304349 360163 304415 360166
rect 499573 360163 499639 360166
rect 118601 359818 118667 359821
rect 115828 359816 118667 359818
rect 67633 359682 67699 359685
rect 70166 359682 70226 359788
rect 115828 359760 118606 359816
rect 118662 359760 118667 359816
rect 115828 359758 118667 359760
rect 118601 359755 118667 359758
rect 67633 359680 70226 359682
rect 67633 359624 67638 359680
rect 67694 359624 70226 359680
rect 67633 359622 70226 359624
rect 271646 359622 277410 359682
rect 67633 359619 67699 359622
rect 146477 359410 146543 359413
rect 173014 359410 173020 359412
rect 146477 359408 173020 359410
rect 146477 359352 146482 359408
rect 146538 359352 173020 359408
rect 146477 359350 173020 359352
rect 146477 359347 146543 359350
rect 173014 359348 173020 359350
rect 173084 359348 173090 359412
rect 173249 359410 173315 359413
rect 271646 359410 271706 359622
rect 271965 359546 272031 359549
rect 271965 359544 272074 359546
rect 271965 359488 271970 359544
rect 272026 359488 272074 359544
rect 271965 359483 272074 359488
rect 173249 359408 271706 359410
rect 173249 359352 173254 359408
rect 173310 359352 271706 359408
rect 173249 359350 271706 359352
rect 173249 359347 173315 359350
rect 134517 359274 134583 359277
rect 272014 359274 272074 359483
rect 277350 359410 277410 359622
rect 317045 359546 317111 359549
rect 354673 359546 354739 359549
rect 317045 359544 354739 359546
rect 317045 359488 317050 359544
rect 317106 359488 354678 359544
rect 354734 359488 354739 359544
rect 317045 359486 354739 359488
rect 317045 359483 317111 359486
rect 354673 359483 354739 359486
rect 321737 359410 321803 359413
rect 277350 359408 321803 359410
rect 277350 359352 321742 359408
rect 321798 359352 321803 359408
rect 277350 359350 321803 359352
rect 321737 359347 321803 359350
rect 134517 359272 272074 359274
rect 134517 359216 134522 359272
rect 134578 359216 272074 359272
rect 134517 359214 272074 359216
rect 134517 359211 134583 359214
rect 118141 359138 118207 359141
rect 321502 359138 321508 359140
rect 115828 359136 118207 359138
rect 115828 359080 118146 359136
rect 118202 359080 118207 359136
rect 115828 359078 118207 359080
rect 319884 359078 321508 359138
rect 118141 359075 118207 359078
rect 321502 359076 321508 359078
rect 321572 359138 321578 359140
rect 321645 359138 321711 359141
rect 321572 359136 321711 359138
rect 321572 359080 321650 359136
rect 321706 359080 321711 359136
rect 321572 359078 321711 359080
rect 321572 359076 321578 359078
rect 321645 359075 321711 359078
rect 198774 358804 198780 358868
rect 198844 358866 198850 358868
rect 199653 358866 199719 358869
rect 198844 358864 199719 358866
rect 198844 358808 199658 358864
rect 199714 358808 199719 358864
rect 198844 358806 199719 358808
rect 198844 358804 198850 358806
rect 199653 358803 199719 358806
rect 319345 358866 319411 358869
rect 320030 358866 320036 358868
rect 319345 358864 320036 358866
rect 319345 358808 319350 358864
rect 319406 358808 320036 358864
rect 319345 358806 320036 358808
rect 319345 358803 319411 358806
rect 320030 358804 320036 358806
rect 320100 358804 320106 358868
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect 118601 358458 118667 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect 115828 358456 118667 358458
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 67541 358186 67607 358189
rect 70166 358186 70226 358428
rect 115828 358400 118606 358456
rect 118662 358400 118667 358456
rect 115828 358398 118667 358400
rect 118601 358395 118667 358398
rect 198089 358322 198155 358325
rect 198089 358320 200100 358322
rect 198089 358264 198094 358320
rect 198150 358264 200100 358320
rect 198089 358262 200100 358264
rect 198089 358259 198155 358262
rect 67541 358184 70226 358186
rect 67541 358128 67546 358184
rect 67602 358128 70226 358184
rect 67541 358126 70226 358128
rect 67541 358123 67607 358126
rect 67633 358050 67699 358053
rect 67633 358048 70226 358050
rect 67633 357992 67638 358048
rect 67694 357992 70226 358048
rect 67633 357990 70226 357992
rect 67633 357987 67699 357990
rect 70166 357748 70226 357990
rect 117589 357098 117655 357101
rect 118601 357098 118667 357101
rect 115828 357096 118667 357098
rect 68001 356962 68067 356965
rect 68870 356962 68876 356964
rect 68001 356960 68876 356962
rect 68001 356904 68006 356960
rect 68062 356904 68876 356960
rect 68001 356902 68876 356904
rect 68001 356899 68067 356902
rect 68870 356900 68876 356902
rect 68940 356962 68946 356964
rect 70166 356962 70226 357068
rect 115828 357040 117594 357096
rect 117650 357040 118606 357096
rect 118662 357040 118667 357096
rect 115828 357038 118667 357040
rect 117589 357035 117655 357038
rect 118601 357035 118667 357038
rect 68940 356902 70226 356962
rect 68940 356900 68946 356902
rect 60457 356690 60523 356693
rect 69606 356690 69612 356692
rect 60457 356688 69612 356690
rect 60457 356632 60462 356688
rect 60518 356632 69612 356688
rect 60457 356630 69612 356632
rect 60457 356627 60523 356630
rect 69606 356628 69612 356630
rect 69676 356628 69682 356692
rect 319302 356421 319362 356932
rect 320030 356628 320036 356692
rect 320100 356690 320106 356692
rect 494094 356690 494100 356692
rect 320100 356630 494100 356690
rect 320100 356628 320106 356630
rect 494094 356628 494100 356630
rect 494164 356628 494170 356692
rect 118601 356418 118667 356421
rect 115828 356416 118667 356418
rect 115828 356360 118606 356416
rect 118662 356360 118667 356416
rect 115828 356358 118667 356360
rect 118601 356355 118667 356358
rect 198273 356418 198339 356421
rect 198273 356416 200100 356418
rect 198273 356360 198278 356416
rect 198334 356360 200100 356416
rect 198273 356358 200100 356360
rect 319302 356416 319411 356421
rect 319302 356360 319350 356416
rect 319406 356360 319411 356416
rect 319302 356358 319411 356360
rect 198273 356355 198339 356358
rect 319345 356355 319411 356358
rect 118509 355738 118575 355741
rect 115828 355736 118575 355738
rect 67725 355602 67791 355605
rect 70166 355602 70226 355708
rect 115828 355680 118514 355736
rect 118570 355680 118575 355736
rect 115828 355678 118575 355680
rect 118509 355675 118575 355678
rect 67725 355600 70226 355602
rect 67725 355544 67730 355600
rect 67786 355544 70226 355600
rect 67725 355542 70226 355544
rect 67725 355539 67791 355542
rect 67633 355194 67699 355197
rect 67633 355192 70226 355194
rect 67633 355136 67638 355192
rect 67694 355136 70226 355192
rect 67633 355134 70226 355136
rect 67633 355131 67699 355134
rect 70166 355028 70226 355134
rect 118601 354378 118667 354381
rect 322841 354378 322907 354381
rect 115828 354376 118667 354378
rect 67541 353834 67607 353837
rect 70166 353834 70226 354348
rect 115828 354320 118606 354376
rect 118662 354320 118667 354376
rect 115828 354318 118667 354320
rect 319884 354376 322907 354378
rect 319884 354320 322846 354376
rect 322902 354320 322907 354376
rect 319884 354318 322907 354320
rect 118601 354315 118667 354318
rect 322841 354315 322907 354318
rect 67541 353832 70226 353834
rect 67541 353776 67546 353832
rect 67602 353776 70226 353832
rect 67541 353774 70226 353776
rect 67541 353771 67607 353774
rect 117773 353698 117839 353701
rect 115828 353696 117839 353698
rect 115828 353640 117778 353696
rect 117834 353640 117839 353696
rect 115828 353638 117839 353640
rect 117773 353635 117839 353638
rect 197997 353698 198063 353701
rect 197997 353696 200100 353698
rect 197997 353640 198002 353696
rect 198058 353640 200100 353696
rect 197997 353638 200100 353640
rect 197997 353635 198063 353638
rect 133873 353428 133939 353429
rect 133822 353426 133828 353428
rect 133782 353366 133828 353426
rect 133892 353424 133939 353428
rect 133934 353368 133939 353424
rect 133822 353364 133828 353366
rect 133892 353364 133939 353368
rect 133873 353363 133939 353364
rect 324497 353426 324563 353429
rect 327022 353426 327028 353428
rect 324497 353424 327028 353426
rect 324497 353368 324502 353424
rect 324558 353368 327028 353424
rect 324497 353366 327028 353368
rect 324497 353363 324563 353366
rect 327022 353364 327028 353366
rect 327092 353364 327098 353428
rect 115841 353290 115907 353293
rect 115798 353288 115907 353290
rect 115798 353232 115846 353288
rect 115902 353232 115907 353288
rect 115798 353227 115907 353232
rect 68921 353154 68987 353157
rect 68921 353152 70226 353154
rect 68921 353096 68926 353152
rect 68982 353096 70226 353152
rect 68921 353094 70226 353096
rect 68921 353091 68987 353094
rect 70166 352988 70226 353094
rect 115798 352988 115858 353227
rect 30281 352610 30347 352613
rect 66662 352610 66668 352612
rect 30281 352608 66668 352610
rect 30281 352552 30286 352608
rect 30342 352552 66668 352608
rect 30281 352550 66668 352552
rect 30281 352547 30347 352550
rect 66662 352548 66668 352550
rect 66732 352610 66738 352612
rect 66732 352550 70226 352610
rect 66732 352548 66738 352550
rect 70166 352308 70226 352550
rect 321553 352202 321619 352205
rect 322197 352202 322263 352205
rect 319884 352200 322263 352202
rect 319884 352144 321558 352200
rect 321614 352144 322202 352200
rect 322258 352144 322263 352200
rect 319884 352142 322263 352144
rect 321553 352139 321619 352142
rect 322197 352139 322263 352142
rect 580257 351930 580323 351933
rect 583520 351930 584960 352020
rect 580257 351928 584960 351930
rect 580257 351872 580262 351928
rect 580318 351872 584960 351928
rect 580257 351870 584960 351872
rect 580257 351867 580323 351870
rect 67633 351794 67699 351797
rect 67633 351792 70226 351794
rect 67633 351736 67638 351792
rect 67694 351736 70226 351792
rect 583520 351780 584960 351870
rect 67633 351734 70226 351736
rect 67633 351731 67699 351734
rect 70166 351628 70226 351734
rect 117405 351658 117471 351661
rect 115828 351656 117471 351658
rect 115828 351600 117410 351656
rect 117466 351600 117471 351656
rect 115828 351598 117471 351600
rect 117405 351595 117471 351598
rect 198273 351522 198339 351525
rect 198273 351520 200100 351522
rect 198273 351464 198278 351520
rect 198334 351464 200100 351520
rect 198273 351462 200100 351464
rect 198273 351459 198339 351462
rect 145189 351114 145255 351117
rect 191046 351114 191052 351116
rect 145189 351112 191052 351114
rect 145189 351056 145194 351112
rect 145250 351056 191052 351112
rect 145189 351054 191052 351056
rect 145189 351051 145255 351054
rect 191046 351052 191052 351054
rect 191116 351052 191122 351116
rect 118601 350978 118667 350981
rect 115828 350976 118667 350978
rect 115828 350920 118606 350976
rect 118662 350920 118667 350976
rect 115828 350918 118667 350920
rect 118601 350915 118667 350918
rect 118601 350298 118667 350301
rect 115828 350296 118667 350298
rect 69657 349890 69723 349893
rect 70166 349890 70226 350268
rect 115828 350240 118606 350296
rect 118662 350240 118667 350296
rect 115828 350238 118667 350240
rect 118601 350235 118667 350238
rect 322657 350162 322723 350165
rect 319884 350160 322723 350162
rect 319884 350104 322662 350160
rect 322718 350104 322723 350160
rect 319884 350102 322723 350104
rect 322657 350099 322723 350102
rect 69657 349888 70226 349890
rect 69657 349832 69662 349888
rect 69718 349832 70226 349888
rect 69657 349830 70226 349832
rect 69657 349827 69723 349830
rect 178534 349692 178540 349756
rect 178604 349754 178610 349756
rect 198774 349754 198780 349756
rect 178604 349694 198780 349754
rect 178604 349692 178610 349694
rect 198774 349692 198780 349694
rect 198844 349692 198850 349756
rect 197353 349618 197419 349621
rect 197353 349616 200100 349618
rect 67633 349210 67699 349213
rect 70166 349210 70226 349588
rect 197353 349560 197358 349616
rect 197414 349560 200100 349616
rect 197353 349558 200100 349560
rect 197353 349555 197419 349558
rect 67633 349208 70226 349210
rect 67633 349152 67638 349208
rect 67694 349152 70226 349208
rect 67633 349150 70226 349152
rect 67633 349147 67699 349150
rect 67633 349074 67699 349077
rect 67633 349072 70226 349074
rect 67633 349016 67638 349072
rect 67694 349016 70226 349072
rect 67633 349014 70226 349016
rect 67633 349011 67699 349014
rect 70166 348908 70226 349014
rect 118601 348938 118667 348941
rect 115828 348936 118667 348938
rect 115828 348880 118606 348936
rect 118662 348880 118667 348936
rect 115828 348878 118667 348880
rect 118601 348875 118667 348878
rect 143441 348530 143507 348533
rect 186814 348530 186820 348532
rect 143441 348528 186820 348530
rect 143441 348472 143446 348528
rect 143502 348472 186820 348528
rect 143441 348470 186820 348472
rect 143441 348467 143507 348470
rect 186814 348468 186820 348470
rect 186884 348468 186890 348532
rect 146201 348394 146267 348397
rect 192334 348394 192340 348396
rect 146201 348392 192340 348394
rect 146201 348336 146206 348392
rect 146262 348336 192340 348392
rect 146201 348334 192340 348336
rect 146201 348331 146267 348334
rect 192334 348332 192340 348334
rect 192404 348332 192410 348396
rect 118509 348258 118575 348261
rect 115828 348256 118575 348258
rect 115828 348200 118514 348256
rect 118570 348200 118575 348256
rect 115828 348198 118575 348200
rect 118509 348195 118575 348198
rect 66161 347716 66227 347717
rect 66110 347714 66116 347716
rect 66070 347654 66116 347714
rect 66180 347712 66227 347716
rect 66222 347656 66227 347712
rect 66110 347652 66116 347654
rect 66180 347652 66227 347656
rect 66161 347651 66227 347652
rect 67633 347714 67699 347717
rect 117497 347714 117563 347717
rect 132585 347716 132651 347717
rect 118734 347714 118740 347716
rect 67633 347712 70226 347714
rect 67633 347656 67638 347712
rect 67694 347656 70226 347712
rect 67633 347654 70226 347656
rect 67633 347651 67699 347654
rect 70166 347548 70226 347654
rect 117497 347712 118740 347714
rect 117497 347656 117502 347712
rect 117558 347656 118740 347712
rect 117497 347654 118740 347656
rect 117497 347651 117563 347654
rect 118734 347652 118740 347654
rect 118804 347652 118810 347716
rect 132534 347714 132540 347716
rect 132494 347654 132540 347714
rect 132604 347712 132651 347716
rect 132646 347656 132651 347712
rect 132534 347652 132540 347654
rect 132604 347652 132651 347656
rect 132585 347651 132651 347652
rect 118601 347578 118667 347581
rect 115828 347576 118667 347578
rect 115828 347520 118606 347576
rect 118662 347520 118667 347576
rect 115828 347518 118667 347520
rect 118601 347515 118667 347518
rect 197353 347442 197419 347445
rect 321829 347442 321895 347445
rect 322289 347442 322355 347445
rect 197353 347440 200100 347442
rect 197353 347384 197358 347440
rect 197414 347384 200100 347440
rect 197353 347382 200100 347384
rect 319884 347440 322355 347442
rect 319884 347384 321834 347440
rect 321890 347384 322294 347440
rect 322350 347384 322355 347440
rect 319884 347382 322355 347384
rect 197353 347379 197419 347382
rect 321829 347379 321895 347382
rect 322289 347379 322355 347382
rect 65374 347244 65380 347308
rect 65444 347306 65450 347308
rect 68921 347306 68987 347309
rect 65444 347304 70226 347306
rect 65444 347248 68926 347304
rect 68982 347248 70226 347304
rect 65444 347246 70226 347248
rect 65444 347244 65450 347246
rect 68921 347243 68987 347246
rect 70166 346868 70226 347246
rect 68829 346354 68895 346357
rect 150525 346354 150591 346357
rect 200614 346354 200620 346356
rect 68829 346352 70226 346354
rect 68829 346296 68834 346352
rect 68890 346296 70226 346352
rect 68829 346294 70226 346296
rect 68829 346291 68895 346294
rect 70166 346188 70226 346294
rect 150525 346352 200620 346354
rect 150525 346296 150530 346352
rect 150586 346296 200620 346352
rect 150525 346294 200620 346296
rect 150525 346291 150591 346294
rect 200614 346292 200620 346294
rect 200684 346292 200690 346356
rect 118509 346218 118575 346221
rect 115828 346216 118575 346218
rect 115828 346160 118514 346216
rect 118570 346160 118575 346216
rect 115828 346158 118575 346160
rect 118509 346155 118575 346158
rect 140865 345674 140931 345677
rect 150525 345674 150591 345677
rect 140865 345672 150591 345674
rect 140865 345616 140870 345672
rect 140926 345616 150530 345672
rect 150586 345616 150591 345672
rect 140865 345614 150591 345616
rect 140865 345611 140931 345614
rect 150525 345611 150591 345614
rect 118601 345538 118667 345541
rect 320265 345538 320331 345541
rect 115828 345536 118667 345538
rect -960 345402 480 345492
rect 115828 345480 118606 345536
rect 118662 345480 118667 345536
rect 115828 345478 118667 345480
rect 319884 345536 320331 345538
rect 319884 345480 320270 345536
rect 320326 345480 320331 345536
rect 319884 345478 320331 345480
rect 118601 345475 118667 345478
rect 320265 345475 320331 345478
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 68645 344994 68711 344997
rect 68645 344992 70226 344994
rect 68645 344936 68650 344992
rect 68706 344936 70226 344992
rect 68645 344934 70226 344936
rect 68645 344931 68711 344934
rect 70166 344828 70226 344934
rect 118601 344858 118667 344861
rect 115828 344856 118667 344858
rect 115828 344800 118606 344856
rect 118662 344800 118667 344856
rect 115828 344798 118667 344800
rect 118601 344795 118667 344798
rect 198181 344722 198247 344725
rect 198181 344720 200100 344722
rect 198181 344664 198186 344720
rect 198242 344664 200100 344720
rect 198181 344662 200100 344664
rect 198181 344659 198247 344662
rect 67633 343770 67699 343773
rect 70166 343770 70226 344148
rect 67633 343768 70226 343770
rect 67633 343712 67638 343768
rect 67694 343712 70226 343768
rect 67633 343710 70226 343712
rect 67633 343707 67699 343710
rect 118601 343498 118667 343501
rect 115828 343496 118667 343498
rect 67633 342954 67699 342957
rect 70166 342954 70226 343468
rect 115828 343440 118606 343496
rect 118662 343440 118667 343496
rect 115828 343438 118667 343440
rect 118601 343435 118667 343438
rect 322473 343362 322539 343365
rect 319884 343360 322539 343362
rect 319884 343304 322478 343360
rect 322534 343304 322539 343360
rect 319884 343302 322539 343304
rect 322473 343299 322539 343302
rect 67633 342952 70226 342954
rect 67633 342896 67638 342952
rect 67694 342896 70226 342952
rect 67633 342894 70226 342896
rect 67633 342891 67699 342894
rect 117773 342818 117839 342821
rect 115828 342816 117839 342818
rect 115828 342760 117778 342816
rect 117834 342760 117839 342816
rect 115828 342758 117839 342760
rect 117773 342755 117839 342758
rect 197997 342682 198063 342685
rect 197997 342680 200100 342682
rect 197997 342624 198002 342680
rect 198058 342624 200100 342680
rect 197997 342622 200100 342624
rect 197997 342619 198063 342622
rect 128721 342274 128787 342277
rect 128854 342274 128860 342276
rect 128721 342272 128860 342274
rect 128721 342216 128726 342272
rect 128782 342216 128860 342272
rect 128721 342214 128860 342216
rect 128721 342211 128787 342214
rect 128854 342212 128860 342214
rect 128924 342274 128930 342276
rect 131757 342274 131823 342277
rect 128924 342272 131823 342274
rect 128924 342216 131762 342272
rect 131818 342216 131823 342272
rect 128924 342214 131823 342216
rect 128924 342212 128930 342214
rect 131757 342211 131823 342214
rect 117313 342138 117379 342141
rect 118509 342138 118575 342141
rect 115828 342136 118575 342138
rect 67909 341730 67975 341733
rect 68737 341730 68803 341733
rect 70166 341730 70226 342108
rect 115828 342080 117318 342136
rect 117374 342080 118514 342136
rect 118570 342080 118575 342136
rect 115828 342078 118575 342080
rect 117313 342075 117379 342078
rect 118509 342075 118575 342078
rect 67909 341728 70226 341730
rect 67909 341672 67914 341728
rect 67970 341672 68742 341728
rect 68798 341672 70226 341728
rect 67909 341670 70226 341672
rect 67909 341667 67975 341670
rect 68737 341667 68803 341670
rect 322841 341458 322907 341461
rect 319884 341456 322907 341458
rect 67633 341050 67699 341053
rect 70166 341050 70226 341428
rect 319884 341400 322846 341456
rect 322902 341400 322907 341456
rect 319884 341398 322907 341400
rect 322841 341395 322907 341398
rect 67633 341048 70226 341050
rect 67633 340992 67638 341048
rect 67694 340992 70226 341048
rect 67633 340990 70226 340992
rect 67633 340987 67699 340990
rect 117405 340778 117471 340781
rect 115828 340776 117471 340778
rect 67633 340234 67699 340237
rect 70166 340234 70226 340748
rect 115828 340720 117410 340776
rect 117466 340720 117471 340776
rect 115828 340718 117471 340720
rect 117405 340715 117471 340718
rect 197353 340642 197419 340645
rect 197353 340640 200100 340642
rect 197353 340584 197358 340640
rect 197414 340584 200100 340640
rect 197353 340582 200100 340584
rect 197353 340579 197419 340582
rect 67633 340232 70226 340234
rect 67633 340176 67638 340232
rect 67694 340176 70226 340232
rect 67633 340174 70226 340176
rect 67633 340171 67699 340174
rect 117313 340098 117379 340101
rect 115828 340096 117379 340098
rect 115828 340068 117318 340096
rect 115798 340040 117318 340068
rect 117374 340040 117379 340096
rect 115798 340038 117379 340040
rect 68921 339962 68987 339965
rect 75177 339962 75243 339965
rect 68921 339960 75243 339962
rect 68921 339904 68926 339960
rect 68982 339904 75182 339960
rect 75238 339904 75243 339960
rect 68921 339902 75243 339904
rect 68921 339899 68987 339902
rect 75177 339899 75243 339902
rect 115657 339826 115723 339829
rect 115798 339826 115858 340038
rect 117313 340035 117379 340038
rect 115657 339824 115858 339826
rect 115657 339768 115662 339824
rect 115718 339768 115858 339824
rect 115657 339766 115858 339768
rect 115657 339763 115723 339766
rect 111241 339690 111307 339693
rect 122598 339690 122604 339692
rect 111241 339688 122604 339690
rect 111241 339632 111246 339688
rect 111302 339632 122604 339688
rect 111241 339630 122604 339632
rect 111241 339627 111307 339630
rect 122598 339628 122604 339630
rect 122668 339628 122674 339692
rect 57789 339418 57855 339421
rect 79685 339418 79751 339421
rect 57789 339416 79751 339418
rect 57789 339360 57794 339416
rect 57850 339360 79690 339416
rect 79746 339360 79751 339416
rect 57789 339358 79751 339360
rect 57789 339355 57855 339358
rect 79685 339355 79751 339358
rect 84837 339418 84903 339421
rect 199326 339418 199332 339420
rect 84837 339416 199332 339418
rect 84837 339360 84842 339416
rect 84898 339360 199332 339416
rect 84837 339358 199332 339360
rect 84837 339355 84903 339358
rect 199326 339356 199332 339358
rect 199396 339356 199402 339420
rect 323025 338738 323091 338741
rect 319884 338736 323091 338738
rect 319884 338680 323030 338736
rect 323086 338680 323091 338736
rect 319884 338678 323091 338680
rect 323025 338675 323091 338678
rect 583520 338452 584960 338692
rect 115749 338058 115815 338061
rect 134149 338058 134215 338061
rect 135161 338058 135227 338061
rect 115749 338056 135227 338058
rect 115749 338000 115754 338056
rect 115810 338000 134154 338056
rect 134210 338000 135166 338056
rect 135222 338000 135227 338056
rect 115749 337998 135227 338000
rect 115749 337995 115815 337998
rect 134149 337995 134215 337998
rect 135161 337995 135227 337998
rect 117221 337922 117287 337925
rect 119705 337922 119771 337925
rect 117221 337920 119771 337922
rect 117221 337864 117226 337920
rect 117282 337864 119710 337920
rect 119766 337864 119771 337920
rect 117221 337862 119771 337864
rect 117221 337859 117287 337862
rect 119705 337859 119771 337862
rect 197353 337922 197419 337925
rect 197353 337920 200100 337922
rect 197353 337864 197358 337920
rect 197414 337864 200100 337920
rect 197353 337862 200100 337864
rect 197353 337859 197419 337862
rect 111793 337378 111859 337381
rect 129733 337378 129799 337381
rect 111793 337376 129799 337378
rect 111793 337320 111798 337376
rect 111854 337320 129738 337376
rect 129794 337320 129799 337376
rect 111793 337318 129799 337320
rect 111793 337315 111859 337318
rect 129733 337315 129799 337318
rect 135161 337378 135227 337381
rect 174537 337378 174603 337381
rect 135161 337376 174603 337378
rect 135161 337320 135166 337376
rect 135222 337320 174542 337376
rect 174598 337320 174603 337376
rect 135161 337318 174603 337320
rect 135161 337315 135227 337318
rect 174537 337315 174603 337318
rect 110229 336834 110295 336837
rect 117221 336834 117287 336837
rect 110229 336832 117287 336834
rect 110229 336776 110234 336832
rect 110290 336776 117226 336832
rect 117282 336776 117287 336832
rect 110229 336774 117287 336776
rect 110229 336771 110295 336774
rect 117221 336771 117287 336774
rect 322473 336698 322539 336701
rect 319884 336696 322539 336698
rect 319884 336640 322478 336696
rect 322534 336640 322539 336696
rect 319884 336638 322539 336640
rect 322473 336635 322539 336638
rect 77385 336018 77451 336021
rect 170397 336018 170463 336021
rect 77385 336016 170463 336018
rect 77385 335960 77390 336016
rect 77446 335960 170402 336016
rect 170458 335960 170463 336016
rect 77385 335958 170463 335960
rect 77385 335955 77451 335958
rect 170397 335955 170463 335958
rect 197353 335882 197419 335885
rect 197353 335880 200100 335882
rect 197353 335824 197358 335880
rect 197414 335824 200100 335880
rect 197353 335822 200100 335824
rect 197353 335819 197419 335822
rect 102041 335338 102107 335341
rect 125726 335338 125732 335340
rect 102041 335336 125732 335338
rect 102041 335280 102046 335336
rect 102102 335280 125732 335336
rect 102041 335278 125732 335280
rect 102041 335275 102107 335278
rect 125726 335276 125732 335278
rect 125796 335276 125802 335340
rect 103605 335202 103671 335205
rect 104801 335202 104867 335205
rect 120022 335202 120028 335204
rect 103605 335200 120028 335202
rect 103605 335144 103610 335200
rect 103666 335144 104806 335200
rect 104862 335144 120028 335200
rect 103605 335142 120028 335144
rect 103605 335139 103671 335142
rect 104801 335139 104867 335142
rect 120022 335140 120028 335142
rect 120092 335140 120098 335204
rect 321737 334658 321803 334661
rect 319884 334656 321803 334658
rect 319884 334600 321742 334656
rect 321798 334600 321803 334656
rect 319884 334598 321803 334600
rect 321737 334595 321803 334598
rect 95785 333978 95851 333981
rect 127014 333978 127020 333980
rect 95785 333976 127020 333978
rect 95785 333920 95790 333976
rect 95846 333920 127020 333976
rect 95785 333918 127020 333920
rect 95785 333915 95851 333918
rect 127014 333916 127020 333918
rect 127084 333916 127090 333980
rect 199009 333842 199075 333845
rect 199009 333840 200100 333842
rect 199009 333784 199014 333840
rect 199070 333784 200100 333840
rect 199009 333782 200100 333784
rect 199009 333779 199075 333782
rect 74625 333298 74691 333301
rect 195094 333298 195100 333300
rect 74625 333296 195100 333298
rect 74625 333240 74630 333296
rect 74686 333240 195100 333296
rect 74625 333238 195100 333240
rect 74625 333235 74691 333238
rect 195094 333236 195100 333238
rect 195164 333236 195170 333300
rect 95785 332618 95851 332621
rect 96521 332618 96587 332621
rect 95785 332616 96587 332618
rect 95785 332560 95790 332616
rect 95846 332560 96526 332616
rect 96582 332560 96587 332616
rect 95785 332558 96587 332560
rect 95785 332555 95851 332558
rect 96521 332555 96587 332558
rect -960 332196 480 332436
rect 197353 331802 197419 331805
rect 321645 331802 321711 331805
rect 322197 331802 322263 331805
rect 197353 331800 200100 331802
rect 197353 331744 197358 331800
rect 197414 331744 200100 331800
rect 197353 331742 200100 331744
rect 319884 331800 322263 331802
rect 319884 331744 321650 331800
rect 321706 331744 322202 331800
rect 322258 331744 322263 331800
rect 319884 331742 322263 331744
rect 197353 331739 197419 331742
rect 321645 331739 321711 331742
rect 322197 331739 322263 331742
rect 188521 331260 188587 331261
rect 69238 331196 69244 331260
rect 69308 331258 69314 331260
rect 188470 331258 188476 331260
rect 69308 331198 188476 331258
rect 188540 331256 188587 331260
rect 188582 331200 188587 331256
rect 69308 331196 69314 331198
rect 188470 331196 188476 331198
rect 188540 331196 188587 331200
rect 188521 331195 188587 331196
rect 322197 329898 322263 329901
rect 319884 329896 322263 329898
rect 319884 329840 322202 329896
rect 322258 329840 322263 329896
rect 319884 329838 322263 329840
rect 322197 329835 322263 329838
rect 197353 329082 197419 329085
rect 197353 329080 200100 329082
rect 197353 329024 197358 329080
rect 197414 329024 200100 329080
rect 197353 329022 200100 329024
rect 197353 329019 197419 329022
rect 107653 327722 107719 327725
rect 121862 327722 121868 327724
rect 107653 327720 121868 327722
rect 107653 327664 107658 327720
rect 107714 327664 121868 327720
rect 107653 327662 121868 327664
rect 107653 327659 107719 327662
rect 121862 327660 121868 327662
rect 121932 327660 121938 327724
rect 322841 327722 322907 327725
rect 319884 327720 322907 327722
rect 319884 327664 322846 327720
rect 322902 327664 322907 327720
rect 319884 327662 322907 327664
rect 322841 327659 322907 327662
rect 197353 327178 197419 327181
rect 197353 327176 200100 327178
rect 197353 327120 197358 327176
rect 197414 327120 200100 327176
rect 197353 327118 200100 327120
rect 197353 327115 197419 327118
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 198089 325002 198155 325005
rect 322749 325002 322815 325005
rect 198089 325000 200100 325002
rect 198089 324944 198094 325000
rect 198150 324944 200100 325000
rect 198089 324942 200100 324944
rect 319884 325000 322815 325002
rect 319884 324944 322754 325000
rect 322810 324944 322815 325000
rect 319884 324942 322815 324944
rect 198089 324939 198155 324942
rect 322749 324939 322815 324942
rect 322473 322962 322539 322965
rect 319884 322960 322539 322962
rect 319884 322904 322478 322960
rect 322534 322904 322539 322960
rect 319884 322902 322539 322904
rect 322473 322899 322539 322902
rect 197353 322418 197419 322421
rect 197353 322416 200100 322418
rect 197353 322360 197358 322416
rect 197414 322360 200100 322416
rect 197353 322358 200100 322360
rect 197353 322355 197419 322358
rect 322197 320922 322263 320925
rect 319884 320920 322263 320922
rect 319884 320864 322202 320920
rect 322258 320864 322263 320920
rect 319884 320862 322263 320864
rect 322197 320859 322263 320862
rect 69054 320724 69060 320788
rect 69124 320786 69130 320788
rect 69124 320726 122850 320786
rect 69124 320724 69130 320726
rect 122790 320242 122850 320726
rect 132493 320242 132559 320245
rect 172421 320242 172487 320245
rect 122790 320240 172487 320242
rect 122790 320184 132498 320240
rect 132554 320184 172426 320240
rect 172482 320184 172487 320240
rect 122790 320182 172487 320184
rect 132493 320179 132559 320182
rect 172421 320179 172487 320182
rect 197353 320242 197419 320245
rect 197353 320240 200100 320242
rect 197353 320184 197358 320240
rect 197414 320184 200100 320240
rect 197353 320182 200100 320184
rect 197353 320179 197419 320182
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 322841 318882 322907 318885
rect 319884 318880 322907 318882
rect 319884 318824 322846 318880
rect 322902 318824 322907 318880
rect 319884 318822 322907 318824
rect 322841 318819 322907 318822
rect 198641 318202 198707 318205
rect 198641 318200 200100 318202
rect 198641 318144 198646 318200
rect 198702 318144 200100 318200
rect 198641 318142 200100 318144
rect 198641 318139 198707 318142
rect 116669 318066 116735 318069
rect 129917 318066 129983 318069
rect 160686 318066 160692 318068
rect 116669 318064 160692 318066
rect 116669 318008 116674 318064
rect 116730 318008 129922 318064
rect 129978 318008 160692 318064
rect 116669 318006 160692 318008
rect 116669 318003 116735 318006
rect 129917 318003 129983 318006
rect 160686 318004 160692 318006
rect 160756 318004 160762 318068
rect 129774 317324 129780 317388
rect 129844 317386 129850 317388
rect 129917 317386 129983 317389
rect 129844 317384 129983 317386
rect 129844 317328 129922 317384
rect 129978 317328 129983 317384
rect 129844 317326 129983 317328
rect 129844 317324 129850 317326
rect 129917 317323 129983 317326
rect 322473 316298 322539 316301
rect 319884 316296 322539 316298
rect 319884 316240 322478 316296
rect 322534 316240 322539 316296
rect 319884 316238 322539 316240
rect 322473 316235 322539 316238
rect 129774 316100 129780 316164
rect 129844 316162 129850 316164
rect 130285 316162 130351 316165
rect 129844 316160 130351 316162
rect 129844 316104 130290 316160
rect 130346 316104 130351 316160
rect 129844 316102 130351 316104
rect 129844 316100 129850 316102
rect 130285 316099 130351 316102
rect 197353 315482 197419 315485
rect 197353 315480 200100 315482
rect 197353 315424 197358 315480
rect 197414 315424 200100 315480
rect 197353 315422 200100 315424
rect 197353 315419 197419 315422
rect 76649 315346 76715 315349
rect 193806 315346 193812 315348
rect 76649 315344 193812 315346
rect 76649 315288 76654 315344
rect 76710 315288 193812 315344
rect 76649 315286 193812 315288
rect 76649 315283 76715 315286
rect 193806 315284 193812 315286
rect 193876 315284 193882 315348
rect 124305 314668 124371 314669
rect 124254 314666 124260 314668
rect 124214 314606 124260 314666
rect 124324 314664 124371 314668
rect 124366 314608 124371 314664
rect 124254 314604 124260 314606
rect 124324 314604 124371 314608
rect 124305 314603 124371 314604
rect 322473 314258 322539 314261
rect 319884 314256 322539 314258
rect 319884 314200 322478 314256
rect 322534 314200 322539 314256
rect 319884 314198 322539 314200
rect 322473 314195 322539 314198
rect 197353 313442 197419 313445
rect 198917 313442 198983 313445
rect 197353 313440 200100 313442
rect 197353 313384 197358 313440
rect 197414 313384 198922 313440
rect 198978 313384 200100 313440
rect 197353 313382 200100 313384
rect 197353 313379 197419 313382
rect 198917 313379 198983 313382
rect 322841 312082 322907 312085
rect 319884 312080 322907 312082
rect 319884 312024 322846 312080
rect 322902 312024 322907 312080
rect 319884 312022 322907 312024
rect 322841 312019 322907 312022
rect 580349 312082 580415 312085
rect 583520 312082 584960 312172
rect 580349 312080 584960 312082
rect 580349 312024 580354 312080
rect 580410 312024 584960 312080
rect 580349 312022 584960 312024
rect 580349 312019 580415 312022
rect 583520 311932 584960 312022
rect 324262 311748 324268 311812
rect 324332 311810 324338 311812
rect 324405 311810 324471 311813
rect 324332 311808 324471 311810
rect 324332 311752 324410 311808
rect 324466 311752 324471 311808
rect 324332 311750 324471 311752
rect 324332 311748 324338 311750
rect 324405 311747 324471 311750
rect 197353 311402 197419 311405
rect 197353 311400 200100 311402
rect 197353 311344 197358 311400
rect 197414 311344 200100 311400
rect 197353 311342 200100 311344
rect 197353 311339 197419 311342
rect 98729 311130 98795 311133
rect 152406 311130 152412 311132
rect 98729 311128 152412 311130
rect 98729 311072 98734 311128
rect 98790 311072 152412 311128
rect 98729 311070 152412 311072
rect 98729 311067 98795 311070
rect 152406 311068 152412 311070
rect 152476 311068 152482 311132
rect 322473 309498 322539 309501
rect 319884 309496 322539 309498
rect 319884 309440 322478 309496
rect 322534 309440 322539 309496
rect 319884 309438 322539 309440
rect 322473 309435 322539 309438
rect 196801 309362 196867 309365
rect 196801 309360 200100 309362
rect 196801 309304 196806 309360
rect 196862 309304 200100 309360
rect 196801 309302 200100 309304
rect 196801 309299 196867 309302
rect 56225 308410 56291 308413
rect 125726 308410 125732 308412
rect 56225 308408 125732 308410
rect 56225 308352 56230 308408
rect 56286 308352 125732 308408
rect 56225 308350 125732 308352
rect 56225 308347 56291 308350
rect 125726 308348 125732 308350
rect 125796 308348 125802 308412
rect 322473 307458 322539 307461
rect 319884 307456 322539 307458
rect 319884 307400 322478 307456
rect 322534 307400 322539 307456
rect 319884 307398 322539 307400
rect 322473 307395 322539 307398
rect 197261 306642 197327 306645
rect 197261 306640 200100 306642
rect 197261 306584 197266 306640
rect 197322 306584 200100 306640
rect 197261 306582 200100 306584
rect 197261 306579 197327 306582
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 88977 305690 89043 305693
rect 195094 305690 195100 305692
rect 88977 305688 195100 305690
rect 88977 305632 88982 305688
rect 89038 305632 195100 305688
rect 88977 305630 195100 305632
rect 88977 305627 89043 305630
rect 195094 305628 195100 305630
rect 195164 305628 195170 305692
rect 322473 305282 322539 305285
rect 319884 305280 322539 305282
rect 319884 305224 322478 305280
rect 322534 305224 322539 305280
rect 319884 305222 322539 305224
rect 322473 305219 322539 305222
rect 197353 304602 197419 304605
rect 197353 304600 200100 304602
rect 197353 304544 197358 304600
rect 197414 304544 200100 304600
rect 197353 304542 200100 304544
rect 197353 304539 197419 304542
rect 322473 303242 322539 303245
rect 319884 303240 322539 303242
rect 319884 303184 322478 303240
rect 322534 303184 322539 303240
rect 319884 303182 322539 303184
rect 322473 303179 322539 303182
rect 97809 302834 97875 302837
rect 144126 302834 144132 302836
rect 97809 302832 144132 302834
rect 97809 302776 97814 302832
rect 97870 302776 144132 302832
rect 97809 302774 144132 302776
rect 97809 302771 97875 302774
rect 144126 302772 144132 302774
rect 144196 302772 144202 302836
rect 197353 302562 197419 302565
rect 197353 302560 200100 302562
rect 197353 302504 197358 302560
rect 197414 302504 200100 302560
rect 197353 302502 200100 302504
rect 197353 302499 197419 302502
rect 197445 301338 197511 301341
rect 197997 301338 198063 301341
rect 197445 301336 198063 301338
rect 197445 301280 197450 301336
rect 197506 301280 198002 301336
rect 198058 301280 198063 301336
rect 197445 301278 198063 301280
rect 197445 301275 197511 301278
rect 197997 301275 198063 301278
rect 70894 300868 70900 300932
rect 70964 300930 70970 300932
rect 197445 300930 197511 300933
rect 70964 300928 197511 300930
rect 70964 300872 197450 300928
rect 197506 300872 197511 300928
rect 70964 300870 197511 300872
rect 70964 300868 70970 300870
rect 197445 300867 197511 300870
rect 322841 300658 322907 300661
rect 319884 300656 322907 300658
rect 319884 300600 322846 300656
rect 322902 300600 322907 300656
rect 319884 300598 322907 300600
rect 322841 300595 322907 300598
rect 53557 300114 53623 300117
rect 138013 300114 138079 300117
rect 53557 300112 138079 300114
rect 53557 300056 53562 300112
rect 53618 300056 138018 300112
rect 138074 300056 138079 300112
rect 53557 300054 138079 300056
rect 53557 300051 53623 300054
rect 138013 300051 138079 300054
rect 197353 299978 197419 299981
rect 197353 299976 200100 299978
rect 197353 299920 197358 299976
rect 197414 299920 200100 299976
rect 197353 299918 200100 299920
rect 197353 299915 197419 299918
rect 49601 298890 49667 298893
rect 67449 298890 67515 298893
rect 49601 298888 67515 298890
rect 49601 298832 49606 298888
rect 49662 298832 67454 298888
rect 67510 298832 67515 298888
rect 49601 298830 67515 298832
rect 49601 298827 49667 298830
rect 67449 298827 67515 298830
rect 53598 298692 53604 298756
rect 53668 298754 53674 298756
rect 91277 298754 91343 298757
rect 53668 298752 91343 298754
rect 53668 298696 91282 298752
rect 91338 298696 91343 298752
rect 53668 298694 91343 298696
rect 53668 298692 53674 298694
rect 91277 298691 91343 298694
rect 580257 298754 580323 298757
rect 583520 298754 584960 298844
rect 580257 298752 584960 298754
rect 580257 298696 580262 298752
rect 580318 298696 584960 298752
rect 580257 298694 584960 298696
rect 580257 298691 580323 298694
rect 322473 298618 322539 298621
rect 319884 298616 322539 298618
rect 319884 298560 322478 298616
rect 322534 298560 322539 298616
rect 583520 298604 584960 298694
rect 319884 298558 322539 298560
rect 322473 298555 322539 298558
rect 67449 298346 67515 298349
rect 69013 298346 69079 298349
rect 67449 298344 69079 298346
rect 67449 298288 67454 298344
rect 67510 298288 69018 298344
rect 69074 298288 69079 298344
rect 67449 298286 69079 298288
rect 67449 298283 67515 298286
rect 69013 298283 69079 298286
rect 91277 298210 91343 298213
rect 162301 298210 162367 298213
rect 91277 298208 162367 298210
rect 91277 298152 91282 298208
rect 91338 298152 162306 298208
rect 162362 298152 162367 298208
rect 91277 298150 162367 298152
rect 91277 298147 91343 298150
rect 162301 298147 162367 298150
rect 197353 297802 197419 297805
rect 197353 297800 200100 297802
rect 197353 297744 197358 297800
rect 197414 297744 200100 297800
rect 197353 297742 200100 297744
rect 197353 297739 197419 297742
rect 102041 297394 102107 297397
rect 127617 297394 127683 297397
rect 102041 297392 127683 297394
rect 102041 297336 102046 297392
rect 102102 297336 127622 297392
rect 127678 297336 127683 297392
rect 102041 297334 127683 297336
rect 102041 297331 102107 297334
rect 127617 297331 127683 297334
rect 322473 296442 322539 296445
rect 319884 296440 322539 296442
rect 319884 296384 322478 296440
rect 322534 296384 322539 296440
rect 319884 296382 322539 296384
rect 322473 296379 322539 296382
rect 96521 296034 96587 296037
rect 141417 296034 141483 296037
rect 96521 296032 141483 296034
rect 96521 295976 96526 296032
rect 96582 295976 141422 296032
rect 141478 295976 141483 296032
rect 96521 295974 141483 295976
rect 96521 295971 96587 295974
rect 141417 295971 141483 295974
rect 197445 295762 197511 295765
rect 197445 295760 200100 295762
rect 197445 295704 197450 295760
rect 197506 295704 200100 295760
rect 197445 295702 200100 295704
rect 197445 295699 197511 295702
rect 118969 295218 119035 295221
rect 123569 295218 123635 295221
rect 118969 295216 123635 295218
rect 118969 295160 118974 295216
rect 119030 295160 123574 295216
rect 123630 295160 123635 295216
rect 118969 295158 123635 295160
rect 118969 295155 119035 295158
rect 123569 295155 123635 295158
rect 88701 294810 88767 294813
rect 119337 294810 119403 294813
rect 88701 294808 119403 294810
rect 88701 294752 88706 294808
rect 88762 294752 119342 294808
rect 119398 294752 119403 294808
rect 88701 294750 119403 294752
rect 88701 294747 88767 294750
rect 119337 294747 119403 294750
rect 81617 294674 81683 294677
rect 119521 294674 119587 294677
rect 81617 294672 119587 294674
rect 81617 294616 81622 294672
rect 81678 294616 119526 294672
rect 119582 294616 119587 294672
rect 81617 294614 119587 294616
rect 81617 294611 81683 294614
rect 119521 294611 119587 294614
rect 73245 294538 73311 294541
rect 80697 294538 80763 294541
rect 73245 294536 80763 294538
rect 73245 294480 73250 294536
rect 73306 294480 80702 294536
rect 80758 294480 80763 294536
rect 73245 294478 80763 294480
rect 73245 294475 73311 294478
rect 80697 294475 80763 294478
rect 104157 294538 104223 294541
rect 196566 294538 196572 294540
rect 104157 294536 196572 294538
rect 104157 294480 104162 294536
rect 104218 294480 196572 294536
rect 104157 294478 196572 294480
rect 104157 294475 104223 294478
rect 196566 294476 196572 294478
rect 196636 294476 196642 294540
rect 197445 293722 197511 293725
rect 322841 293722 322907 293725
rect 197445 293720 200100 293722
rect 197445 293664 197450 293720
rect 197506 293664 200100 293720
rect 197445 293662 200100 293664
rect 319884 293720 322907 293722
rect 319884 293664 322846 293720
rect 322902 293664 322907 293720
rect 319884 293662 322907 293664
rect 197445 293659 197511 293662
rect 322841 293659 322907 293662
rect 117129 293314 117195 293317
rect 125593 293314 125659 293317
rect 117129 293312 125659 293314
rect -960 293178 480 293268
rect 117129 293256 117134 293312
rect 117190 293256 125598 293312
rect 125654 293256 125659 293312
rect 117129 293254 125659 293256
rect 117129 293251 117195 293254
rect 125593 293251 125659 293254
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 97901 293178 97967 293181
rect 126237 293178 126303 293181
rect 97901 293176 126303 293178
rect 97901 293120 97906 293176
rect 97962 293120 126242 293176
rect 126298 293120 126303 293176
rect 97901 293118 126303 293120
rect 97901 293115 97967 293118
rect 126237 293115 126303 293118
rect 80973 292634 81039 292637
rect 124806 292634 124812 292636
rect 80973 292632 124812 292634
rect 80973 292576 80978 292632
rect 81034 292576 124812 292632
rect 80973 292574 124812 292576
rect 80973 292571 81039 292574
rect 124806 292572 124812 292574
rect 124876 292572 124882 292636
rect 71681 292362 71747 292365
rect 70718 292360 71747 292362
rect 70718 292304 71686 292360
rect 71742 292304 71747 292360
rect 70718 292302 71747 292304
rect 70718 291788 70778 292302
rect 71681 292299 71747 292302
rect 116577 292090 116643 292093
rect 130469 292090 130535 292093
rect 116577 292088 130535 292090
rect 116577 292032 116582 292088
rect 116638 292032 130474 292088
rect 130530 292032 130535 292088
rect 116577 292030 130535 292032
rect 116577 292027 116643 292030
rect 130469 292027 130535 292030
rect 121453 291818 121519 291821
rect 119876 291816 121519 291818
rect 119876 291760 121458 291816
rect 121514 291760 121519 291816
rect 119876 291758 121519 291760
rect 121453 291755 121519 291758
rect 322841 291682 322907 291685
rect 319884 291680 322907 291682
rect 319884 291624 322846 291680
rect 322902 291624 322907 291680
rect 319884 291622 322907 291624
rect 322841 291619 322907 291622
rect 121545 291138 121611 291141
rect 119876 291136 121611 291138
rect 67633 290866 67699 290869
rect 70350 290866 70410 291108
rect 119876 291080 121550 291136
rect 121606 291080 121611 291136
rect 119876 291078 121611 291080
rect 121545 291075 121611 291078
rect 197445 291002 197511 291005
rect 197445 291000 200100 291002
rect 197445 290944 197450 291000
rect 197506 290944 200100 291000
rect 197445 290942 200100 290944
rect 197445 290939 197511 290942
rect 67633 290864 70410 290866
rect 67633 290808 67638 290864
rect 67694 290808 70410 290864
rect 67633 290806 70410 290808
rect 67633 290803 67699 290806
rect 121453 290458 121519 290461
rect 119876 290456 121519 290458
rect 67633 290186 67699 290189
rect 70166 290186 70226 290428
rect 119876 290400 121458 290456
rect 121514 290400 121519 290456
rect 119876 290398 121519 290400
rect 121453 290395 121519 290398
rect 67633 290184 70226 290186
rect 67633 290128 67638 290184
rect 67694 290128 70226 290184
rect 67633 290126 70226 290128
rect 67633 290123 67699 290126
rect 120809 289778 120875 289781
rect 119876 289776 120875 289778
rect 69238 289444 69244 289508
rect 69308 289506 69314 289508
rect 70350 289506 70410 289748
rect 119876 289720 120814 289776
rect 120870 289720 120875 289776
rect 119876 289718 120875 289720
rect 120809 289715 120875 289718
rect 322841 289642 322907 289645
rect 319884 289640 322907 289642
rect 319884 289584 322846 289640
rect 322902 289584 322907 289640
rect 319884 289582 322907 289584
rect 322841 289579 322907 289582
rect 69308 289446 70410 289506
rect 69308 289444 69314 289446
rect 121545 289098 121611 289101
rect 119876 289096 121611 289098
rect 67633 288826 67699 288829
rect 70166 288826 70226 289068
rect 119876 289040 121550 289096
rect 121606 289040 121611 289096
rect 119876 289038 121611 289040
rect 121545 289035 121611 289038
rect 197445 288962 197511 288965
rect 197445 288960 200100 288962
rect 197445 288904 197450 288960
rect 197506 288904 200100 288960
rect 197445 288902 200100 288904
rect 197445 288899 197511 288902
rect 67633 288824 70226 288826
rect 67633 288768 67638 288824
rect 67694 288768 70226 288824
rect 67633 288766 70226 288768
rect 67633 288763 67699 288766
rect 121453 288418 121519 288421
rect 119876 288416 121519 288418
rect 68645 288146 68711 288149
rect 70350 288146 70410 288388
rect 119876 288360 121458 288416
rect 121514 288360 121519 288416
rect 119876 288358 121519 288360
rect 121453 288355 121519 288358
rect 68645 288144 70410 288146
rect 68645 288088 68650 288144
rect 68706 288088 70410 288144
rect 68645 288086 70410 288088
rect 68645 288083 68711 288086
rect 121545 287738 121611 287741
rect 119876 287736 121611 287738
rect 67633 287466 67699 287469
rect 70166 287466 70226 287708
rect 119876 287680 121550 287736
rect 121606 287680 121611 287736
rect 119876 287678 121611 287680
rect 121545 287675 121611 287678
rect 67633 287464 70226 287466
rect 67633 287408 67638 287464
rect 67694 287408 70226 287464
rect 67633 287406 70226 287408
rect 67633 287403 67699 287406
rect 67817 287058 67883 287061
rect 69982 287058 70226 287070
rect 120717 287058 120783 287061
rect 67817 287056 70226 287058
rect 67817 287000 67822 287056
rect 67878 287010 70226 287056
rect 119876 287056 120783 287058
rect 67878 287000 70042 287010
rect 67817 286998 70042 287000
rect 119876 287000 120722 287056
rect 120778 287000 120783 287056
rect 119876 286998 120783 287000
rect 67817 286995 67883 286998
rect 120717 286995 120783 286998
rect 197445 286922 197511 286925
rect 321553 286922 321619 286925
rect 197445 286920 200100 286922
rect 197445 286864 197450 286920
rect 197506 286864 200100 286920
rect 197445 286862 200100 286864
rect 319884 286920 321619 286922
rect 319884 286864 321558 286920
rect 321614 286864 321619 286920
rect 319884 286862 321619 286864
rect 197445 286859 197511 286862
rect 321553 286859 321619 286862
rect 67725 286786 67791 286789
rect 67725 286784 70226 286786
rect 67725 286728 67730 286784
rect 67786 286728 70226 286784
rect 67725 286726 70226 286728
rect 67725 286723 67791 286726
rect 70166 286348 70226 286726
rect 122741 286378 122807 286381
rect 119876 286376 122807 286378
rect 119876 286320 122746 286376
rect 122802 286320 122807 286376
rect 119876 286318 122807 286320
rect 122741 286315 122807 286318
rect 67633 286106 67699 286109
rect 67633 286104 70226 286106
rect 67633 286048 67638 286104
rect 67694 286048 70226 286104
rect 67633 286046 70226 286048
rect 67633 286043 67699 286046
rect 70166 285668 70226 286046
rect 121545 285698 121611 285701
rect 119876 285696 121611 285698
rect 119876 285640 121550 285696
rect 121606 285640 121611 285696
rect 119876 285638 121611 285640
rect 121545 285635 121611 285638
rect 67633 285426 67699 285429
rect 67633 285424 70226 285426
rect 67633 285368 67638 285424
rect 67694 285368 70226 285424
rect 67633 285366 70226 285368
rect 67633 285363 67699 285366
rect 70166 284988 70226 285366
rect 583520 285276 584960 285516
rect 121453 285018 121519 285021
rect 322197 285018 322263 285021
rect 119876 285016 121519 285018
rect 119876 284960 121458 285016
rect 121514 284960 121519 285016
rect 119876 284958 121519 284960
rect 319884 285016 322263 285018
rect 319884 284960 322202 285016
rect 322258 284960 322263 285016
rect 319884 284958 322263 284960
rect 121453 284955 121519 284958
rect 322197 284955 322263 284958
rect 153193 284882 153259 284885
rect 196566 284882 196572 284884
rect 153193 284880 196572 284882
rect 153193 284824 153198 284880
rect 153254 284824 196572 284880
rect 153193 284822 196572 284824
rect 153193 284819 153259 284822
rect 196566 284820 196572 284822
rect 196636 284820 196642 284884
rect 67633 284474 67699 284477
rect 67633 284472 70226 284474
rect 67633 284416 67638 284472
rect 67694 284416 70226 284472
rect 67633 284414 70226 284416
rect 67633 284411 67699 284414
rect 70166 284308 70226 284414
rect 121545 284338 121611 284341
rect 119876 284336 121611 284338
rect 119876 284280 121550 284336
rect 121606 284280 121611 284336
rect 119876 284278 121611 284280
rect 121545 284275 121611 284278
rect 197445 284202 197511 284205
rect 197445 284200 200100 284202
rect 197445 284144 197450 284200
rect 197506 284144 200100 284200
rect 197445 284142 200100 284144
rect 197445 284139 197511 284142
rect 70526 284004 70532 284068
rect 70596 284004 70602 284068
rect 70534 283628 70594 284004
rect 121453 283658 121519 283661
rect 119876 283656 121519 283658
rect 119876 283600 121458 283656
rect 121514 283600 121519 283656
rect 119876 283598 121519 283600
rect 121453 283595 121519 283598
rect 67449 283386 67515 283389
rect 67449 283384 70226 283386
rect 67449 283328 67454 283384
rect 67510 283328 70226 283384
rect 67449 283326 70226 283328
rect 67449 283323 67515 283326
rect 70166 282948 70226 283326
rect 121453 282978 121519 282981
rect 322473 282978 322539 282981
rect 119876 282976 121519 282978
rect 119876 282920 121458 282976
rect 121514 282920 121519 282976
rect 119876 282918 121519 282920
rect 319884 282976 322539 282978
rect 319884 282920 322478 282976
rect 322534 282920 322539 282976
rect 319884 282918 322539 282920
rect 121453 282915 121519 282918
rect 322473 282915 322539 282918
rect 122189 282298 122255 282301
rect 119876 282296 122255 282298
rect 119876 282240 122194 282296
rect 122250 282240 122255 282296
rect 119876 282238 122255 282240
rect 122189 282235 122255 282238
rect 67633 282162 67699 282165
rect 197445 282162 197511 282165
rect 67633 282160 70226 282162
rect 67633 282104 67638 282160
rect 67694 282104 70226 282160
rect 67633 282102 70226 282104
rect 67633 282099 67699 282102
rect 70166 281588 70226 282102
rect 197445 282160 200100 282162
rect 197445 282104 197450 282160
rect 197506 282104 200100 282160
rect 197445 282102 200100 282104
rect 197445 282099 197511 282102
rect 121453 281618 121519 281621
rect 119876 281616 121519 281618
rect 119876 281560 121458 281616
rect 121514 281560 121519 281616
rect 119876 281558 121519 281560
rect 121453 281555 121519 281558
rect 69197 281346 69263 281349
rect 69197 281344 70226 281346
rect 69197 281288 69202 281344
rect 69258 281288 70226 281344
rect 69197 281286 70226 281288
rect 69197 281283 69263 281286
rect 70166 280908 70226 281286
rect 121545 280938 121611 280941
rect 119876 280936 121611 280938
rect 119876 280880 121550 280936
rect 121606 280880 121611 280936
rect 119876 280878 121611 280880
rect 121545 280875 121611 280878
rect 322473 280802 322539 280805
rect 319884 280800 322539 280802
rect 319884 280744 322478 280800
rect 322534 280744 322539 280800
rect 319884 280742 322539 280744
rect 322473 280739 322539 280742
rect 67633 280394 67699 280397
rect 67633 280392 70226 280394
rect 67633 280336 67638 280392
rect 67694 280336 70226 280392
rect 67633 280334 70226 280336
rect 67633 280331 67699 280334
rect 70166 280228 70226 280334
rect 121453 280258 121519 280261
rect 119876 280256 121519 280258
rect -960 279972 480 280212
rect 119876 280200 121458 280256
rect 121514 280200 121519 280256
rect 119876 280198 121519 280200
rect 121453 280195 121519 280198
rect 197445 280258 197511 280261
rect 197445 280256 200100 280258
rect 197445 280200 197450 280256
rect 197506 280200 200100 280256
rect 197445 280198 200100 280200
rect 197445 280195 197511 280198
rect 67725 279850 67791 279853
rect 67725 279848 70226 279850
rect 67725 279792 67730 279848
rect 67786 279792 70226 279848
rect 67725 279790 70226 279792
rect 67725 279787 67791 279790
rect 70166 279548 70226 279790
rect 121545 279578 121611 279581
rect 119876 279576 121611 279578
rect 119876 279520 121550 279576
rect 121606 279520 121611 279576
rect 119876 279518 121611 279520
rect 121545 279515 121611 279518
rect 123334 279380 123340 279444
rect 123404 279442 123410 279444
rect 151813 279442 151879 279445
rect 123404 279440 151879 279442
rect 123404 279384 151818 279440
rect 151874 279384 151879 279440
rect 123404 279382 151879 279384
rect 123404 279380 123410 279382
rect 151813 279379 151879 279382
rect 67633 279306 67699 279309
rect 67633 279304 70226 279306
rect 67633 279248 67638 279304
rect 67694 279248 70226 279304
rect 67633 279246 70226 279248
rect 67633 279243 67699 279246
rect 57789 278900 57855 278901
rect 57789 278896 57836 278900
rect 57900 278898 57906 278900
rect 57789 278840 57794 278896
rect 57789 278836 57836 278840
rect 57900 278838 57946 278898
rect 70166 278868 70226 279246
rect 121453 278898 121519 278901
rect 119876 278896 121519 278898
rect 119876 278840 121458 278896
rect 121514 278840 121519 278896
rect 119876 278838 121519 278840
rect 57900 278836 57906 278838
rect 57789 278835 57855 278836
rect 121453 278835 121519 278838
rect 68829 278626 68895 278629
rect 68829 278624 70226 278626
rect 68829 278568 68834 278624
rect 68890 278568 70226 278624
rect 68829 278566 70226 278568
rect 68829 278563 68895 278566
rect 70166 278188 70226 278566
rect 121545 278218 121611 278221
rect 119876 278216 121611 278218
rect 119876 278160 121550 278216
rect 121606 278160 121611 278216
rect 119876 278158 121611 278160
rect 121545 278155 121611 278158
rect 322197 278082 322263 278085
rect 319884 278080 322263 278082
rect 319884 278024 322202 278080
rect 322258 278024 322263 278080
rect 319884 278022 322263 278024
rect 322197 278019 322263 278022
rect 67633 277674 67699 277677
rect 67633 277672 70226 277674
rect 67633 277616 67638 277672
rect 67694 277616 70226 277672
rect 67633 277614 70226 277616
rect 67633 277611 67699 277614
rect 70166 277508 70226 277614
rect 120809 277538 120875 277541
rect 119876 277536 120875 277538
rect 119876 277480 120814 277536
rect 120870 277480 120875 277536
rect 119876 277478 120875 277480
rect 120809 277475 120875 277478
rect 197445 277538 197511 277541
rect 197445 277536 200100 277538
rect 197445 277480 197450 277536
rect 197506 277480 200100 277536
rect 197445 277478 200100 277480
rect 197445 277475 197511 277478
rect 67817 276994 67883 276997
rect 67817 276992 70226 276994
rect 67817 276936 67822 276992
rect 67878 276936 70226 276992
rect 67817 276934 70226 276936
rect 67817 276931 67883 276934
rect 70166 276828 70226 276934
rect 121453 276858 121519 276861
rect 119876 276856 121519 276858
rect 119876 276800 121458 276856
rect 121514 276800 121519 276856
rect 119876 276798 121519 276800
rect 121453 276795 121519 276798
rect 68737 276586 68803 276589
rect 68737 276584 70226 276586
rect 68737 276528 68742 276584
rect 68798 276528 70226 276584
rect 68737 276526 70226 276528
rect 68737 276523 68803 276526
rect 70166 276148 70226 276526
rect 121453 276178 121519 276181
rect 119876 276176 121519 276178
rect 119876 276120 121458 276176
rect 121514 276120 121519 276176
rect 119876 276118 121519 276120
rect 121453 276115 121519 276118
rect 322841 276042 322907 276045
rect 319884 276040 322907 276042
rect 319884 275984 322846 276040
rect 322902 275984 322907 276040
rect 319884 275982 322907 275984
rect 322841 275979 322907 275982
rect 67633 275906 67699 275909
rect 67633 275904 70226 275906
rect 67633 275848 67638 275904
rect 67694 275848 70226 275904
rect 67633 275846 70226 275848
rect 67633 275843 67699 275846
rect 70166 275468 70226 275846
rect 121545 275498 121611 275501
rect 119876 275496 121611 275498
rect 119876 275440 121550 275496
rect 121606 275440 121611 275496
rect 119876 275438 121611 275440
rect 121545 275435 121611 275438
rect 197353 275362 197419 275365
rect 197353 275360 200100 275362
rect 197353 275304 197358 275360
rect 197414 275304 200100 275360
rect 197353 275302 200100 275304
rect 197353 275299 197419 275302
rect 67633 274954 67699 274957
rect 67633 274952 70226 274954
rect 67633 274896 67638 274952
rect 67694 274896 70226 274952
rect 67633 274894 70226 274896
rect 67633 274891 67699 274894
rect 70166 274788 70226 274894
rect 121453 274818 121519 274821
rect 119876 274816 121519 274818
rect 119876 274760 121458 274816
rect 121514 274760 121519 274816
rect 119876 274758 121519 274760
rect 121453 274755 121519 274758
rect 67725 274546 67791 274549
rect 67725 274544 70226 274546
rect 67725 274488 67730 274544
rect 67786 274488 70226 274544
rect 67725 274486 70226 274488
rect 67725 274483 67791 274486
rect 70166 274108 70226 274486
rect 121545 274138 121611 274141
rect 322381 274138 322447 274141
rect 119876 274136 121611 274138
rect 119876 274080 121550 274136
rect 121606 274080 121611 274136
rect 119876 274078 121611 274080
rect 319884 274136 322447 274138
rect 319884 274080 322386 274136
rect 322442 274080 322447 274136
rect 319884 274078 322447 274080
rect 121545 274075 121611 274078
rect 322381 274075 322447 274078
rect 67633 273594 67699 273597
rect 67633 273592 70226 273594
rect 67633 273536 67638 273592
rect 67694 273536 70226 273592
rect 67633 273534 70226 273536
rect 67633 273531 67699 273534
rect 70166 273428 70226 273534
rect 121453 273458 121519 273461
rect 119876 273456 121519 273458
rect 119876 273400 121458 273456
rect 121514 273400 121519 273456
rect 119876 273398 121519 273400
rect 121453 273395 121519 273398
rect 197353 273322 197419 273325
rect 197353 273320 200100 273322
rect 197353 273264 197358 273320
rect 197414 273264 200100 273320
rect 197353 273262 200100 273264
rect 197353 273259 197419 273262
rect 121453 272778 121519 272781
rect 119876 272776 121519 272778
rect 68737 272234 68803 272237
rect 70166 272234 70226 272748
rect 119876 272720 121458 272776
rect 121514 272720 121519 272776
rect 119876 272718 121519 272720
rect 121453 272715 121519 272718
rect 68737 272232 70226 272234
rect 68737 272176 68742 272232
rect 68798 272176 70226 272232
rect 68737 272174 70226 272176
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 68737 272171 68803 272174
rect 580165 272171 580231 272174
rect 122281 272098 122347 272101
rect 119876 272096 122347 272098
rect 67449 271962 67515 271965
rect 67449 271960 69858 271962
rect 67449 271904 67454 271960
rect 67510 271904 69858 271960
rect 67449 271902 69858 271904
rect 67449 271899 67515 271902
rect 69798 271826 69858 271902
rect 70350 271826 70410 272068
rect 119876 272040 122286 272096
rect 122342 272040 122347 272096
rect 583520 272084 584960 272174
rect 119876 272038 122347 272040
rect 122281 272035 122347 272038
rect 69798 271766 70410 271826
rect 121453 271418 121519 271421
rect 119876 271416 121519 271418
rect 67633 271010 67699 271013
rect 70166 271010 70226 271388
rect 119876 271360 121458 271416
rect 121514 271360 121519 271416
rect 119876 271358 121519 271360
rect 121453 271355 121519 271358
rect 197353 271282 197419 271285
rect 198641 271282 198707 271285
rect 322841 271282 322907 271285
rect 197353 271280 200100 271282
rect 197353 271224 197358 271280
rect 197414 271224 198646 271280
rect 198702 271224 200100 271280
rect 197353 271222 200100 271224
rect 319884 271280 322907 271282
rect 319884 271224 322846 271280
rect 322902 271224 322907 271280
rect 319884 271222 322907 271224
rect 197353 271219 197419 271222
rect 198641 271219 198707 271222
rect 322841 271219 322907 271222
rect 67633 271008 70226 271010
rect 67633 270952 67638 271008
rect 67694 270952 70226 271008
rect 67633 270950 70226 270952
rect 67633 270947 67699 270950
rect 67725 270874 67791 270877
rect 67725 270872 70226 270874
rect 67725 270816 67730 270872
rect 67786 270816 70226 270872
rect 67725 270814 70226 270816
rect 67725 270811 67791 270814
rect 70166 270708 70226 270814
rect 68185 270194 68251 270197
rect 68185 270192 70226 270194
rect 68185 270136 68190 270192
rect 68246 270136 70226 270192
rect 68185 270134 70226 270136
rect 68185 270131 68251 270134
rect 70166 270028 70226 270134
rect 121545 270058 121611 270061
rect 119876 270056 121611 270058
rect 119876 270000 121550 270056
rect 121606 270000 121611 270056
rect 119876 269998 121611 270000
rect 121545 269995 121611 269998
rect 67725 269786 67791 269789
rect 67725 269784 70226 269786
rect 67725 269728 67730 269784
rect 67786 269728 70226 269784
rect 67725 269726 70226 269728
rect 67725 269723 67791 269726
rect 70166 269348 70226 269726
rect 120717 269378 120783 269381
rect 119876 269376 120783 269378
rect 119876 269320 120722 269376
rect 120778 269320 120783 269376
rect 119876 269318 120783 269320
rect 120717 269315 120783 269318
rect 322841 269242 322907 269245
rect 319884 269240 322907 269242
rect 319884 269184 322846 269240
rect 322902 269184 322907 269240
rect 319884 269182 322907 269184
rect 322841 269179 322907 269182
rect 68553 268834 68619 268837
rect 68553 268832 70226 268834
rect 68553 268776 68558 268832
rect 68614 268776 70226 268832
rect 68553 268774 70226 268776
rect 68553 268771 68619 268774
rect 70166 268668 70226 268774
rect 121453 268698 121519 268701
rect 119876 268696 121519 268698
rect 119876 268640 121458 268696
rect 121514 268640 121519 268696
rect 119876 268638 121519 268640
rect 121453 268635 121519 268638
rect 197353 268562 197419 268565
rect 197353 268560 200100 268562
rect 197353 268504 197358 268560
rect 197414 268504 200100 268560
rect 197353 268502 200100 268504
rect 197353 268499 197419 268502
rect 67633 268426 67699 268429
rect 67633 268424 70226 268426
rect 67633 268368 67638 268424
rect 67694 268368 70226 268424
rect 67633 268366 70226 268368
rect 67633 268363 67699 268366
rect 70166 267988 70226 268366
rect 121453 268018 121519 268021
rect 119876 268016 121519 268018
rect 119876 267960 121458 268016
rect 121514 267960 121519 268016
rect 119876 267958 121519 267960
rect 121453 267955 121519 267958
rect 121545 267338 121611 267341
rect 322473 267338 322539 267341
rect 119876 267336 121611 267338
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 67633 267066 67699 267069
rect 70166 267066 70226 267308
rect 119876 267280 121550 267336
rect 121606 267280 121611 267336
rect 119876 267278 121611 267280
rect 319884 267336 322539 267338
rect 319884 267280 322478 267336
rect 322534 267280 322539 267336
rect 319884 267278 322539 267280
rect 121545 267275 121611 267278
rect 322473 267275 322539 267278
rect 67633 267064 70226 267066
rect 67633 267008 67638 267064
rect 67694 267008 70226 267064
rect 67633 267006 70226 267008
rect 67633 267003 67699 267006
rect 67725 266930 67791 266933
rect 67725 266928 70226 266930
rect 67725 266872 67730 266928
rect 67786 266872 70226 266928
rect 67725 266870 70226 266872
rect 67725 266867 67791 266870
rect 70166 266628 70226 266870
rect 121453 266658 121519 266661
rect 119876 266656 121519 266658
rect 119876 266600 121458 266656
rect 121514 266600 121519 266656
rect 119876 266598 121519 266600
rect 121453 266595 121519 266598
rect 197353 266522 197419 266525
rect 197353 266520 200100 266522
rect 197353 266464 197358 266520
rect 197414 266464 200100 266520
rect 197353 266462 200100 266464
rect 197353 266459 197419 266462
rect 121545 265978 121611 265981
rect 119876 265976 121611 265978
rect 67633 265434 67699 265437
rect 70166 265434 70226 265948
rect 119876 265920 121550 265976
rect 121606 265920 121611 265976
rect 119876 265918 121611 265920
rect 121545 265915 121611 265918
rect 67633 265432 70226 265434
rect 67633 265376 67638 265432
rect 67694 265376 70226 265432
rect 67633 265374 70226 265376
rect 67633 265371 67699 265374
rect 121453 265298 121519 265301
rect 119876 265296 121519 265298
rect 67725 265026 67791 265029
rect 70350 265026 70410 265268
rect 119876 265240 121458 265296
rect 121514 265240 121519 265296
rect 119876 265238 121519 265240
rect 121453 265235 121519 265238
rect 322473 265162 322539 265165
rect 319884 265160 322539 265162
rect 319884 265104 322478 265160
rect 322534 265104 322539 265160
rect 319884 265102 322539 265104
rect 322473 265099 322539 265102
rect 67725 265024 70410 265026
rect 67725 264968 67730 265024
rect 67786 264968 70410 265024
rect 67725 264966 70410 264968
rect 67725 264963 67791 264966
rect 67725 264210 67791 264213
rect 70166 264210 70226 264588
rect 67725 264208 70226 264210
rect 67725 264152 67730 264208
rect 67786 264152 70226 264208
rect 67725 264150 70226 264152
rect 67725 264147 67791 264150
rect 119846 264074 119906 264588
rect 197353 264482 197419 264485
rect 197353 264480 200100 264482
rect 197353 264424 197358 264480
rect 197414 264424 200100 264480
rect 197353 264422 200100 264424
rect 197353 264419 197419 264422
rect 125726 264074 125732 264076
rect 119846 264014 125732 264074
rect 125726 264012 125732 264014
rect 125796 264012 125802 264076
rect 121545 263938 121611 263941
rect 119876 263936 121611 263938
rect 67633 263666 67699 263669
rect 70350 263666 70410 263908
rect 119876 263880 121550 263936
rect 121606 263880 121611 263936
rect 119876 263878 121611 263880
rect 121545 263875 121611 263878
rect 67633 263664 70410 263666
rect 67633 263608 67638 263664
rect 67694 263608 70410 263664
rect 67633 263606 70410 263608
rect 67633 263603 67699 263606
rect 67633 263530 67699 263533
rect 67633 263528 70226 263530
rect 67633 263472 67638 263528
rect 67694 263472 70226 263528
rect 67633 263470 70226 263472
rect 67633 263467 67699 263470
rect 70166 263228 70226 263470
rect 121453 263258 121519 263261
rect 119876 263256 121519 263258
rect 119876 263200 121458 263256
rect 121514 263200 121519 263256
rect 119876 263198 121519 263200
rect 121453 263195 121519 263198
rect 121453 262578 121519 262581
rect 119876 262576 121519 262578
rect 67633 262306 67699 262309
rect 70166 262306 70226 262548
rect 119876 262520 121458 262576
rect 121514 262520 121519 262576
rect 119876 262518 121519 262520
rect 121453 262515 121519 262518
rect 322473 262442 322539 262445
rect 319884 262440 322539 262442
rect 319884 262384 322478 262440
rect 322534 262384 322539 262440
rect 319884 262382 322539 262384
rect 322473 262379 322539 262382
rect 67633 262304 70226 262306
rect 67633 262248 67638 262304
rect 67694 262248 70226 262304
rect 67633 262246 70226 262248
rect 67633 262243 67699 262246
rect 67725 262170 67791 262173
rect 67725 262168 70226 262170
rect 67725 262112 67730 262168
rect 67786 262112 70226 262168
rect 67725 262110 70226 262112
rect 67725 262107 67791 262110
rect 70166 261868 70226 262110
rect 121453 261898 121519 261901
rect 119876 261896 121519 261898
rect 119876 261840 121458 261896
rect 121514 261840 121519 261896
rect 119876 261838 121519 261840
rect 121453 261835 121519 261838
rect 197353 261762 197419 261765
rect 197353 261760 200100 261762
rect 197353 261704 197358 261760
rect 197414 261704 200100 261760
rect 197353 261702 200100 261704
rect 197353 261699 197419 261702
rect 67357 261626 67423 261629
rect 67357 261624 70226 261626
rect 67357 261568 67362 261624
rect 67418 261568 70226 261624
rect 67357 261566 70226 261568
rect 67357 261563 67423 261566
rect 70166 261188 70226 261566
rect 121545 261218 121611 261221
rect 119876 261216 121611 261218
rect 119876 261160 121550 261216
rect 121606 261160 121611 261216
rect 119876 261158 121611 261160
rect 121545 261155 121611 261158
rect 67633 260810 67699 260813
rect 67633 260808 70226 260810
rect 67633 260752 67638 260808
rect 67694 260752 70226 260808
rect 67633 260750 70226 260752
rect 67633 260747 67699 260750
rect 70166 260508 70226 260750
rect 121453 260538 121519 260541
rect 119876 260536 121519 260538
rect 119876 260480 121458 260536
rect 121514 260480 121519 260536
rect 119876 260478 121519 260480
rect 121453 260475 121519 260478
rect 322565 260402 322631 260405
rect 319884 260400 322631 260402
rect 319884 260344 322570 260400
rect 322626 260344 322631 260400
rect 319884 260342 322631 260344
rect 322565 260339 322631 260342
rect 69105 260266 69171 260269
rect 69105 260264 70226 260266
rect 69105 260208 69110 260264
rect 69166 260208 70226 260264
rect 69105 260206 70226 260208
rect 69105 260203 69171 260206
rect 70166 259828 70226 260206
rect 121453 259858 121519 259861
rect 119876 259856 121519 259858
rect 119876 259800 121458 259856
rect 121514 259800 121519 259856
rect 119876 259798 121519 259800
rect 121453 259795 121519 259798
rect 197353 259722 197419 259725
rect 197353 259720 200100 259722
rect 197353 259664 197358 259720
rect 197414 259664 200100 259720
rect 197353 259662 200100 259664
rect 197353 259659 197419 259662
rect 121637 259178 121703 259181
rect 119876 259176 121703 259178
rect 67725 258634 67791 258637
rect 70166 258634 70226 259148
rect 119876 259120 121642 259176
rect 121698 259120 121703 259176
rect 119876 259118 121703 259120
rect 121637 259115 121703 259118
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect 67725 258632 70226 258634
rect 67725 258576 67730 258632
rect 67786 258576 70226 258632
rect 67725 258574 70226 258576
rect 67725 258571 67791 258574
rect 121545 258498 121611 258501
rect 119876 258496 121611 258498
rect 70166 258092 70226 258468
rect 119876 258440 121550 258496
rect 121606 258440 121611 258496
rect 119876 258438 121611 258440
rect 121545 258435 121611 258438
rect 324262 258362 324268 258364
rect 319884 258302 324268 258362
rect 324262 258300 324268 258302
rect 324332 258362 324338 258364
rect 324405 258362 324471 258365
rect 324332 258360 324471 258362
rect 324332 258304 324410 258360
rect 324466 258304 324471 258360
rect 324332 258302 324471 258304
rect 324332 258300 324338 258302
rect 324405 258299 324471 258302
rect 70158 258028 70164 258092
rect 70228 258028 70234 258092
rect 67633 257954 67699 257957
rect 67633 257952 70226 257954
rect 67633 257896 67638 257952
rect 67694 257896 70226 257952
rect 67633 257894 70226 257896
rect 67633 257891 67699 257894
rect 70166 257788 70226 257894
rect 121545 257818 121611 257821
rect 119876 257816 121611 257818
rect 119876 257760 121550 257816
rect 121606 257760 121611 257816
rect 119876 257758 121611 257760
rect 121545 257755 121611 257758
rect 197353 257682 197419 257685
rect 197353 257680 200100 257682
rect 197353 257624 197358 257680
rect 197414 257624 200100 257680
rect 197353 257622 200100 257624
rect 197353 257619 197419 257622
rect 121453 257138 121519 257141
rect 119876 257136 121519 257138
rect 68001 256866 68067 256869
rect 70166 256866 70226 257108
rect 119876 257080 121458 257136
rect 121514 257080 121519 257136
rect 119876 257078 121519 257080
rect 121453 257075 121519 257078
rect 68001 256864 70226 256866
rect 68001 256808 68006 256864
rect 68062 256808 70226 256864
rect 68001 256806 70226 256808
rect 68001 256803 68067 256806
rect 121453 256458 121519 256461
rect 119876 256456 121519 256458
rect 69197 255914 69263 255917
rect 70166 255914 70226 256428
rect 119876 256400 121458 256456
rect 121514 256400 121519 256456
rect 119876 256398 121519 256400
rect 121453 256395 121519 256398
rect 69197 255912 70226 255914
rect 69197 255856 69202 255912
rect 69258 255856 70226 255912
rect 69197 255854 70226 255856
rect 69197 255851 69263 255854
rect 121545 255778 121611 255781
rect 119876 255776 121611 255778
rect 67633 255370 67699 255373
rect 70166 255370 70226 255748
rect 119876 255720 121550 255776
rect 121606 255720 121611 255776
rect 119876 255718 121611 255720
rect 121545 255715 121611 255718
rect 197353 255642 197419 255645
rect 321645 255642 321711 255645
rect 197353 255640 200100 255642
rect 197353 255584 197358 255640
rect 197414 255584 200100 255640
rect 197353 255582 200100 255584
rect 319884 255640 321711 255642
rect 319884 255584 321650 255640
rect 321706 255584 321711 255640
rect 319884 255582 321711 255584
rect 197353 255579 197419 255582
rect 321645 255579 321711 255582
rect 67633 255368 70226 255370
rect 67633 255312 67638 255368
rect 67694 255312 70226 255368
rect 67633 255310 70226 255312
rect 67633 255307 67699 255310
rect 67725 255234 67791 255237
rect 67725 255232 70226 255234
rect 67725 255176 67730 255232
rect 67786 255176 70226 255232
rect 67725 255174 70226 255176
rect 67725 255171 67791 255174
rect 70166 255068 70226 255174
rect 121453 255098 121519 255101
rect 119876 255096 121519 255098
rect 119876 255040 121458 255096
rect 121514 255040 121519 255096
rect 119876 255038 121519 255040
rect 121453 255035 121519 255038
rect 67633 254826 67699 254829
rect 67633 254824 70226 254826
rect 67633 254768 67638 254824
rect 67694 254768 70226 254824
rect 67633 254766 70226 254768
rect 67633 254763 67699 254766
rect 70166 254388 70226 254766
rect 122097 254418 122163 254421
rect 119876 254416 122163 254418
rect 119876 254360 122102 254416
rect 122158 254360 122163 254416
rect 119876 254358 122163 254360
rect 122097 254355 122163 254358
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 67633 253874 67699 253877
rect 67633 253872 70226 253874
rect 67633 253816 67638 253872
rect 67694 253816 70226 253872
rect 67633 253814 70226 253816
rect 67633 253811 67699 253814
rect 70166 253708 70226 253814
rect 121453 253738 121519 253741
rect 119876 253736 121519 253738
rect 119876 253680 121458 253736
rect 121514 253680 121519 253736
rect 119876 253678 121519 253680
rect 121453 253675 121519 253678
rect 120574 253132 120580 253196
rect 120644 253194 120650 253196
rect 143717 253194 143783 253197
rect 120644 253192 143783 253194
rect 120644 253136 143722 253192
rect 143778 253136 143783 253192
rect 120644 253134 143783 253136
rect 120644 253132 120650 253134
rect 143717 253131 143783 253134
rect 121545 253058 121611 253061
rect 319302 253060 319362 253572
rect 119876 253056 121611 253058
rect 61694 252724 61700 252788
rect 61764 252786 61770 252788
rect 70166 252786 70226 253028
rect 119876 253000 121550 253056
rect 121606 253000 121611 253056
rect 119876 252998 121611 253000
rect 121545 252995 121611 252998
rect 319294 252996 319300 253060
rect 319364 252996 319370 253060
rect 197353 252922 197419 252925
rect 197353 252920 200100 252922
rect 197353 252864 197358 252920
rect 197414 252864 200100 252920
rect 197353 252862 200100 252864
rect 197353 252859 197419 252862
rect 61764 252726 70226 252786
rect 61764 252724 61770 252726
rect 121453 252378 121519 252381
rect 119876 252376 121519 252378
rect 67633 251834 67699 251837
rect 70166 251834 70226 252348
rect 119876 252320 121458 252376
rect 121514 252320 121519 252376
rect 119876 252318 121519 252320
rect 121453 252315 121519 252318
rect 67633 251832 70226 251834
rect 67633 251776 67638 251832
rect 67694 251776 70226 251832
rect 67633 251774 70226 251776
rect 67633 251771 67699 251774
rect 121453 251698 121519 251701
rect 119876 251696 121519 251698
rect 68553 251426 68619 251429
rect 70350 251426 70410 251668
rect 119876 251640 121458 251696
rect 121514 251640 121519 251696
rect 119876 251638 121519 251640
rect 121453 251635 121519 251638
rect 322473 251562 322539 251565
rect 319884 251560 322539 251562
rect 319884 251504 322478 251560
rect 322534 251504 322539 251560
rect 319884 251502 322539 251504
rect 322473 251499 322539 251502
rect 68553 251424 70410 251426
rect 68553 251368 68558 251424
rect 68614 251368 70410 251424
rect 68553 251366 70410 251368
rect 68553 251363 68619 251366
rect 67725 251154 67791 251157
rect 67725 251152 70226 251154
rect 67725 251096 67730 251152
rect 67786 251096 70226 251152
rect 67725 251094 70226 251096
rect 67725 251091 67791 251094
rect 70166 250988 70226 251094
rect 120165 251018 120231 251021
rect 120625 251018 120691 251021
rect 119876 251016 120691 251018
rect 119876 250960 120170 251016
rect 120226 250960 120630 251016
rect 120686 250960 120691 251016
rect 119876 250958 120691 250960
rect 120165 250955 120231 250958
rect 120625 250955 120691 250958
rect 195830 250820 195836 250884
rect 195900 250882 195906 250884
rect 195900 250822 200100 250882
rect 195900 250820 195906 250822
rect 166441 250474 166507 250477
rect 195830 250474 195836 250476
rect 166441 250472 195836 250474
rect 166441 250416 166446 250472
rect 166502 250416 195836 250472
rect 166441 250414 195836 250416
rect 166441 250411 166507 250414
rect 195830 250412 195836 250414
rect 195900 250412 195906 250476
rect 121453 250338 121519 250341
rect 119876 250336 121519 250338
rect 68461 249930 68527 249933
rect 70166 249930 70226 250308
rect 119876 250280 121458 250336
rect 121514 250280 121519 250336
rect 119876 250278 121519 250280
rect 121453 250275 121519 250278
rect 68461 249928 70226 249930
rect 68461 249872 68466 249928
rect 68522 249872 70226 249928
rect 68461 249870 70226 249872
rect 68461 249867 68527 249870
rect 120073 249658 120139 249661
rect 119876 249656 120139 249658
rect 67633 249114 67699 249117
rect 70166 249114 70226 249628
rect 119876 249600 120078 249656
rect 120134 249600 120139 249656
rect 119876 249598 120139 249600
rect 120073 249595 120139 249598
rect 67633 249112 70226 249114
rect 67633 249056 67638 249112
rect 67694 249056 70226 249112
rect 67633 249054 70226 249056
rect 67633 249051 67699 249054
rect 121545 248978 121611 248981
rect 119876 248976 121611 248978
rect 67357 248706 67423 248709
rect 70166 248706 70226 248948
rect 119876 248920 121550 248976
rect 121606 248920 121611 248976
rect 119876 248918 121611 248920
rect 121545 248915 121611 248918
rect 197353 248842 197419 248845
rect 320265 248842 320331 248845
rect 197353 248840 200100 248842
rect 197353 248784 197358 248840
rect 197414 248784 200100 248840
rect 197353 248782 200100 248784
rect 319884 248840 320331 248842
rect 319884 248784 320270 248840
rect 320326 248784 320331 248840
rect 319884 248782 320331 248784
rect 197353 248779 197419 248782
rect 320265 248779 320331 248782
rect 67357 248704 70226 248706
rect 67357 248648 67362 248704
rect 67418 248648 70226 248704
rect 67357 248646 70226 248648
rect 67357 248643 67423 248646
rect 121453 248298 121519 248301
rect 119876 248296 121519 248298
rect 67725 247754 67791 247757
rect 70166 247754 70226 248268
rect 119876 248240 121458 248296
rect 121514 248240 121519 248296
rect 119876 248238 121519 248240
rect 121453 248235 121519 248238
rect 67725 247752 70226 247754
rect 67725 247696 67730 247752
rect 67786 247696 70226 247752
rect 67725 247694 70226 247696
rect 67725 247691 67791 247694
rect 121545 247618 121611 247621
rect 119876 247616 121611 247618
rect 67633 247210 67699 247213
rect 70166 247210 70226 247588
rect 119876 247560 121550 247616
rect 121606 247560 121611 247616
rect 119876 247558 121611 247560
rect 121545 247555 121611 247558
rect 67633 247208 70226 247210
rect 67633 247152 67638 247208
rect 67694 247152 70226 247208
rect 67633 247150 70226 247152
rect 67633 247147 67699 247150
rect 121545 246938 121611 246941
rect 119876 246936 121611 246938
rect 67725 246394 67791 246397
rect 70166 246394 70226 246908
rect 119876 246880 121550 246936
rect 121606 246880 121611 246936
rect 119876 246878 121611 246880
rect 121545 246875 121611 246878
rect 320357 246802 320423 246805
rect 319884 246800 320423 246802
rect 319884 246744 320362 246800
rect 320418 246744 320423 246800
rect 319884 246742 320423 246744
rect 320357 246739 320423 246742
rect 67725 246392 70226 246394
rect 67725 246336 67730 246392
rect 67786 246336 70226 246392
rect 67725 246334 70226 246336
rect 67725 246331 67791 246334
rect 121453 246258 121519 246261
rect 119876 246256 121519 246258
rect 67633 245850 67699 245853
rect 70166 245850 70226 246228
rect 119876 246200 121458 246256
rect 121514 246200 121519 246256
rect 119876 246198 121519 246200
rect 121453 246195 121519 246198
rect 197353 246258 197419 246261
rect 197353 246256 200100 246258
rect 197353 246200 197358 246256
rect 197414 246200 200100 246256
rect 197353 246198 200100 246200
rect 197353 246195 197419 246198
rect 67633 245848 70226 245850
rect 67633 245792 67638 245848
rect 67694 245792 70226 245848
rect 67633 245790 70226 245792
rect 67633 245787 67699 245790
rect 121453 245578 121519 245581
rect 119876 245576 121519 245578
rect 67633 245306 67699 245309
rect 70350 245306 70410 245548
rect 119876 245520 121458 245576
rect 121514 245520 121519 245576
rect 119876 245518 121519 245520
rect 121453 245515 121519 245518
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 67633 245304 70410 245306
rect 67633 245248 67638 245304
rect 67694 245248 70410 245304
rect 67633 245246 70410 245248
rect 67633 245243 67699 245246
rect 121545 244898 121611 244901
rect 119876 244896 121611 244898
rect 69105 244354 69171 244357
rect 70166 244354 70226 244868
rect 119876 244840 121550 244896
rect 121606 244840 121611 244896
rect 119876 244838 121611 244840
rect 121545 244835 121611 244838
rect 322841 244762 322907 244765
rect 319884 244760 322907 244762
rect 319884 244704 322846 244760
rect 322902 244704 322907 244760
rect 319884 244702 322907 244704
rect 322841 244699 322907 244702
rect 69105 244352 70226 244354
rect 69105 244296 69110 244352
rect 69166 244296 70226 244352
rect 69105 244294 70226 244296
rect 69105 244291 69171 244294
rect 121453 244218 121519 244221
rect 119876 244216 121519 244218
rect 67633 243810 67699 243813
rect 70350 243810 70410 244188
rect 119876 244160 121458 244216
rect 121514 244160 121519 244216
rect 119876 244158 121519 244160
rect 121453 244155 121519 244158
rect 197118 244020 197124 244084
rect 197188 244082 197194 244084
rect 197188 244022 200100 244082
rect 197188 244020 197194 244022
rect 67633 243808 70410 243810
rect 67633 243752 67638 243808
rect 67694 243752 70410 243808
rect 67633 243750 70410 243752
rect 67633 243747 67699 243750
rect 67725 243674 67791 243677
rect 67725 243672 70226 243674
rect 67725 243616 67730 243672
rect 67786 243616 70226 243672
rect 67725 243614 70226 243616
rect 67725 243611 67791 243614
rect 70166 243508 70226 243614
rect 123334 243538 123340 243540
rect 119876 243478 123340 243538
rect 123334 243476 123340 243478
rect 123404 243476 123410 243540
rect 121453 242858 121519 242861
rect 119876 242856 121519 242858
rect 70534 242452 70594 242828
rect 119876 242800 121458 242856
rect 121514 242800 121519 242856
rect 119876 242798 121519 242800
rect 121453 242795 121519 242798
rect 319345 242586 319411 242589
rect 319854 242586 319914 242692
rect 321737 242586 321803 242589
rect 319345 242584 321803 242586
rect 319345 242528 319350 242584
rect 319406 242528 321742 242584
rect 321798 242528 321803 242584
rect 319345 242526 321803 242528
rect 319345 242523 319411 242526
rect 321737 242523 321803 242526
rect 70526 242388 70532 242452
rect 70596 242388 70602 242452
rect 121545 242178 121611 242181
rect 119876 242176 121611 242178
rect 69841 241634 69907 241637
rect 70166 241634 70226 242148
rect 119876 242120 121550 242176
rect 121606 242120 121611 242176
rect 119876 242118 121611 242120
rect 121545 242115 121611 242118
rect 133781 242178 133847 242181
rect 196014 242178 196020 242180
rect 133781 242176 196020 242178
rect 133781 242120 133786 242176
rect 133842 242120 196020 242176
rect 133781 242118 196020 242120
rect 133781 242115 133847 242118
rect 196014 242116 196020 242118
rect 196084 242116 196090 242180
rect 198457 242178 198523 242181
rect 198457 242176 200100 242178
rect 198457 242120 198462 242176
rect 198518 242120 200100 242176
rect 198457 242118 200100 242120
rect 198457 242115 198523 242118
rect 69841 241632 70226 241634
rect 69841 241576 69846 241632
rect 69902 241576 70226 241632
rect 69841 241574 70226 241576
rect 69841 241571 69907 241574
rect 120574 241498 120580 241500
rect 119876 241468 120580 241498
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 68645 240954 68711 240957
rect 70166 240954 70226 241468
rect 119846 241438 120580 241468
rect 119846 241226 119906 241438
rect 120574 241436 120580 241438
rect 120644 241436 120650 241500
rect 120022 241226 120028 241228
rect 119846 241166 120028 241226
rect 120022 241164 120028 241166
rect 120092 241164 120098 241228
rect 68645 240952 70226 240954
rect 68645 240896 68650 240952
rect 68706 240896 70226 240952
rect 68645 240894 70226 240896
rect 68645 240891 68711 240894
rect 121453 240818 121519 240821
rect 119876 240816 121519 240818
rect 70534 240276 70594 240788
rect 119876 240760 121458 240816
rect 121514 240760 121519 240816
rect 119876 240758 121519 240760
rect 121453 240755 121519 240758
rect 147213 240818 147279 240821
rect 200614 240818 200620 240820
rect 147213 240816 200620 240818
rect 147213 240760 147218 240816
rect 147274 240760 200620 240816
rect 147213 240758 200620 240760
rect 147213 240755 147279 240758
rect 200614 240756 200620 240758
rect 200684 240756 200690 240820
rect 70526 240212 70532 240276
rect 70596 240212 70602 240276
rect 121453 240138 121519 240141
rect 119876 240136 121519 240138
rect 119876 240080 121458 240136
rect 121514 240080 121519 240136
rect 119876 240078 121519 240080
rect 121453 240075 121519 240078
rect 329833 240138 329899 240141
rect 330334 240138 330340 240140
rect 329833 240136 330340 240138
rect 329833 240080 329838 240136
rect 329894 240080 330340 240136
rect 329833 240078 330340 240080
rect 329833 240075 329899 240078
rect 330334 240076 330340 240078
rect 330404 240076 330410 240140
rect 321737 240002 321803 240005
rect 319884 240000 321803 240002
rect 319884 239944 321742 240000
rect 321798 239944 321803 240000
rect 319884 239942 321803 239944
rect 321737 239939 321803 239942
rect 327073 240002 327139 240005
rect 327206 240002 327212 240004
rect 327073 240000 327212 240002
rect 327073 239944 327078 240000
rect 327134 239944 327212 240000
rect 327073 239942 327212 239944
rect 327073 239939 327139 239942
rect 327206 239940 327212 239942
rect 327276 239940 327282 240004
rect 152549 239866 152615 239869
rect 201401 239866 201467 239869
rect 152549 239864 201467 239866
rect 152549 239808 152554 239864
rect 152610 239808 201406 239864
rect 201462 239808 201467 239864
rect 152549 239806 201467 239808
rect 152549 239803 152615 239806
rect 201401 239803 201467 239806
rect 197169 239458 197235 239461
rect 204897 239458 204963 239461
rect 197169 239456 204963 239458
rect 197169 239400 197174 239456
rect 197230 239400 204902 239456
rect 204958 239400 204963 239456
rect 197169 239398 204963 239400
rect 197169 239395 197235 239398
rect 204897 239395 204963 239398
rect 196014 238716 196020 238780
rect 196084 238778 196090 238780
rect 252829 238778 252895 238781
rect 196084 238776 252895 238778
rect 196084 238720 252834 238776
rect 252890 238720 252895 238776
rect 196084 238718 252895 238720
rect 196084 238716 196090 238718
rect 252829 238715 252895 238718
rect 71078 238580 71084 238644
rect 71148 238642 71154 238644
rect 140865 238642 140931 238645
rect 71148 238640 140931 238642
rect 71148 238584 140870 238640
rect 140926 238584 140931 238640
rect 71148 238582 140931 238584
rect 71148 238580 71154 238582
rect 140865 238579 140931 238582
rect 144913 238642 144979 238645
rect 305637 238642 305703 238645
rect 144913 238640 305703 238642
rect 144913 238584 144918 238640
rect 144974 238584 305642 238640
rect 305698 238584 305703 238640
rect 144913 238582 305703 238584
rect 144913 238579 144979 238582
rect 305637 238579 305703 238582
rect 184381 238506 184447 238509
rect 244457 238506 244523 238509
rect 184381 238504 244523 238506
rect 184381 238448 184386 238504
rect 184442 238448 244462 238504
rect 244518 238448 244523 238504
rect 184381 238446 244523 238448
rect 184381 238443 184447 238446
rect 244457 238443 244523 238446
rect 188470 237900 188476 237964
rect 188540 237962 188546 237964
rect 207657 237962 207723 237965
rect 188540 237960 207723 237962
rect 188540 237904 207662 237960
rect 207718 237904 207723 237960
rect 188540 237902 207723 237904
rect 188540 237900 188546 237902
rect 207657 237899 207723 237902
rect 140865 237418 140931 237421
rect 141509 237418 141575 237421
rect 140865 237416 141575 237418
rect 140865 237360 140870 237416
rect 140926 237360 141514 237416
rect 141570 237360 141575 237416
rect 140865 237358 141575 237360
rect 140865 237355 140931 237358
rect 141509 237355 141575 237358
rect 63217 237282 63283 237285
rect 323669 237282 323735 237285
rect 63217 237280 323735 237282
rect 63217 237224 63222 237280
rect 63278 237224 323674 237280
rect 323730 237224 323735 237280
rect 63217 237222 323735 237224
rect 63217 237219 63283 237222
rect 323669 237219 323735 237222
rect 86125 237146 86191 237149
rect 325049 237146 325115 237149
rect 86125 237144 325115 237146
rect 86125 237088 86130 237144
rect 86186 237088 325054 237144
rect 325110 237088 325115 237144
rect 86125 237086 325115 237088
rect 86125 237083 86191 237086
rect 325049 237083 325115 237086
rect 68737 236602 68803 236605
rect 255262 236602 255268 236604
rect 68737 236600 255268 236602
rect 68737 236544 68742 236600
rect 68798 236544 255268 236600
rect 68737 236542 255268 236544
rect 68737 236539 68803 236542
rect 255262 236540 255268 236542
rect 255332 236540 255338 236604
rect 160686 235860 160692 235924
rect 160756 235922 160762 235924
rect 227069 235922 227135 235925
rect 160756 235920 227135 235922
rect 160756 235864 227074 235920
rect 227130 235864 227135 235920
rect 160756 235862 227135 235864
rect 160756 235860 160762 235862
rect 227069 235859 227135 235862
rect 56225 235242 56291 235245
rect 211613 235242 211679 235245
rect 56225 235240 211679 235242
rect 56225 235184 56230 235240
rect 56286 235184 211618 235240
rect 211674 235184 211679 235240
rect 56225 235182 211679 235184
rect 56225 235179 56291 235182
rect 211613 235179 211679 235182
rect 57830 234500 57836 234564
rect 57900 234562 57906 234564
rect 293217 234562 293283 234565
rect 57900 234560 293283 234562
rect 57900 234504 293222 234560
rect 293278 234504 293283 234560
rect 57900 234502 293283 234504
rect 57900 234500 57906 234502
rect 293217 234499 293283 234502
rect 75821 234426 75887 234429
rect 133822 234426 133828 234428
rect 75821 234424 133828 234426
rect 75821 234368 75826 234424
rect 75882 234368 133828 234424
rect 75821 234366 133828 234368
rect 75821 234363 75887 234366
rect 133822 234364 133828 234366
rect 133892 234364 133898 234428
rect 163589 234426 163655 234429
rect 333973 234426 334039 234429
rect 163589 234424 334039 234426
rect 163589 234368 163594 234424
rect 163650 234368 333978 234424
rect 334034 234368 334039 234424
rect 163589 234366 334039 234368
rect 163589 234363 163655 234366
rect 333973 234363 334039 234366
rect 200614 234228 200620 234292
rect 200684 234290 200690 234292
rect 327257 234290 327323 234293
rect 327441 234290 327507 234293
rect 200684 234288 327507 234290
rect 200684 234232 327262 234288
rect 327318 234232 327446 234288
rect 327502 234232 327507 234288
rect 200684 234230 327507 234232
rect 200684 234228 200690 234230
rect 327257 234227 327323 234230
rect 327441 234227 327507 234230
rect 71773 233202 71839 233205
rect 289445 233202 289511 233205
rect 71773 233200 289511 233202
rect 71773 233144 71778 233200
rect 71834 233144 289450 233200
rect 289506 233144 289511 233200
rect 71773 233142 289511 233144
rect 71773 233139 71839 233142
rect 289445 233139 289511 233142
rect 176193 233066 176259 233069
rect 265617 233066 265683 233069
rect 176193 233064 265683 233066
rect 176193 233008 176198 233064
rect 176254 233008 265622 233064
rect 265678 233008 265683 233064
rect 176193 233006 265683 233008
rect 176193 233003 176259 233006
rect 265617 233003 265683 233006
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect 91737 231842 91803 231845
rect 299197 231842 299263 231845
rect 91737 231840 299263 231842
rect 91737 231784 91742 231840
rect 91798 231784 299202 231840
rect 299258 231784 299263 231840
rect 91737 231782 299263 231784
rect 91737 231779 91803 231782
rect 299197 231779 299263 231782
rect 162301 231706 162367 231709
rect 318742 231706 318748 231708
rect 162301 231704 318748 231706
rect 162301 231648 162306 231704
rect 162362 231648 318748 231704
rect 162301 231646 318748 231648
rect 162301 231643 162367 231646
rect 318742 231644 318748 231646
rect 318812 231644 318818 231708
rect 166349 230482 166415 230485
rect 324262 230482 324268 230484
rect 166349 230480 324268 230482
rect 166349 230424 166354 230480
rect 166410 230424 324268 230480
rect 166349 230422 324268 230424
rect 166349 230419 166415 230422
rect 324262 230420 324268 230422
rect 324332 230420 324338 230484
rect 70894 228924 70900 228988
rect 70964 228986 70970 228988
rect 198590 228986 198596 228988
rect 70964 228926 198596 228986
rect 70964 228924 70970 228926
rect 198590 228924 198596 228926
rect 198660 228924 198666 228988
rect 198590 228244 198596 228308
rect 198660 228306 198666 228308
rect 251909 228306 251975 228309
rect 198660 228304 251975 228306
rect 198660 228248 251914 228304
rect 251970 228248 251975 228304
rect 198660 228246 251975 228248
rect 198660 228244 198666 228246
rect 251909 228243 251975 228246
rect -960 227884 480 228124
rect 180006 227020 180012 227084
rect 180076 227082 180082 227084
rect 215937 227082 216003 227085
rect 180076 227080 216003 227082
rect 180076 227024 215942 227080
rect 215998 227024 216003 227080
rect 180076 227022 216003 227024
rect 180076 227020 180082 227022
rect 215937 227019 216003 227022
rect 68829 226946 68895 226949
rect 252502 226946 252508 226948
rect 68829 226944 252508 226946
rect 68829 226888 68834 226944
rect 68890 226888 252508 226944
rect 68829 226886 252508 226888
rect 68829 226883 68895 226886
rect 252502 226884 252508 226886
rect 252572 226884 252578 226948
rect 152641 226266 152707 226269
rect 331213 226266 331279 226269
rect 152641 226264 331279 226266
rect 152641 226208 152646 226264
rect 152702 226208 331218 226264
rect 331274 226208 331279 226264
rect 152641 226206 331279 226208
rect 152641 226203 152707 226206
rect 331213 226203 331279 226206
rect 66069 225586 66135 225589
rect 252001 225586 252067 225589
rect 66069 225584 252067 225586
rect 66069 225528 66074 225584
rect 66130 225528 252006 225584
rect 252062 225528 252067 225584
rect 66069 225526 252067 225528
rect 66069 225523 66135 225526
rect 252001 225523 252067 225526
rect 1301 224226 1367 224229
rect 120022 224226 120028 224228
rect 1301 224224 120028 224226
rect 1301 224168 1306 224224
rect 1362 224168 120028 224224
rect 1301 224166 120028 224168
rect 1301 224163 1367 224166
rect 120022 224164 120028 224166
rect 120092 224164 120098 224228
rect 169017 222866 169083 222869
rect 271086 222866 271092 222868
rect 169017 222864 271092 222866
rect 169017 222808 169022 222864
rect 169078 222808 271092 222864
rect 169017 222806 271092 222808
rect 169017 222803 169083 222806
rect 271086 222804 271092 222806
rect 271156 222804 271162 222868
rect 173157 221506 173223 221509
rect 362953 221506 363019 221509
rect 173157 221504 363019 221506
rect 173157 221448 173162 221504
rect 173218 221448 362958 221504
rect 363014 221448 363019 221504
rect 173157 221446 363019 221448
rect 173157 221443 173223 221446
rect 362953 221443 363019 221446
rect 579797 219058 579863 219061
rect 583520 219058 584960 219148
rect 579797 219056 584960 219058
rect 579797 219000 579802 219056
rect 579858 219000 584960 219056
rect 579797 218998 584960 219000
rect 579797 218995 579863 218998
rect 583520 218908 584960 218998
rect 195830 218588 195836 218652
rect 195900 218650 195906 218652
rect 517605 218650 517671 218653
rect 195900 218648 517671 218650
rect 195900 218592 517610 218648
rect 517666 218592 517671 218648
rect 195900 218590 517671 218592
rect 195900 218588 195906 218590
rect 517605 218587 517671 218590
rect 130469 215930 130535 215933
rect 335854 215930 335860 215932
rect 130469 215928 335860 215930
rect 130469 215872 130474 215928
rect 130530 215872 335860 215928
rect 130469 215870 335860 215872
rect 130469 215867 130535 215870
rect 335854 215868 335860 215870
rect 335924 215868 335930 215932
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 170254 211924 170260 211988
rect 170324 211986 170330 211988
rect 287697 211986 287763 211989
rect 170324 211984 287763 211986
rect 170324 211928 287702 211984
rect 287758 211928 287763 211984
rect 170324 211926 287763 211928
rect 170324 211924 170330 211926
rect 287697 211923 287763 211926
rect 197118 211788 197124 211852
rect 197188 211850 197194 211852
rect 511993 211850 512059 211853
rect 197188 211848 512059 211850
rect 197188 211792 511998 211848
rect 512054 211792 512059 211848
rect 197188 211790 512059 211792
rect 197188 211788 197194 211790
rect 511993 211787 512059 211790
rect 144126 210428 144132 210492
rect 144196 210490 144202 210492
rect 268326 210490 268332 210492
rect 144196 210430 268332 210490
rect 144196 210428 144202 210430
rect 268326 210428 268332 210430
rect 268396 210428 268402 210492
rect 49601 210354 49667 210357
rect 263542 210354 263548 210356
rect 49601 210352 263548 210354
rect 49601 210296 49606 210352
rect 49662 210296 263548 210352
rect 49601 210294 263548 210296
rect 49601 210291 49667 210294
rect 263542 210292 263548 210294
rect 263612 210292 263618 210356
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 167637 204914 167703 204917
rect 273846 204914 273852 204916
rect 167637 204912 273852 204914
rect 167637 204856 167642 204912
rect 167698 204856 273852 204912
rect 167637 204854 273852 204856
rect 167637 204851 167703 204854
rect 273846 204852 273852 204854
rect 273916 204852 273922 204916
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 124806 200636 124812 200700
rect 124876 200698 124882 200700
rect 263726 200698 263732 200700
rect 124876 200638 263732 200698
rect 124876 200636 124882 200638
rect 263726 200636 263732 200638
rect 263796 200636 263802 200700
rect 120717 199338 120783 199341
rect 259494 199338 259500 199340
rect 120717 199336 259500 199338
rect 120717 199280 120722 199336
rect 120778 199280 259500 199336
rect 120717 199278 259500 199280
rect 120717 199275 120783 199278
rect 259494 199276 259500 199278
rect 259564 199276 259570 199340
rect 69054 195196 69060 195260
rect 69124 195258 69130 195260
rect 271873 195258 271939 195261
rect 69124 195256 271939 195258
rect 69124 195200 271878 195256
rect 271934 195200 271939 195256
rect 69124 195198 271939 195200
rect 69124 195196 69130 195198
rect 271873 195195 271939 195198
rect 135989 192674 136055 192677
rect 258574 192674 258580 192676
rect 135989 192672 258580 192674
rect 135989 192616 135994 192672
rect 136050 192616 258580 192672
rect 135989 192614 258580 192616
rect 135989 192611 136055 192614
rect 258574 192612 258580 192614
rect 258644 192612 258650 192676
rect 57513 192538 57579 192541
rect 258390 192538 258396 192540
rect 57513 192536 258396 192538
rect 57513 192480 57518 192536
rect 57574 192480 258396 192536
rect 57513 192478 258396 192480
rect 57513 192475 57579 192478
rect 258390 192476 258396 192478
rect 258460 192476 258466 192540
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect 152406 191116 152412 191180
rect 152476 191178 152482 191180
rect 209129 191178 209195 191181
rect 152476 191176 209195 191178
rect 152476 191120 209134 191176
rect 209190 191120 209195 191176
rect 152476 191118 209195 191120
rect 152476 191116 152482 191118
rect 209129 191115 209195 191118
rect 118601 191042 118667 191045
rect 503662 191042 503668 191044
rect 118601 191040 503668 191042
rect 118601 190984 118606 191040
rect 118662 190984 503668 191040
rect 118601 190982 503668 190984
rect 118601 190979 118667 190982
rect 503662 190980 503668 190982
rect 503732 190980 503738 191044
rect 148409 189682 148475 189685
rect 259678 189682 259684 189684
rect 148409 189680 259684 189682
rect 148409 189624 148414 189680
rect 148470 189624 259684 189680
rect 148409 189622 259684 189624
rect 148409 189619 148475 189622
rect 259678 189620 259684 189622
rect 259748 189620 259754 189684
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 252001 188322 252067 188325
rect 266302 188322 266308 188324
rect 252001 188320 266308 188322
rect 252001 188264 252006 188320
rect 252062 188264 266308 188320
rect 252001 188262 266308 188264
rect 252001 188259 252067 188262
rect 266302 188260 266308 188262
rect 266372 188260 266378 188324
rect 69013 186962 69079 186965
rect 249374 186962 249380 186964
rect 69013 186960 249380 186962
rect 69013 186904 69018 186960
rect 69074 186904 249380 186960
rect 69013 186902 249380 186904
rect 69013 186899 69079 186902
rect 249374 186900 249380 186902
rect 249444 186900 249450 186964
rect 240961 185602 241027 185605
rect 262254 185602 262260 185604
rect 240961 185600 262260 185602
rect 240961 185544 240966 185600
rect 241022 185544 262260 185600
rect 240961 185542 262260 185544
rect 240961 185539 241027 185542
rect 262254 185540 262260 185542
rect 262324 185540 262330 185604
rect 153837 184242 153903 184245
rect 188429 184242 188495 184245
rect 153837 184240 188495 184242
rect 153837 184184 153842 184240
rect 153898 184184 188434 184240
rect 188490 184184 188495 184240
rect 153837 184182 188495 184184
rect 153837 184179 153903 184182
rect 188429 184179 188495 184182
rect 209037 184242 209103 184245
rect 321318 184242 321324 184244
rect 209037 184240 321324 184242
rect 209037 184184 209042 184240
rect 209098 184184 321324 184240
rect 209037 184182 321324 184184
rect 209037 184179 209103 184182
rect 321318 184180 321324 184182
rect 321388 184180 321394 184244
rect 164877 181658 164943 181661
rect 182909 181658 182975 181661
rect 164877 181656 182975 181658
rect 164877 181600 164882 181656
rect 164938 181600 182914 181656
rect 182970 181600 182975 181656
rect 164877 181598 182975 181600
rect 164877 181595 164943 181598
rect 182909 181595 182975 181598
rect 166206 181460 166212 181524
rect 166276 181522 166282 181524
rect 206277 181522 206343 181525
rect 166276 181520 206343 181522
rect 166276 181464 206282 181520
rect 206338 181464 206343 181520
rect 166276 181462 206343 181464
rect 166276 181460 166282 181462
rect 206277 181459 206343 181462
rect 206461 181522 206527 181525
rect 279417 181522 279483 181525
rect 206461 181520 279483 181522
rect 206461 181464 206466 181520
rect 206522 181464 279422 181520
rect 279478 181464 279483 181520
rect 206461 181462 279483 181464
rect 206461 181459 206527 181462
rect 279417 181459 279483 181462
rect 324957 181522 325023 181525
rect 331438 181522 331444 181524
rect 324957 181520 331444 181522
rect 324957 181464 324962 181520
rect 325018 181464 331444 181520
rect 324957 181462 331444 181464
rect 324957 181459 325023 181462
rect 331438 181460 331444 181462
rect 331508 181460 331514 181524
rect 175181 181386 175247 181389
rect 347957 181386 348023 181389
rect 175181 181384 348023 181386
rect 175181 181328 175186 181384
rect 175242 181328 347962 181384
rect 348018 181328 348023 181384
rect 175181 181326 348023 181328
rect 175181 181323 175247 181326
rect 347957 181323 348023 181326
rect 232497 180162 232563 180165
rect 260966 180162 260972 180164
rect 232497 180160 260972 180162
rect 232497 180104 232502 180160
rect 232558 180104 260972 180160
rect 232497 180102 260972 180104
rect 232497 180099 232563 180102
rect 260966 180100 260972 180102
rect 261036 180100 261042 180164
rect 169109 180026 169175 180029
rect 269062 180026 269068 180028
rect 169109 180024 269068 180026
rect 169109 179968 169114 180024
rect 169170 179968 269068 180024
rect 169109 179966 269068 179968
rect 169109 179963 169175 179966
rect 269062 179964 269068 179966
rect 269132 179964 269138 180028
rect 494053 179346 494119 179349
rect 494053 179344 494162 179346
rect 494053 179288 494058 179344
rect 494114 179288 494162 179344
rect 494053 179283 494162 179288
rect 243537 178938 243603 178941
rect 255446 178938 255452 178940
rect 243537 178936 255452 178938
rect 243537 178880 243542 178936
rect 243598 178880 255452 178936
rect 243537 178878 255452 178880
rect 243537 178875 243603 178878
rect 255446 178876 255452 178878
rect 255516 178876 255522 178940
rect 494102 178908 494162 179283
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 240869 178802 240935 178805
rect 256734 178802 256740 178804
rect 240869 178800 256740 178802
rect 240869 178744 240874 178800
rect 240930 178744 256740 178800
rect 240869 178742 256740 178744
rect 240869 178739 240935 178742
rect 256734 178740 256740 178742
rect 256804 178740 256810 178804
rect 214557 178666 214623 178669
rect 262438 178666 262444 178668
rect 214557 178664 262444 178666
rect 214557 178608 214562 178664
rect 214618 178608 262444 178664
rect 214557 178606 262444 178608
rect 214557 178603 214623 178606
rect 262438 178604 262444 178606
rect 262508 178604 262514 178668
rect 416773 178666 416839 178669
rect 493869 178666 493935 178669
rect 502374 178666 502380 178668
rect 416773 178664 420164 178666
rect 416773 178608 416778 178664
rect 416834 178608 420164 178664
rect 416773 178606 420164 178608
rect 493869 178664 502380 178666
rect 493869 178608 493874 178664
rect 493930 178608 502380 178664
rect 493869 178606 502380 178608
rect 416773 178603 416839 178606
rect 493869 178603 493935 178606
rect 502374 178604 502380 178606
rect 502444 178604 502450 178668
rect 166390 178122 166396 178124
rect 113222 178062 166396 178122
rect 113222 177988 113282 178062
rect 166390 178060 166396 178062
rect 166460 178060 166466 178124
rect 308489 178122 308555 178125
rect 316033 178122 316099 178125
rect 316401 178122 316467 178125
rect 308489 178120 316467 178122
rect 308489 178064 308494 178120
rect 308550 178064 316038 178120
rect 316094 178064 316406 178120
rect 316462 178064 316467 178120
rect 308489 178062 316467 178064
rect 308489 178059 308555 178062
rect 316033 178059 316099 178062
rect 316401 178059 316467 178062
rect 113214 177924 113220 177988
rect 113284 177924 113290 177988
rect 496905 177850 496971 177853
rect 494316 177848 496971 177850
rect 494316 177792 496910 177848
rect 496966 177792 496971 177848
rect 494316 177790 496971 177792
rect 496905 177787 496971 177790
rect 100702 177652 100708 177716
rect 100772 177714 100778 177716
rect 102041 177714 102107 177717
rect 105721 177716 105787 177717
rect 105670 177714 105676 177716
rect 100772 177712 102107 177714
rect 100772 177656 102046 177712
rect 102102 177656 102107 177712
rect 100772 177654 102107 177656
rect 105630 177654 105676 177714
rect 105740 177712 105787 177716
rect 105782 177656 105787 177712
rect 100772 177652 100778 177654
rect 102041 177651 102107 177654
rect 105670 177652 105676 177654
rect 105740 177652 105787 177656
rect 106958 177652 106964 177716
rect 107028 177714 107034 177716
rect 107561 177714 107627 177717
rect 110689 177716 110755 177717
rect 116945 177716 117011 177717
rect 110638 177714 110644 177716
rect 107028 177712 107627 177714
rect 107028 177656 107566 177712
rect 107622 177656 107627 177712
rect 107028 177654 107627 177656
rect 110598 177654 110644 177714
rect 110708 177712 110755 177716
rect 116894 177714 116900 177716
rect 110750 177656 110755 177712
rect 107028 177652 107034 177654
rect 105721 177651 105787 177652
rect 107561 177651 107627 177654
rect 110638 177652 110644 177654
rect 110708 177652 110755 177656
rect 116854 177654 116900 177714
rect 116964 177712 117011 177716
rect 117006 177656 117011 177712
rect 116894 177652 116900 177654
rect 116964 177652 117011 177656
rect 119470 177652 119476 177716
rect 119540 177714 119546 177716
rect 119705 177714 119771 177717
rect 119540 177712 119771 177714
rect 119540 177656 119710 177712
rect 119766 177656 119771 177712
rect 119540 177654 119771 177656
rect 119540 177652 119546 177654
rect 110689 177651 110755 177652
rect 116945 177651 117011 177652
rect 119705 177651 119771 177654
rect 120758 177652 120764 177716
rect 120828 177714 120834 177716
rect 121177 177714 121243 177717
rect 120828 177712 121243 177714
rect 120828 177656 121182 177712
rect 121238 177656 121243 177712
rect 120828 177654 121243 177656
rect 120828 177652 120834 177654
rect 121177 177651 121243 177654
rect 123150 177652 123156 177716
rect 123220 177714 123226 177716
rect 123293 177714 123359 177717
rect 123220 177712 123359 177714
rect 123220 177656 123298 177712
rect 123354 177656 123359 177712
rect 123220 177654 123359 177656
rect 123220 177652 123226 177654
rect 123293 177651 123359 177654
rect 127014 177652 127020 177716
rect 127084 177714 127090 177716
rect 128261 177714 128327 177717
rect 129457 177716 129523 177717
rect 129406 177714 129412 177716
rect 127084 177712 128327 177714
rect 127084 177656 128266 177712
rect 128322 177656 128327 177712
rect 127084 177654 128327 177656
rect 129366 177654 129412 177714
rect 129476 177712 129523 177716
rect 129518 177656 129523 177712
rect 127084 177652 127090 177654
rect 128261 177651 128327 177654
rect 129406 177652 129412 177654
rect 129476 177652 129523 177656
rect 130694 177652 130700 177716
rect 130764 177714 130770 177716
rect 130929 177714 130995 177717
rect 132401 177716 132467 177717
rect 132350 177714 132356 177716
rect 130764 177712 130995 177714
rect 130764 177656 130934 177712
rect 130990 177656 130995 177712
rect 130764 177654 130995 177656
rect 132310 177654 132356 177714
rect 132420 177712 132467 177716
rect 132462 177656 132467 177712
rect 130764 177652 130770 177654
rect 129457 177651 129523 177652
rect 130929 177651 130995 177654
rect 132350 177652 132356 177654
rect 132420 177652 132467 177656
rect 132401 177651 132467 177652
rect 159449 177442 159515 177445
rect 187049 177442 187115 177445
rect 159449 177440 187115 177442
rect 159449 177384 159454 177440
rect 159510 177384 187054 177440
rect 187110 177384 187115 177440
rect 159449 177382 187115 177384
rect 159449 177379 159515 177382
rect 187049 177379 187115 177382
rect 198089 177442 198155 177445
rect 321686 177442 321692 177444
rect 198089 177440 321692 177442
rect 198089 177384 198094 177440
rect 198150 177384 321692 177440
rect 198089 177382 321692 177384
rect 198089 177379 198155 177382
rect 321686 177380 321692 177382
rect 321756 177380 321762 177444
rect 170581 177306 170647 177309
rect 345105 177306 345171 177309
rect 170581 177304 345171 177306
rect 170581 177248 170586 177304
rect 170642 177248 345110 177304
rect 345166 177248 345171 177304
rect 170581 177246 345171 177248
rect 170581 177243 170647 177246
rect 345105 177243 345171 177246
rect 115841 177172 115907 177173
rect 104566 177108 104572 177172
rect 104636 177170 104642 177172
rect 115790 177170 115796 177172
rect 104636 177110 113190 177170
rect 115750 177110 115796 177170
rect 115860 177168 115907 177172
rect 115902 177112 115907 177168
rect 104636 177108 104642 177110
rect 109534 176972 109540 177036
rect 109604 177034 109610 177036
rect 109953 177034 110019 177037
rect 109604 177032 110019 177034
rect 109604 176976 109958 177032
rect 110014 176976 110019 177032
rect 109604 176974 110019 176976
rect 113130 177034 113190 177110
rect 115790 177108 115796 177110
rect 115860 177108 115907 177112
rect 125726 177108 125732 177172
rect 125796 177170 125802 177172
rect 126053 177170 126119 177173
rect 125796 177168 126119 177170
rect 125796 177112 126058 177168
rect 126114 177112 126119 177168
rect 125796 177110 126119 177112
rect 125796 177108 125802 177110
rect 115841 177107 115907 177108
rect 126053 177107 126119 177110
rect 134374 177108 134380 177172
rect 134444 177170 134450 177172
rect 134701 177170 134767 177173
rect 134444 177168 134767 177170
rect 134444 177112 134706 177168
rect 134762 177112 134767 177168
rect 134444 177110 134767 177112
rect 134444 177108 134450 177110
rect 134701 177107 134767 177110
rect 167729 177034 167795 177037
rect 113130 177032 167795 177034
rect 113130 176976 167734 177032
rect 167790 176976 167795 177032
rect 113130 176974 167795 176976
rect 109604 176972 109610 176974
rect 109953 176971 110019 176974
rect 167729 176971 167795 176974
rect 416773 177034 416839 177037
rect 416773 177032 420164 177034
rect 416773 176976 416778 177032
rect 416834 176976 420164 177032
rect 416773 176974 420164 176976
rect 416773 176971 416839 176974
rect 166206 176898 166212 176900
rect 103470 176838 166212 176898
rect 97022 176700 97028 176764
rect 97092 176762 97098 176764
rect 97809 176762 97875 176765
rect 100661 176762 100727 176765
rect 103470 176762 103530 176838
rect 166206 176836 166212 176838
rect 166276 176836 166282 176900
rect 108113 176764 108179 176765
rect 108062 176762 108068 176764
rect 97092 176760 97875 176762
rect 97092 176704 97814 176760
rect 97870 176704 97875 176760
rect 97092 176702 97875 176704
rect 97092 176700 97098 176702
rect 97809 176699 97875 176702
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 103286 176702 103530 176762
rect 108022 176702 108068 176762
rect 108132 176760 108179 176764
rect 108174 176704 108179 176760
rect 103286 176492 103346 176702
rect 108062 176700 108068 176702
rect 108132 176700 108179 176704
rect 112110 176700 112116 176764
rect 112180 176762 112186 176764
rect 112253 176762 112319 176765
rect 114369 176764 114435 176765
rect 124489 176764 124555 176765
rect 114318 176762 114324 176764
rect 112180 176760 112319 176762
rect 112180 176704 112258 176760
rect 112314 176704 112319 176760
rect 112180 176702 112319 176704
rect 114278 176702 114324 176762
rect 114388 176760 114435 176764
rect 124438 176762 124444 176764
rect 114430 176704 114435 176760
rect 112180 176700 112186 176702
rect 108113 176699 108179 176700
rect 112253 176699 112319 176702
rect 114318 176700 114324 176702
rect 114388 176700 114435 176704
rect 124398 176702 124444 176762
rect 124508 176760 124555 176764
rect 128169 176762 128235 176765
rect 133137 176764 133203 176765
rect 136081 176764 136147 176765
rect 148225 176764 148291 176765
rect 158897 176764 158963 176765
rect 133086 176762 133092 176764
rect 124550 176704 124555 176760
rect 124438 176700 124444 176702
rect 124508 176700 124555 176704
rect 114369 176699 114435 176700
rect 124489 176699 124555 176700
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 133046 176702 133092 176762
rect 133156 176760 133203 176764
rect 136030 176762 136036 176764
rect 133198 176704 133203 176760
rect 133086 176700 133092 176702
rect 133156 176700 133203 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 148174 176762 148180 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 148134 176702 148180 176762
rect 148244 176760 148291 176764
rect 158846 176762 158852 176764
rect 148286 176704 148291 176760
rect 148174 176700 148180 176702
rect 148244 176700 148291 176704
rect 158806 176702 158852 176762
rect 158916 176760 158963 176764
rect 496813 176762 496879 176765
rect 158958 176704 158963 176760
rect 158846 176700 158852 176702
rect 158916 176700 158963 176704
rect 494316 176760 496879 176762
rect 494316 176704 496818 176760
rect 496874 176704 496879 176760
rect 494316 176702 496879 176704
rect 133137 176699 133203 176700
rect 136081 176699 136147 176700
rect 148225 176699 148291 176700
rect 158897 176699 158963 176700
rect 496813 176699 496879 176702
rect 128126 176492 128186 176699
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 213913 176218 213979 176221
rect 318609 176218 318675 176221
rect 324589 176218 324655 176221
rect 213913 176216 217242 176218
rect 213913 176160 213918 176216
rect 213974 176160 217242 176216
rect 213913 176158 217242 176160
rect 213913 176155 213979 176158
rect -960 175796 480 176036
rect 160829 175946 160895 175949
rect 166942 175946 166948 175948
rect 160829 175944 166948 175946
rect 160829 175888 160834 175944
rect 160890 175888 166948 175944
rect 160829 175886 166948 175888
rect 160829 175883 160895 175886
rect 166942 175884 166948 175886
rect 167012 175884 167018 175948
rect 217182 175644 217242 176158
rect 318609 176216 324655 176218
rect 318609 176160 318614 176216
rect 318670 176160 324594 176216
rect 324650 176160 324655 176216
rect 318609 176158 324655 176160
rect 318609 176155 318675 176158
rect 324589 176155 324655 176158
rect 245101 176082 245167 176085
rect 259637 176082 259703 176085
rect 245101 176080 259703 176082
rect 245101 176024 245106 176080
rect 245162 176024 259642 176080
rect 259698 176024 259703 176080
rect 245101 176022 259703 176024
rect 245101 176019 245167 176022
rect 259637 176019 259703 176022
rect 321461 176082 321527 176085
rect 321461 176080 321570 176082
rect 321461 176024 321466 176080
rect 321522 176024 321570 176080
rect 321461 176019 321570 176024
rect 224217 175946 224283 175949
rect 249190 175946 249196 175948
rect 224217 175944 249196 175946
rect 224217 175888 224222 175944
rect 224278 175888 249196 175944
rect 224217 175886 249196 175888
rect 224217 175883 224283 175886
rect 249190 175884 249196 175886
rect 249260 175884 249266 175948
rect 248045 175810 248111 175813
rect 248045 175808 248338 175810
rect 248045 175752 248050 175808
rect 248106 175752 248338 175808
rect 248045 175750 248338 175752
rect 248045 175747 248111 175750
rect 248278 175644 248338 175750
rect 320214 175748 320220 175812
rect 320284 175810 320290 175812
rect 321369 175810 321435 175813
rect 320284 175808 321435 175810
rect 320284 175752 321374 175808
rect 321430 175752 321435 175808
rect 320284 175750 321435 175752
rect 320284 175748 320290 175750
rect 321369 175747 321435 175750
rect 306966 175612 306972 175676
rect 307036 175674 307042 175676
rect 307036 175614 310132 175674
rect 307036 175612 307042 175614
rect 321510 175508 321570 176019
rect 496813 175674 496879 175677
rect 494316 175672 496879 175674
rect 494316 175616 496818 175672
rect 496874 175616 496879 175672
rect 494316 175614 496879 175616
rect 496813 175611 496879 175614
rect 98361 175404 98427 175405
rect 102041 175404 102107 175405
rect 118417 175404 118483 175405
rect 121913 175404 121979 175405
rect 98310 175402 98316 175404
rect 98270 175342 98316 175402
rect 98380 175400 98427 175404
rect 101990 175402 101996 175404
rect 98422 175344 98427 175400
rect 98310 175340 98316 175342
rect 98380 175340 98427 175344
rect 101950 175342 101996 175402
rect 102060 175400 102107 175404
rect 118366 175402 118372 175404
rect 102102 175344 102107 175400
rect 101990 175340 101996 175342
rect 102060 175340 102107 175344
rect 118326 175342 118372 175402
rect 118436 175400 118483 175404
rect 121862 175402 121868 175404
rect 118478 175344 118483 175400
rect 118366 175340 118372 175342
rect 118436 175340 118483 175344
rect 121822 175342 121868 175402
rect 121932 175400 121979 175404
rect 121974 175344 121979 175400
rect 121862 175340 121868 175342
rect 121932 175340 121979 175344
rect 98361 175339 98427 175340
rect 102041 175339 102107 175340
rect 118417 175339 118483 175340
rect 121913 175339 121979 175340
rect 249149 175266 249215 175269
rect 248952 175264 249215 175266
rect 248952 175208 249154 175264
rect 249210 175208 249215 175264
rect 248952 175206 249215 175208
rect 249149 175203 249215 175206
rect 307385 175266 307451 175269
rect 416773 175266 416839 175269
rect 307385 175264 310040 175266
rect 307385 175208 307390 175264
rect 307446 175208 310040 175264
rect 307385 175206 310040 175208
rect 416773 175264 420164 175266
rect 416773 175208 416778 175264
rect 416834 175208 420164 175264
rect 416773 175206 420164 175208
rect 307385 175203 307451 175206
rect 416773 175203 416839 175206
rect 213913 175130 213979 175133
rect 213913 175128 217242 175130
rect 213913 175072 213918 175128
rect 213974 175072 217242 175128
rect 213913 175070 217242 175072
rect 213913 175067 213979 175070
rect 217182 174964 217242 175070
rect 307569 174858 307635 174861
rect 307569 174856 310040 174858
rect 307569 174800 307574 174856
rect 307630 174800 310040 174856
rect 307569 174798 310040 174800
rect 307569 174795 307635 174798
rect 214005 174722 214071 174725
rect 252461 174722 252527 174725
rect 323209 174722 323275 174725
rect 214005 174720 217242 174722
rect 214005 174664 214010 174720
rect 214066 174664 217242 174720
rect 214005 174662 217242 174664
rect 248952 174720 252527 174722
rect 248952 174664 252466 174720
rect 252522 174664 252527 174720
rect 248952 174662 252527 174664
rect 321908 174720 323275 174722
rect 321908 174664 323214 174720
rect 323270 174664 323275 174720
rect 321908 174662 323275 174664
rect 214005 174659 214071 174662
rect 217182 174284 217242 174662
rect 252461 174659 252527 174662
rect 323209 174659 323275 174662
rect 307477 174450 307543 174453
rect 496854 174450 496860 174452
rect 307477 174448 310040 174450
rect 307477 174392 307482 174448
rect 307538 174392 310040 174448
rect 307477 174390 310040 174392
rect 494316 174390 496860 174450
rect 307477 174387 307543 174390
rect 496854 174388 496860 174390
rect 496924 174388 496930 174452
rect 249374 174314 249380 174316
rect 248952 174254 249380 174314
rect 249374 174252 249380 174254
rect 249444 174252 249450 174316
rect 307661 174042 307727 174045
rect 324405 174042 324471 174045
rect 307661 174040 310040 174042
rect 307661 173984 307666 174040
rect 307722 173984 310040 174040
rect 307661 173982 310040 173984
rect 321908 174040 324471 174042
rect 321908 173984 324410 174040
rect 324466 173984 324471 174040
rect 321908 173982 324471 173984
rect 307661 173979 307727 173982
rect 324405 173979 324471 173982
rect 213913 173770 213979 173773
rect 252461 173770 252527 173773
rect 321369 173770 321435 173773
rect 213913 173768 217242 173770
rect 213913 173712 213918 173768
rect 213974 173712 217242 173768
rect 213913 173710 217242 173712
rect 248952 173768 252527 173770
rect 248952 173712 252466 173768
rect 252522 173712 252527 173768
rect 248952 173710 252527 173712
rect 213913 173707 213979 173710
rect 217182 173604 217242 173710
rect 252461 173707 252527 173710
rect 321326 173768 321435 173770
rect 321326 173712 321374 173768
rect 321430 173712 321435 173768
rect 321326 173707 321435 173712
rect 307293 173634 307359 173637
rect 307293 173632 310040 173634
rect 307293 173576 307298 173632
rect 307354 173576 310040 173632
rect 307293 173574 310040 173576
rect 307293 173571 307359 173574
rect 214005 173362 214071 173365
rect 249190 173362 249196 173364
rect 214005 173360 217242 173362
rect 214005 173304 214010 173360
rect 214066 173304 217242 173360
rect 214005 173302 217242 173304
rect 248952 173302 249196 173362
rect 214005 173299 214071 173302
rect 217182 172924 217242 173302
rect 249190 173300 249196 173302
rect 249260 173300 249266 173364
rect 307477 173226 307543 173229
rect 307477 173224 310040 173226
rect 307477 173168 307482 173224
rect 307538 173168 310040 173224
rect 321326 173196 321386 173707
rect 307477 173166 310040 173168
rect 307477 173163 307543 173166
rect 249241 172818 249307 172821
rect 248952 172816 249307 172818
rect 248952 172760 249246 172816
rect 249302 172760 249307 172816
rect 248952 172758 249307 172760
rect 249241 172755 249307 172758
rect 307661 172682 307727 172685
rect 321829 172682 321895 172685
rect 307661 172680 310040 172682
rect 307661 172624 307666 172680
rect 307722 172624 310040 172680
rect 307661 172622 310040 172624
rect 321829 172680 321938 172682
rect 321829 172624 321834 172680
rect 321890 172624 321938 172680
rect 307661 172619 307727 172622
rect 321829 172619 321938 172624
rect 213913 172410 213979 172413
rect 252461 172410 252527 172413
rect 213913 172408 217242 172410
rect 213913 172352 213918 172408
rect 213974 172352 217242 172408
rect 213913 172350 217242 172352
rect 248952 172408 252527 172410
rect 248952 172352 252466 172408
rect 252522 172352 252527 172408
rect 321878 172380 321938 172619
rect 334566 172484 334572 172548
rect 334636 172546 334642 172548
rect 420134 172546 420194 173604
rect 495525 173362 495591 173365
rect 494316 173360 495591 173362
rect 494316 173304 495530 173360
rect 495586 173304 495591 173360
rect 494316 173302 495591 173304
rect 495525 173299 495591 173302
rect 334636 172486 420194 172546
rect 334636 172484 334642 172486
rect 248952 172350 252527 172352
rect 213913 172347 213979 172350
rect 217182 172244 217242 172350
rect 252461 172347 252527 172350
rect 306741 172274 306807 172277
rect 495934 172274 495940 172276
rect 306741 172272 310040 172274
rect 306741 172216 306746 172272
rect 306802 172216 310040 172272
rect 306741 172214 310040 172216
rect 494316 172214 495940 172274
rect 306741 172211 306807 172214
rect 495934 172212 495940 172214
rect 496004 172212 496010 172276
rect 214097 172002 214163 172005
rect 214097 172000 217242 172002
rect 214097 171944 214102 172000
rect 214158 171944 217242 172000
rect 214097 171942 217242 171944
rect 214097 171939 214163 171942
rect 167637 171594 167703 171597
rect 164694 171592 167703 171594
rect 164694 171536 167642 171592
rect 167698 171536 167703 171592
rect 217182 171564 217242 171942
rect 252369 171866 252435 171869
rect 248952 171864 252435 171866
rect 248952 171808 252374 171864
rect 252430 171808 252435 171864
rect 248952 171806 252435 171808
rect 252369 171803 252435 171806
rect 307109 171866 307175 171869
rect 416773 171866 416839 171869
rect 307109 171864 310040 171866
rect 307109 171808 307114 171864
rect 307170 171808 310040 171864
rect 307109 171806 310040 171808
rect 416773 171864 420164 171866
rect 416773 171808 416778 171864
rect 416834 171808 420164 171864
rect 416773 171806 420164 171808
rect 307109 171803 307175 171806
rect 416773 171803 416839 171806
rect 164694 171534 167703 171536
rect 167637 171531 167703 171534
rect 249333 171458 249399 171461
rect 248952 171456 249399 171458
rect 248952 171400 249338 171456
rect 249394 171400 249399 171456
rect 248952 171398 249399 171400
rect 249333 171395 249399 171398
rect 307661 171458 307727 171461
rect 307661 171456 310040 171458
rect 307661 171400 307666 171456
rect 307722 171400 310040 171456
rect 307661 171398 310040 171400
rect 307661 171395 307727 171398
rect 321878 171186 321938 171700
rect 331438 171186 331444 171188
rect 216998 171126 217242 171186
rect 321878 171126 331444 171186
rect 213913 171050 213979 171053
rect 216998 171050 217058 171126
rect 213913 171048 217058 171050
rect 213913 170992 213918 171048
rect 213974 170992 217058 171048
rect 217182 171020 217242 171126
rect 331438 171124 331444 171126
rect 331508 171124 331514 171188
rect 498101 171186 498167 171189
rect 494316 171184 498167 171186
rect 494316 171128 498106 171184
rect 498162 171128 498167 171184
rect 494316 171126 498167 171128
rect 498101 171123 498167 171126
rect 306741 171050 306807 171053
rect 306741 171048 310040 171050
rect 213913 170990 217058 170992
rect 306741 170992 306746 171048
rect 306802 170992 310040 171048
rect 306741 170990 310040 170992
rect 213913 170987 213979 170990
rect 306741 170987 306807 170990
rect 252461 170914 252527 170917
rect 324589 170914 324655 170917
rect 248952 170912 252527 170914
rect 248952 170856 252466 170912
rect 252522 170856 252527 170912
rect 248952 170854 252527 170856
rect 321908 170912 324655 170914
rect 321908 170856 324594 170912
rect 324650 170856 324655 170912
rect 321908 170854 324655 170856
rect 252461 170851 252527 170854
rect 324589 170851 324655 170854
rect 214005 170778 214071 170781
rect 214005 170776 217242 170778
rect 214005 170720 214010 170776
rect 214066 170720 217242 170776
rect 214005 170718 217242 170720
rect 214005 170715 214071 170718
rect 217182 170340 217242 170718
rect 306925 170642 306991 170645
rect 306925 170640 310040 170642
rect 306925 170584 306930 170640
rect 306986 170584 310040 170640
rect 306925 170582 310040 170584
rect 306925 170579 306991 170582
rect 321318 170580 321324 170644
rect 321388 170580 321394 170644
rect 252369 170506 252435 170509
rect 248952 170504 252435 170506
rect 248952 170448 252374 170504
rect 252430 170448 252435 170504
rect 248952 170446 252435 170448
rect 252369 170443 252435 170446
rect 307661 170234 307727 170237
rect 307661 170232 310040 170234
rect 307661 170176 307666 170232
rect 307722 170176 310040 170232
rect 307661 170174 310040 170176
rect 307661 170171 307727 170174
rect 252461 170098 252527 170101
rect 248952 170096 252527 170098
rect 248952 170040 252466 170096
rect 252522 170040 252527 170096
rect 321326 170068 321386 170580
rect 248952 170038 252527 170040
rect 252461 170035 252527 170038
rect 307477 169826 307543 169829
rect 216998 169766 217242 169826
rect 214925 169690 214991 169693
rect 216998 169690 217058 169766
rect 214925 169688 217058 169690
rect 214925 169632 214930 169688
rect 214986 169632 217058 169688
rect 217182 169660 217242 169766
rect 307477 169824 310040 169826
rect 307477 169768 307482 169824
rect 307538 169768 310040 169824
rect 307477 169766 310040 169768
rect 307477 169763 307543 169766
rect 336038 169764 336044 169828
rect 336108 169826 336114 169828
rect 420134 169826 420194 170204
rect 494286 169828 494346 169932
rect 336108 169766 420194 169826
rect 336108 169764 336114 169766
rect 494278 169764 494284 169828
rect 494348 169764 494354 169828
rect 321277 169690 321343 169693
rect 321277 169688 321386 169690
rect 214925 169630 217058 169632
rect 321277 169632 321282 169688
rect 321338 169632 321386 169688
rect 214925 169627 214991 169630
rect 321277 169627 321386 169632
rect 250253 169554 250319 169557
rect 248952 169552 250319 169554
rect 248952 169496 250258 169552
rect 250314 169496 250319 169552
rect 248952 169494 250319 169496
rect 250253 169491 250319 169494
rect 214649 169418 214715 169421
rect 214649 169416 217242 169418
rect 214649 169360 214654 169416
rect 214710 169360 217242 169416
rect 321326 169388 321386 169627
rect 214649 169358 217242 169360
rect 214649 169355 214715 169358
rect 217182 168980 217242 169358
rect 307569 169282 307635 169285
rect 307569 169280 310040 169282
rect 307569 169224 307574 169280
rect 307630 169224 310040 169280
rect 307569 169222 310040 169224
rect 307569 169219 307635 169222
rect 252829 169146 252895 169149
rect 248952 169144 252895 169146
rect 248952 169088 252834 169144
rect 252890 169088 252895 169144
rect 248952 169086 252895 169088
rect 252829 169083 252895 169086
rect 306557 168874 306623 168877
rect 306557 168872 310040 168874
rect 306557 168816 306562 168872
rect 306618 168816 310040 168872
rect 306557 168814 310040 168816
rect 306557 168811 306623 168814
rect 324313 168602 324379 168605
rect 321908 168600 324379 168602
rect 248860 168498 249442 168558
rect 321908 168544 324318 168600
rect 324374 168544 324379 168600
rect 321908 168542 324379 168544
rect 324313 168539 324379 168542
rect 249382 168466 249442 168498
rect 494102 168469 494162 168844
rect 258390 168466 258396 168468
rect 216998 168406 217242 168466
rect 249382 168406 258396 168466
rect 213913 168330 213979 168333
rect 216998 168330 217058 168406
rect 213913 168328 217058 168330
rect 213913 168272 213918 168328
rect 213974 168272 217058 168328
rect 217182 168300 217242 168406
rect 258390 168404 258396 168406
rect 258460 168404 258466 168468
rect 307661 168466 307727 168469
rect 416773 168466 416839 168469
rect 307661 168464 310040 168466
rect 307661 168408 307666 168464
rect 307722 168408 310040 168464
rect 307661 168406 310040 168408
rect 416773 168464 420164 168466
rect 416773 168408 416778 168464
rect 416834 168408 420164 168464
rect 416773 168406 420164 168408
rect 494053 168464 494162 168469
rect 494053 168408 494058 168464
rect 494114 168408 494162 168464
rect 494053 168406 494162 168408
rect 307661 168403 307727 168406
rect 416773 168403 416839 168406
rect 494053 168403 494119 168406
rect 213913 168270 217058 168272
rect 213913 168267 213979 168270
rect 252461 168194 252527 168197
rect 248952 168192 252527 168194
rect 248952 168136 252466 168192
rect 252522 168136 252527 168192
rect 248952 168134 252527 168136
rect 252461 168131 252527 168134
rect 214005 168058 214071 168061
rect 307293 168058 307359 168061
rect 214005 168056 217242 168058
rect 214005 168000 214010 168056
rect 214066 168000 217242 168056
rect 214005 167998 217242 168000
rect 214005 167995 214071 167998
rect 217182 167620 217242 167998
rect 307293 168056 310040 168058
rect 307293 168000 307298 168056
rect 307354 168000 310040 168056
rect 307293 167998 310040 168000
rect 307293 167995 307359 167998
rect 324313 167786 324379 167789
rect 496813 167786 496879 167789
rect 321908 167784 324379 167786
rect 321908 167728 324318 167784
rect 324374 167728 324379 167784
rect 321908 167726 324379 167728
rect 494316 167784 496879 167786
rect 494316 167728 496818 167784
rect 496874 167728 496879 167784
rect 494316 167726 496879 167728
rect 324313 167723 324379 167726
rect 496813 167723 496879 167726
rect 307569 167650 307635 167653
rect 307569 167648 310040 167650
rect 248860 167546 249442 167606
rect 307569 167592 307574 167648
rect 307630 167592 310040 167648
rect 307569 167590 310040 167592
rect 307569 167587 307635 167590
rect 249382 167378 249442 167546
rect 260966 167378 260972 167380
rect 249382 167318 260972 167378
rect 260966 167316 260972 167318
rect 261036 167316 261042 167380
rect 252369 167242 252435 167245
rect 248952 167240 252435 167242
rect 248952 167184 252374 167240
rect 252430 167184 252435 167240
rect 248952 167182 252435 167184
rect 252369 167179 252435 167182
rect 307661 167242 307727 167245
rect 307661 167240 310040 167242
rect 307661 167184 307666 167240
rect 307722 167184 310040 167240
rect 307661 167182 310040 167184
rect 307661 167179 307727 167182
rect 349102 167106 349108 167108
rect 321908 167046 349108 167106
rect 349102 167044 349108 167046
rect 349172 167044 349178 167108
rect 213913 166970 213979 166973
rect 216998 166970 217242 167010
rect 213913 166968 217242 166970
rect 213913 166912 213918 166968
rect 213974 166950 217242 166968
rect 213974 166912 217058 166950
rect 217182 166940 217242 166950
rect 213913 166910 217058 166912
rect 213913 166907 213979 166910
rect 503662 166908 503668 166972
rect 503732 166970 503738 166972
rect 504081 166970 504147 166973
rect 503732 166968 504147 166970
rect 503732 166912 504086 166968
rect 504142 166912 504147 166968
rect 503732 166910 504147 166912
rect 503732 166908 503738 166910
rect 504081 166907 504147 166910
rect 306741 166834 306807 166837
rect 306741 166832 310040 166834
rect 306741 166776 306746 166832
rect 306802 166776 310040 166832
rect 306741 166774 310040 166776
rect 306741 166771 306807 166774
rect 321686 166772 321692 166836
rect 321756 166772 321762 166836
rect 416773 166834 416839 166837
rect 416773 166832 420164 166834
rect 416773 166776 416778 166832
rect 416834 166776 420164 166832
rect 416773 166774 420164 166776
rect 214097 166698 214163 166701
rect 252461 166698 252527 166701
rect 214097 166696 217242 166698
rect 214097 166640 214102 166696
rect 214158 166640 217242 166696
rect 214097 166638 217242 166640
rect 248952 166696 252527 166698
rect 248952 166640 252466 166696
rect 252522 166640 252527 166696
rect 248952 166638 252527 166640
rect 214097 166635 214163 166638
rect 217182 166396 217242 166638
rect 252461 166635 252527 166638
rect 306557 166426 306623 166429
rect 306557 166424 310040 166426
rect 306557 166368 306562 166424
rect 306618 166368 310040 166424
rect 306557 166366 310040 166368
rect 306557 166363 306623 166366
rect 252369 166290 252435 166293
rect 248952 166288 252435 166290
rect 248952 166232 252374 166288
rect 252430 166232 252435 166288
rect 321694 166260 321754 166772
rect 416773 166771 416839 166774
rect 496813 166698 496879 166701
rect 494316 166696 496879 166698
rect 494316 166640 496818 166696
rect 496874 166640 496879 166696
rect 494316 166638 496879 166640
rect 496813 166635 496879 166638
rect 248952 166230 252435 166232
rect 252369 166227 252435 166230
rect 214005 166154 214071 166157
rect 214005 166152 217242 166154
rect 214005 166096 214010 166152
rect 214066 166096 217242 166152
rect 214005 166094 217242 166096
rect 214005 166091 214071 166094
rect 217182 165716 217242 166094
rect 307477 165882 307543 165885
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 307477 165880 310040 165882
rect 307477 165824 307482 165880
rect 307538 165824 310040 165880
rect 307477 165822 310040 165824
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 307477 165819 307543 165822
rect 580165 165819 580231 165822
rect 252461 165746 252527 165749
rect 248952 165744 252527 165746
rect 248952 165688 252466 165744
rect 252522 165688 252527 165744
rect 583520 165732 584960 165822
rect 248952 165686 252527 165688
rect 252461 165683 252527 165686
rect 307201 165474 307267 165477
rect 324313 165474 324379 165477
rect 496813 165474 496879 165477
rect 307201 165472 310040 165474
rect 307201 165416 307206 165472
rect 307262 165416 310040 165472
rect 307201 165414 310040 165416
rect 321908 165472 324379 165474
rect 321908 165416 324318 165472
rect 324374 165416 324379 165472
rect 321908 165414 324379 165416
rect 494316 165472 496879 165474
rect 494316 165416 496818 165472
rect 496874 165416 496879 165472
rect 494316 165414 496879 165416
rect 307201 165411 307267 165414
rect 324313 165411 324379 165414
rect 496813 165411 496879 165414
rect 213913 165338 213979 165341
rect 252461 165338 252527 165341
rect 213913 165336 217242 165338
rect 213913 165280 213918 165336
rect 213974 165280 217242 165336
rect 213913 165278 217242 165280
rect 248952 165336 252527 165338
rect 248952 165280 252466 165336
rect 252522 165280 252527 165336
rect 248952 165278 252527 165280
rect 213913 165275 213979 165278
rect 217182 165036 217242 165278
rect 252461 165275 252527 165278
rect 307017 165066 307083 165069
rect 416773 165066 416839 165069
rect 307017 165064 310040 165066
rect 307017 165008 307022 165064
rect 307078 165008 310040 165064
rect 307017 165006 310040 165008
rect 416773 165064 420164 165066
rect 416773 165008 416778 165064
rect 416834 165008 420164 165064
rect 416773 165006 420164 165008
rect 307017 165003 307083 165006
rect 416773 165003 416839 165006
rect 214005 164794 214071 164797
rect 252369 164794 252435 164797
rect 324405 164794 324471 164797
rect 214005 164792 217242 164794
rect 214005 164736 214010 164792
rect 214066 164736 217242 164792
rect 214005 164734 217242 164736
rect 248952 164792 252435 164794
rect 248952 164736 252374 164792
rect 252430 164736 252435 164792
rect 248952 164734 252435 164736
rect 321908 164792 324471 164794
rect 321908 164736 324410 164792
rect 324466 164736 324471 164792
rect 321908 164734 324471 164736
rect 214005 164731 214071 164734
rect 217182 164356 217242 164734
rect 252369 164731 252435 164734
rect 324405 164731 324471 164734
rect 307661 164658 307727 164661
rect 307661 164656 310040 164658
rect 307661 164600 307666 164656
rect 307722 164600 310040 164656
rect 307661 164598 310040 164600
rect 307661 164595 307727 164598
rect 252737 164386 252803 164389
rect 495709 164386 495775 164389
rect 496353 164386 496419 164389
rect 248952 164384 252803 164386
rect 248952 164328 252742 164384
rect 252798 164328 252803 164384
rect 248952 164326 252803 164328
rect 494316 164384 496419 164386
rect 494316 164328 495714 164384
rect 495770 164328 496358 164384
rect 496414 164328 496419 164384
rect 494316 164326 496419 164328
rect 252737 164323 252803 164326
rect 495709 164323 495775 164326
rect 496353 164323 496419 164326
rect 307109 164250 307175 164253
rect 307109 164248 310040 164250
rect 307109 164192 307114 164248
rect 307170 164192 310040 164248
rect 307109 164190 310040 164192
rect 307109 164187 307175 164190
rect 252461 163978 252527 163981
rect 324313 163978 324379 163981
rect 248952 163976 252527 163978
rect 248952 163920 252466 163976
rect 252522 163920 252527 163976
rect 248952 163918 252527 163920
rect 321908 163976 324379 163978
rect 321908 163920 324318 163976
rect 324374 163920 324379 163976
rect 321908 163918 324379 163920
rect 252461 163915 252527 163918
rect 324313 163915 324379 163918
rect 306925 163842 306991 163845
rect 200070 163782 217242 163842
rect 166390 163100 166396 163164
rect 166460 163162 166466 163164
rect 200070 163162 200130 163782
rect 217182 163676 217242 163782
rect 306925 163840 310040 163842
rect 306925 163784 306930 163840
rect 306986 163784 310040 163840
rect 306925 163782 310040 163784
rect 306925 163779 306991 163782
rect 213913 163434 213979 163437
rect 307385 163434 307451 163437
rect 416773 163434 416839 163437
rect 213913 163432 217426 163434
rect 213913 163376 213918 163432
rect 213974 163376 217426 163432
rect 307385 163432 310040 163434
rect 213913 163374 217426 163376
rect 213913 163371 213979 163374
rect 166460 163102 200130 163162
rect 166460 163100 166466 163102
rect 217366 162996 217426 163374
rect 248860 163330 249442 163390
rect 307385 163376 307390 163432
rect 307446 163376 310040 163432
rect 307385 163374 310040 163376
rect 416773 163432 420164 163434
rect 416773 163376 416778 163432
rect 416834 163376 420164 163432
rect 416773 163374 420164 163376
rect 307385 163371 307451 163374
rect 416773 163371 416839 163374
rect 249382 163162 249442 163330
rect 496813 163298 496879 163301
rect 494316 163296 496879 163298
rect 494316 163240 496818 163296
rect 496874 163240 496879 163296
rect 494316 163238 496879 163240
rect 496813 163235 496879 163238
rect 262438 163162 262444 163164
rect 249382 163102 262444 163162
rect 262438 163100 262444 163102
rect 262508 163100 262514 163164
rect 324405 163162 324471 163165
rect 321908 163160 324471 163162
rect 321908 163104 324410 163160
rect 324466 163104 324471 163160
rect 321908 163102 324471 163104
rect 324405 163099 324471 163102
rect 252369 163026 252435 163029
rect 248952 163024 252435 163026
rect -960 162890 480 162980
rect 248952 162968 252374 163024
rect 252430 162968 252435 163024
rect 248952 162966 252435 162968
rect 252369 162963 252435 162966
rect 305637 163026 305703 163029
rect 306925 163026 306991 163029
rect 305637 163024 306991 163026
rect 305637 162968 305642 163024
rect 305698 162968 306930 163024
rect 306986 162968 306991 163024
rect 305637 162966 306991 162968
rect 305637 162963 305703 162966
rect 306925 162963 306991 162966
rect 307661 163026 307727 163029
rect 307661 163024 310040 163026
rect 307661 162968 307666 163024
rect 307722 162968 310040 163024
rect 307661 162966 310040 162968
rect 307661 162963 307727 162966
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 213913 162754 213979 162757
rect 213913 162752 217242 162754
rect 213913 162696 213918 162752
rect 213974 162696 217242 162752
rect 213913 162694 217242 162696
rect 213913 162691 213979 162694
rect 217182 162316 217242 162694
rect 252461 162482 252527 162485
rect 248952 162480 252527 162482
rect 248952 162424 252466 162480
rect 252522 162424 252527 162480
rect 248952 162422 252527 162424
rect 252461 162419 252527 162422
rect 307477 162482 307543 162485
rect 324313 162482 324379 162485
rect 307477 162480 310040 162482
rect 307477 162424 307482 162480
rect 307538 162424 310040 162480
rect 307477 162422 310040 162424
rect 321908 162480 324379 162482
rect 321908 162424 324318 162480
rect 324374 162424 324379 162480
rect 321908 162422 324379 162424
rect 307477 162419 307543 162422
rect 324313 162419 324379 162422
rect 321645 162210 321711 162213
rect 496813 162210 496879 162213
rect 321645 162208 321754 162210
rect 321645 162152 321650 162208
rect 321706 162152 321754 162208
rect 321645 162147 321754 162152
rect 494316 162208 496879 162210
rect 494316 162152 496818 162208
rect 496874 162152 496879 162208
rect 494316 162150 496879 162152
rect 496813 162147 496879 162150
rect 214005 162074 214071 162077
rect 252369 162074 252435 162077
rect 214005 162072 217242 162074
rect 214005 162016 214010 162072
rect 214066 162016 217242 162072
rect 214005 162014 217242 162016
rect 248952 162072 252435 162074
rect 248952 162016 252374 162072
rect 252430 162016 252435 162072
rect 248952 162014 252435 162016
rect 214005 162011 214071 162014
rect 217182 161772 217242 162014
rect 252369 162011 252435 162014
rect 307569 162074 307635 162077
rect 307569 162072 310040 162074
rect 307569 162016 307574 162072
rect 307630 162016 310040 162072
rect 307569 162014 310040 162016
rect 307569 162011 307635 162014
rect 307661 161666 307727 161669
rect 307661 161664 310040 161666
rect 307661 161608 307666 161664
rect 307722 161608 310040 161664
rect 321694 161636 321754 162147
rect 416773 161802 416839 161805
rect 416773 161800 420164 161802
rect 416773 161744 416778 161800
rect 416834 161744 420164 161800
rect 416773 161742 420164 161744
rect 416773 161739 416839 161742
rect 307661 161606 310040 161608
rect 307661 161603 307727 161606
rect 249149 161530 249215 161533
rect 248952 161528 249215 161530
rect 248952 161472 249154 161528
rect 249210 161472 249215 161528
rect 248952 161470 249215 161472
rect 249149 161467 249215 161470
rect 213913 161394 213979 161397
rect 213913 161392 217242 161394
rect 213913 161336 213918 161392
rect 213974 161336 217242 161392
rect 213913 161334 217242 161336
rect 213913 161331 213979 161334
rect 217182 161092 217242 161334
rect 306557 161258 306623 161261
rect 306557 161256 310040 161258
rect 306557 161200 306562 161256
rect 306618 161200 310040 161256
rect 306557 161198 310040 161200
rect 306557 161195 306623 161198
rect 256734 161122 256740 161124
rect 248952 161062 256740 161122
rect 256734 161060 256740 161062
rect 256804 161060 256810 161124
rect 496905 160986 496971 160989
rect 494316 160984 496971 160986
rect 494316 160928 496910 160984
rect 496966 160928 496971 160984
rect 494316 160926 496971 160928
rect 496905 160923 496971 160926
rect 214005 160850 214071 160853
rect 307569 160850 307635 160853
rect 322933 160850 322999 160853
rect 214005 160848 217242 160850
rect 214005 160792 214010 160848
rect 214066 160792 217242 160848
rect 214005 160790 217242 160792
rect 214005 160787 214071 160790
rect 217182 160412 217242 160790
rect 307569 160848 310040 160850
rect 307569 160792 307574 160848
rect 307630 160792 310040 160848
rect 307569 160790 310040 160792
rect 321908 160848 322999 160850
rect 321908 160792 322938 160848
rect 322994 160792 322999 160848
rect 321908 160790 322999 160792
rect 307569 160787 307635 160790
rect 322933 160787 322999 160790
rect 252461 160578 252527 160581
rect 248952 160576 252527 160578
rect 248952 160520 252466 160576
rect 252522 160520 252527 160576
rect 248952 160518 252527 160520
rect 252461 160515 252527 160518
rect 307661 160442 307727 160445
rect 307661 160440 310040 160442
rect 307661 160384 307666 160440
rect 307722 160384 310040 160440
rect 307661 160382 310040 160384
rect 307661 160379 307727 160382
rect 251449 160170 251515 160173
rect 325601 160170 325667 160173
rect 248952 160168 251515 160170
rect 248952 160112 251454 160168
rect 251510 160112 251515 160168
rect 248952 160110 251515 160112
rect 321908 160168 325667 160170
rect 321908 160112 325606 160168
rect 325662 160112 325667 160168
rect 321908 160110 325667 160112
rect 251449 160107 251515 160110
rect 325601 160107 325667 160110
rect 306925 160034 306991 160037
rect 416773 160034 416839 160037
rect 306925 160032 310040 160034
rect 306925 159976 306930 160032
rect 306986 159976 310040 160032
rect 306925 159974 310040 159976
rect 416773 160032 420164 160034
rect 416773 159976 416778 160032
rect 416834 159976 420164 160032
rect 416773 159974 420164 159976
rect 306925 159971 306991 159974
rect 416773 159971 416839 159974
rect 213913 159898 213979 159901
rect 496905 159898 496971 159901
rect 213913 159896 217242 159898
rect 213913 159840 213918 159896
rect 213974 159840 217242 159896
rect 213913 159838 217242 159840
rect 494316 159896 496971 159898
rect 494316 159840 496910 159896
rect 496966 159840 496971 159896
rect 494316 159838 496971 159840
rect 213913 159835 213979 159838
rect 217182 159732 217242 159838
rect 496905 159835 496971 159838
rect 252461 159626 252527 159629
rect 248952 159624 252527 159626
rect 248952 159568 252466 159624
rect 252522 159568 252527 159624
rect 248952 159566 252527 159568
rect 252461 159563 252527 159566
rect 307569 159626 307635 159629
rect 307569 159624 310040 159626
rect 307569 159568 307574 159624
rect 307630 159568 310040 159624
rect 307569 159566 310040 159568
rect 307569 159563 307635 159566
rect 214005 159490 214071 159493
rect 214005 159488 217242 159490
rect 214005 159432 214010 159488
rect 214066 159432 217242 159488
rect 214005 159430 217242 159432
rect 214005 159427 214071 159430
rect 217182 159052 217242 159430
rect 323117 159354 323183 159357
rect 321908 159352 323183 159354
rect 321908 159296 323122 159352
rect 323178 159296 323183 159352
rect 321908 159294 323183 159296
rect 323117 159291 323183 159294
rect 251357 159218 251423 159221
rect 248952 159216 251423 159218
rect 248952 159160 251362 159216
rect 251418 159160 251423 159216
rect 248952 159158 251423 159160
rect 251357 159155 251423 159158
rect 307661 159082 307727 159085
rect 307661 159080 310040 159082
rect 307661 159024 307666 159080
rect 307722 159024 310040 159080
rect 307661 159022 310040 159024
rect 307661 159019 307727 159022
rect 252502 158810 252508 158812
rect 248952 158750 252508 158810
rect 252502 158748 252508 158750
rect 252572 158748 252578 158812
rect 496997 158810 497063 158813
rect 494316 158808 497063 158810
rect 494316 158752 497002 158808
rect 497058 158752 497063 158808
rect 494316 158750 497063 158752
rect 496997 158747 497063 158750
rect 307385 158674 307451 158677
rect 307385 158672 310040 158674
rect 307385 158616 307390 158672
rect 307446 158616 310040 158672
rect 307385 158614 310040 158616
rect 307385 158611 307451 158614
rect 324313 158538 324379 158541
rect 321908 158536 324379 158538
rect 321908 158480 324318 158536
rect 324374 158480 324379 158536
rect 321908 158478 324379 158480
rect 324313 158475 324379 158478
rect 217182 157858 217242 158372
rect 252369 158266 252435 158269
rect 248952 158264 252435 158266
rect 248952 158208 252374 158264
rect 252430 158208 252435 158264
rect 248952 158206 252435 158208
rect 252369 158203 252435 158206
rect 306741 158266 306807 158269
rect 306741 158264 310040 158266
rect 306741 158208 306746 158264
rect 306802 158208 310040 158264
rect 306741 158206 310040 158208
rect 306741 158203 306807 158206
rect 252461 157858 252527 157861
rect 200070 157798 217242 157858
rect 248952 157856 252527 157858
rect 248952 157800 252466 157856
rect 252522 157800 252527 157856
rect 248952 157798 252527 157800
rect 166206 157388 166212 157452
rect 166276 157450 166282 157452
rect 200070 157450 200130 157798
rect 252461 157795 252527 157798
rect 307477 157858 307543 157861
rect 324405 157858 324471 157861
rect 307477 157856 310040 157858
rect 307477 157800 307482 157856
rect 307538 157800 310040 157856
rect 307477 157798 310040 157800
rect 321908 157856 324471 157858
rect 321908 157800 324410 157856
rect 324466 157800 324471 157856
rect 321908 157798 324471 157800
rect 307477 157795 307543 157798
rect 324405 157795 324471 157798
rect 166276 157390 200130 157450
rect 213913 157450 213979 157453
rect 217366 157450 217426 157692
rect 213913 157448 217426 157450
rect 213913 157392 213918 157448
rect 213974 157392 217426 157448
rect 213913 157390 217426 157392
rect 307109 157450 307175 157453
rect 307109 157448 310040 157450
rect 307109 157392 307114 157448
rect 307170 157392 310040 157448
rect 307109 157390 310040 157392
rect 166276 157388 166282 157390
rect 213913 157387 213979 157390
rect 307109 157387 307175 157390
rect 338614 157388 338620 157452
rect 338684 157450 338690 157452
rect 420134 157450 420194 158372
rect 496905 157722 496971 157725
rect 494316 157720 496971 157722
rect 494316 157664 496910 157720
rect 496966 157664 496971 157720
rect 494316 157662 496971 157664
rect 496905 157659 496971 157662
rect 338684 157390 420194 157450
rect 338684 157388 338690 157390
rect 213913 157314 213979 157317
rect 252461 157314 252527 157317
rect 213913 157312 217242 157314
rect 213913 157256 213918 157312
rect 213974 157256 217242 157312
rect 213913 157254 217242 157256
rect 248952 157312 252527 157314
rect 248952 157256 252466 157312
rect 252522 157256 252527 157312
rect 248952 157254 252527 157256
rect 213913 157251 213979 157254
rect 217182 157148 217242 157254
rect 252461 157251 252527 157254
rect 306557 157042 306623 157045
rect 306557 157040 310040 157042
rect 306557 156984 306562 157040
rect 306618 156984 310040 157040
rect 306557 156982 310040 156984
rect 306557 156979 306623 156982
rect 214005 156906 214071 156909
rect 251541 156906 251607 156909
rect 214005 156904 217242 156906
rect 214005 156848 214010 156904
rect 214066 156848 217242 156904
rect 214005 156846 217242 156848
rect 248952 156904 251607 156906
rect 248952 156848 251546 156904
rect 251602 156848 251607 156904
rect 248952 156846 251607 156848
rect 214005 156843 214071 156846
rect 217182 156468 217242 156846
rect 251541 156843 251607 156846
rect 307569 156634 307635 156637
rect 307569 156632 310040 156634
rect 307569 156576 307574 156632
rect 307630 156576 310040 156632
rect 307569 156574 310040 156576
rect 307569 156571 307635 156574
rect 321878 156498 321938 157012
rect 416773 156634 416839 156637
rect 416773 156632 420164 156634
rect 416773 156576 416778 156632
rect 416834 156576 420164 156632
rect 416773 156574 420164 156576
rect 416773 156571 416839 156574
rect 334014 156498 334020 156500
rect 321878 156438 334020 156498
rect 334014 156436 334020 156438
rect 334084 156436 334090 156500
rect 496905 156498 496971 156501
rect 494316 156496 496971 156498
rect 494316 156440 496910 156496
rect 496966 156440 496971 156496
rect 494316 156438 496971 156440
rect 496905 156435 496971 156438
rect 251173 156362 251239 156365
rect 324313 156362 324379 156365
rect 248952 156360 251239 156362
rect 248952 156304 251178 156360
rect 251234 156304 251239 156360
rect 248952 156302 251239 156304
rect 321908 156360 324379 156362
rect 321908 156304 324318 156360
rect 324374 156304 324379 156360
rect 321908 156302 324379 156304
rect 251173 156299 251239 156302
rect 324313 156299 324379 156302
rect 307661 156226 307727 156229
rect 307661 156224 310040 156226
rect 307661 156168 307666 156224
rect 307722 156168 310040 156224
rect 307661 156166 310040 156168
rect 307661 156163 307727 156166
rect 213913 155954 213979 155957
rect 252369 155954 252435 155957
rect 213913 155952 217242 155954
rect 213913 155896 213918 155952
rect 213974 155896 217242 155952
rect 213913 155894 217242 155896
rect 248952 155952 252435 155954
rect 248952 155896 252374 155952
rect 252430 155896 252435 155952
rect 248952 155894 252435 155896
rect 213913 155891 213979 155894
rect 217182 155788 217242 155894
rect 252369 155891 252435 155894
rect 306557 155682 306623 155685
rect 306557 155680 310040 155682
rect 306557 155624 306562 155680
rect 306618 155624 310040 155680
rect 306557 155622 310040 155624
rect 306557 155619 306623 155622
rect 214005 155410 214071 155413
rect 250069 155410 250135 155413
rect 214005 155408 217242 155410
rect 214005 155352 214010 155408
rect 214066 155352 217242 155408
rect 214005 155350 217242 155352
rect 248952 155408 250135 155410
rect 248952 155352 250074 155408
rect 250130 155352 250135 155408
rect 248952 155350 250135 155352
rect 214005 155347 214071 155350
rect 217182 155108 217242 155350
rect 250069 155347 250135 155350
rect 307661 155274 307727 155277
rect 307661 155272 310040 155274
rect 307661 155216 307666 155272
rect 307722 155216 310040 155272
rect 307661 155214 310040 155216
rect 307661 155211 307727 155214
rect 252461 155002 252527 155005
rect 248952 155000 252527 155002
rect 248952 154944 252466 155000
rect 252522 154944 252527 155000
rect 248952 154942 252527 154944
rect 252461 154939 252527 154942
rect 307293 154866 307359 154869
rect 321878 154866 321938 155516
rect 496905 155410 496971 155413
rect 494316 155408 496971 155410
rect 494316 155352 496910 155408
rect 496966 155352 496971 155408
rect 494316 155350 496971 155352
rect 496905 155347 496971 155350
rect 416773 155002 416839 155005
rect 416773 155000 420164 155002
rect 416773 154944 416778 155000
rect 416834 154944 420164 155000
rect 416773 154942 420164 154944
rect 416773 154939 416839 154942
rect 330334 154866 330340 154868
rect 307293 154864 310040 154866
rect 307293 154808 307298 154864
rect 307354 154808 310040 154864
rect 307293 154806 310040 154808
rect 321878 154806 330340 154866
rect 307293 154803 307359 154806
rect 330334 154804 330340 154806
rect 330404 154804 330410 154868
rect 323025 154730 323091 154733
rect 321908 154728 323091 154730
rect 321908 154672 323030 154728
rect 323086 154672 323091 154728
rect 321908 154670 323091 154672
rect 323025 154667 323091 154670
rect 252461 154458 252527 154461
rect 248952 154456 252527 154458
rect 213913 153914 213979 153917
rect 217182 153914 217242 154428
rect 248952 154400 252466 154456
rect 252522 154400 252527 154456
rect 248952 154398 252527 154400
rect 252461 154395 252527 154398
rect 307293 154458 307359 154461
rect 307293 154456 310040 154458
rect 307293 154400 307298 154456
rect 307354 154400 310040 154456
rect 307293 154398 310040 154400
rect 307293 154395 307359 154398
rect 496905 154322 496971 154325
rect 494316 154320 496971 154322
rect 494316 154264 496910 154320
rect 496966 154264 496971 154320
rect 494316 154262 496971 154264
rect 496905 154259 496971 154262
rect 307569 154050 307635 154053
rect 324313 154050 324379 154053
rect 307569 154048 310040 154050
rect 248860 153946 249442 154006
rect 307569 153992 307574 154048
rect 307630 153992 310040 154048
rect 307569 153990 310040 153992
rect 321908 154048 324379 154050
rect 321908 153992 324318 154048
rect 324374 153992 324379 154048
rect 321908 153990 324379 153992
rect 307569 153987 307635 153990
rect 324313 153987 324379 153990
rect 213913 153912 217242 153914
rect 213913 153856 213918 153912
rect 213974 153856 217242 153912
rect 213913 153854 217242 153856
rect 213913 153851 213979 153854
rect 213361 153234 213427 153237
rect 217182 153234 217242 153748
rect 249382 153506 249442 153946
rect 306649 153642 306715 153645
rect 306649 153640 310040 153642
rect 306649 153584 306654 153640
rect 306710 153584 310040 153640
rect 306649 153582 310040 153584
rect 306649 153579 306715 153582
rect 266302 153506 266308 153508
rect 248860 153402 249258 153462
rect 249382 153446 266308 153506
rect 266302 153444 266308 153446
rect 266372 153444 266378 153508
rect 249198 153370 249258 153402
rect 251449 153370 251515 153373
rect 249198 153368 251515 153370
rect 249198 153312 251454 153368
rect 251510 153312 251515 153368
rect 249198 153310 251515 153312
rect 251449 153307 251515 153310
rect 213361 153232 217242 153234
rect 213361 153176 213366 153232
rect 213422 153176 217242 153232
rect 213361 153174 217242 153176
rect 307661 153234 307727 153237
rect 324405 153234 324471 153237
rect 307661 153232 310040 153234
rect 307661 153176 307666 153232
rect 307722 153176 310040 153232
rect 307661 153174 310040 153176
rect 321908 153232 324471 153234
rect 321908 153176 324410 153232
rect 324466 153176 324471 153232
rect 321908 153174 324471 153176
rect 213361 153171 213427 153174
rect 307661 153171 307727 153174
rect 324405 153171 324471 153174
rect 416773 153234 416839 153237
rect 496997 153234 497063 153237
rect 416773 153232 420164 153234
rect 416773 153176 416778 153232
rect 416834 153176 420164 153232
rect 416773 153174 420164 153176
rect 494316 153232 497063 153234
rect 494316 153176 497002 153232
rect 497058 153176 497063 153232
rect 494316 153174 497063 153176
rect 416773 153171 416839 153174
rect 496997 153171 497063 153174
rect 252461 153098 252527 153101
rect 248952 153096 252527 153098
rect 214005 152690 214071 152693
rect 217182 152690 217242 153068
rect 248952 153040 252466 153096
rect 252522 153040 252527 153096
rect 248952 153038 252527 153040
rect 252461 153035 252527 153038
rect 252369 152690 252435 152693
rect 214005 152688 217242 152690
rect 214005 152632 214010 152688
rect 214066 152632 217242 152688
rect 214005 152630 217242 152632
rect 248952 152688 252435 152690
rect 248952 152632 252374 152688
rect 252430 152632 252435 152688
rect 248952 152630 252435 152632
rect 214005 152627 214071 152630
rect 252369 152627 252435 152630
rect 307477 152690 307543 152693
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 307477 152688 310040 152690
rect 307477 152632 307482 152688
rect 307538 152632 310040 152688
rect 307477 152630 310040 152632
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 307477 152627 307543 152630
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect 213913 152010 213979 152013
rect 217182 152010 217242 152524
rect 324313 152418 324379 152421
rect 321908 152416 324379 152418
rect 321908 152360 324318 152416
rect 324374 152360 324379 152416
rect 321908 152358 324379 152360
rect 324313 152355 324379 152358
rect 307569 152282 307635 152285
rect 307569 152280 310040 152282
rect 307569 152224 307574 152280
rect 307630 152224 310040 152280
rect 307569 152222 310040 152224
rect 307569 152219 307635 152222
rect 252277 152146 252343 152149
rect 496905 152146 496971 152149
rect 248952 152144 252343 152146
rect 248952 152088 252282 152144
rect 252338 152088 252343 152144
rect 248952 152086 252343 152088
rect 494316 152144 496971 152146
rect 494316 152088 496910 152144
rect 496966 152088 496971 152144
rect 494316 152086 496971 152088
rect 252277 152083 252343 152086
rect 496905 152083 496971 152086
rect 213913 152008 217242 152010
rect 213913 151952 213918 152008
rect 213974 151952 217242 152008
rect 213913 151950 217242 151952
rect 213913 151947 213979 151950
rect 215017 151874 215083 151877
rect 307661 151874 307727 151877
rect 215017 151872 217058 151874
rect 215017 151816 215022 151872
rect 215078 151830 217058 151872
rect 307661 151872 310040 151874
rect 217182 151830 217242 151844
rect 215078 151816 217242 151830
rect 215017 151814 217242 151816
rect 215017 151811 215083 151814
rect 216998 151770 217242 151814
rect 307661 151816 307666 151872
rect 307722 151816 310040 151872
rect 307661 151814 310040 151816
rect 307661 151811 307727 151814
rect 252645 151738 252711 151741
rect 324313 151738 324379 151741
rect 248952 151736 252711 151738
rect 248952 151680 252650 151736
rect 252706 151680 252711 151736
rect 248952 151678 252711 151680
rect 321908 151736 324379 151738
rect 321908 151680 324318 151736
rect 324374 151680 324379 151736
rect 321908 151678 324379 151680
rect 252645 151675 252711 151678
rect 324313 151675 324379 151678
rect 416773 151602 416839 151605
rect 416773 151600 420164 151602
rect 416773 151544 416778 151600
rect 416834 151544 420164 151600
rect 416773 151542 420164 151544
rect 416773 151539 416839 151542
rect 307569 151466 307635 151469
rect 307569 151464 310040 151466
rect 307569 151408 307574 151464
rect 307630 151408 310040 151464
rect 307569 151406 310040 151408
rect 307569 151403 307635 151406
rect 252461 151194 252527 151197
rect 248952 151192 252527 151194
rect 214005 150922 214071 150925
rect 217182 150922 217242 151164
rect 248952 151136 252466 151192
rect 252522 151136 252527 151192
rect 248952 151134 252527 151136
rect 252461 151131 252527 151134
rect 307661 151058 307727 151061
rect 307661 151056 310040 151058
rect 307661 151000 307666 151056
rect 307722 151000 310040 151056
rect 307661 150998 310040 151000
rect 307661 150995 307727 150998
rect 324405 150922 324471 150925
rect 496813 150922 496879 150925
rect 214005 150920 217242 150922
rect 214005 150864 214010 150920
rect 214066 150864 217242 150920
rect 214005 150862 217242 150864
rect 321908 150920 324471 150922
rect 321908 150864 324410 150920
rect 324466 150864 324471 150920
rect 321908 150862 324471 150864
rect 494316 150920 496879 150922
rect 494316 150864 496818 150920
rect 496874 150864 496879 150920
rect 494316 150862 496879 150864
rect 214005 150859 214071 150862
rect 324405 150859 324471 150862
rect 496813 150859 496879 150862
rect 251449 150786 251515 150789
rect 248952 150784 251515 150786
rect 248952 150728 251454 150784
rect 251510 150728 251515 150784
rect 248952 150726 251515 150728
rect 251449 150723 251515 150726
rect 213913 150650 213979 150653
rect 305821 150650 305887 150653
rect 213913 150648 217242 150650
rect 213913 150592 213918 150648
rect 213974 150592 217242 150648
rect 213913 150590 217242 150592
rect 213913 150587 213979 150590
rect 217182 150484 217242 150590
rect 305821 150648 310040 150650
rect 305821 150592 305826 150648
rect 305882 150592 310040 150648
rect 305821 150590 310040 150592
rect 305821 150587 305887 150590
rect 252461 150242 252527 150245
rect 248952 150240 252527 150242
rect 248952 150184 252466 150240
rect 252522 150184 252527 150240
rect 248952 150182 252527 150184
rect 252461 150179 252527 150182
rect 306741 150242 306807 150245
rect 306741 150240 310040 150242
rect 306741 150184 306746 150240
rect 306802 150184 310040 150240
rect 306741 150182 310040 150184
rect 306741 150179 306807 150182
rect 214005 150106 214071 150109
rect 324313 150106 324379 150109
rect 214005 150104 217242 150106
rect 214005 150048 214010 150104
rect 214066 150048 217242 150104
rect 214005 150046 217242 150048
rect 321908 150104 324379 150106
rect 321908 150048 324318 150104
rect 324374 150048 324379 150104
rect 321908 150046 324379 150048
rect 214005 150043 214071 150046
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect 217182 149804 217242 150046
rect 324313 150043 324379 150046
rect 249885 149834 249951 149837
rect 248952 149832 249951 149834
rect -960 149774 3483 149776
rect 248952 149776 249890 149832
rect 249946 149776 249951 149832
rect 248952 149774 249951 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 249885 149771 249951 149774
rect 307661 149834 307727 149837
rect 416773 149834 416839 149837
rect 496813 149834 496879 149837
rect 307661 149832 310040 149834
rect 307661 149776 307666 149832
rect 307722 149776 310040 149832
rect 307661 149774 310040 149776
rect 416773 149832 420164 149834
rect 416773 149776 416778 149832
rect 416834 149776 420164 149832
rect 416773 149774 420164 149776
rect 494316 149832 496879 149834
rect 494316 149776 496818 149832
rect 496874 149776 496879 149832
rect 494316 149774 496879 149776
rect 307661 149771 307727 149774
rect 416773 149771 416839 149774
rect 496813 149771 496879 149774
rect 251766 149636 251772 149700
rect 251836 149698 251842 149700
rect 304349 149698 304415 149701
rect 251836 149696 304415 149698
rect 251836 149640 304354 149696
rect 304410 149640 304415 149696
rect 251836 149638 304415 149640
rect 251836 149636 251842 149638
rect 304349 149635 304415 149638
rect 213913 149562 213979 149565
rect 213913 149560 217242 149562
rect 213913 149504 213918 149560
rect 213974 149504 217242 149560
rect 213913 149502 217242 149504
rect 213913 149499 213979 149502
rect 217182 149124 217242 149502
rect 324405 149426 324471 149429
rect 321908 149424 324471 149426
rect 321908 149368 324410 149424
rect 324466 149368 324471 149424
rect 321908 149366 324471 149368
rect 324405 149363 324471 149366
rect 251357 149290 251423 149293
rect 248952 149288 251423 149290
rect 248952 149232 251362 149288
rect 251418 149232 251423 149288
rect 248952 149230 251423 149232
rect 251357 149227 251423 149230
rect 307569 149290 307635 149293
rect 307569 149288 310040 149290
rect 307569 149232 307574 149288
rect 307630 149232 310040 149288
rect 307569 149230 310040 149232
rect 307569 149227 307635 149230
rect 494145 149018 494211 149021
rect 494102 149016 494211 149018
rect 494102 148960 494150 149016
rect 494206 148960 494211 149016
rect 494102 148955 494211 148960
rect 214741 148882 214807 148885
rect 252461 148882 252527 148885
rect 214741 148880 217242 148882
rect 214741 148824 214746 148880
rect 214802 148824 217242 148880
rect 214741 148822 217242 148824
rect 248952 148880 252527 148882
rect 248952 148824 252466 148880
rect 252522 148824 252527 148880
rect 248952 148822 252527 148824
rect 214741 148819 214807 148822
rect 217182 148444 217242 148822
rect 252461 148819 252527 148822
rect 307569 148882 307635 148885
rect 307569 148880 310040 148882
rect 307569 148824 307574 148880
rect 307630 148824 310040 148880
rect 307569 148822 310040 148824
rect 307569 148819 307635 148822
rect 494102 148716 494162 148955
rect 324313 148610 324379 148613
rect 321908 148608 324379 148610
rect 321908 148552 324318 148608
rect 324374 148552 324379 148608
rect 321908 148550 324379 148552
rect 324313 148547 324379 148550
rect 306925 148474 306991 148477
rect 306925 148472 310040 148474
rect 306925 148416 306930 148472
rect 306986 148416 310040 148472
rect 306925 148414 310040 148416
rect 306925 148411 306991 148414
rect 252369 148338 252435 148341
rect 248952 148336 252435 148338
rect 248952 148280 252374 148336
rect 252430 148280 252435 148336
rect 248952 148278 252435 148280
rect 252369 148275 252435 148278
rect 254526 148276 254532 148340
rect 254596 148338 254602 148340
rect 273345 148338 273411 148341
rect 254596 148336 273411 148338
rect 254596 148280 273350 148336
rect 273406 148280 273411 148336
rect 254596 148278 273411 148280
rect 254596 148276 254602 148278
rect 273345 148275 273411 148278
rect 416773 148202 416839 148205
rect 416773 148200 420164 148202
rect 416773 148144 416778 148200
rect 416834 148144 420164 148200
rect 416773 148142 420164 148144
rect 416773 148139 416839 148142
rect 214557 148066 214623 148069
rect 307661 148066 307727 148069
rect 214557 148064 217242 148066
rect 214557 148008 214562 148064
rect 214618 148008 217242 148064
rect 214557 148006 217242 148008
rect 214557 148003 214623 148006
rect 217182 147900 217242 148006
rect 307661 148064 310040 148066
rect 307661 148008 307666 148064
rect 307722 148008 310040 148064
rect 307661 148006 310040 148008
rect 307661 148003 307727 148006
rect 255262 147930 255268 147932
rect 248952 147870 255268 147930
rect 255262 147868 255268 147870
rect 255332 147868 255338 147932
rect 324405 147794 324471 147797
rect 321908 147792 324471 147794
rect 321908 147736 324410 147792
rect 324466 147736 324471 147792
rect 321908 147734 324471 147736
rect 324405 147731 324471 147734
rect 331254 147732 331260 147796
rect 331324 147794 331330 147796
rect 331857 147794 331923 147797
rect 332501 147794 332567 147797
rect 331324 147792 332567 147794
rect 331324 147736 331862 147792
rect 331918 147736 332506 147792
rect 332562 147736 332567 147792
rect 331324 147734 332567 147736
rect 331324 147732 331330 147734
rect 331857 147731 331923 147734
rect 332501 147731 332567 147734
rect 307385 147658 307451 147661
rect 496813 147658 496879 147661
rect 307385 147656 310040 147658
rect 307385 147600 307390 147656
rect 307446 147600 310040 147656
rect 307385 147598 310040 147600
rect 494316 147656 496879 147658
rect 494316 147600 496818 147656
rect 496874 147600 496879 147656
rect 494316 147598 496879 147600
rect 307385 147595 307451 147598
rect 496813 147595 496879 147598
rect 252461 147522 252527 147525
rect 248952 147520 252527 147522
rect 248952 147464 252466 147520
rect 252522 147464 252527 147520
rect 248952 147462 252527 147464
rect 252461 147459 252527 147462
rect 307569 147250 307635 147253
rect 307569 147248 310040 147250
rect 214005 146706 214071 146709
rect 217182 146706 217242 147220
rect 307569 147192 307574 147248
rect 307630 147192 310040 147248
rect 307569 147190 310040 147192
rect 307569 147187 307635 147190
rect 324313 147114 324379 147117
rect 321908 147112 324379 147114
rect 321908 147056 324318 147112
rect 324374 147056 324379 147112
rect 321908 147054 324379 147056
rect 324313 147051 324379 147054
rect 252093 146978 252159 146981
rect 248952 146976 252159 146978
rect 248952 146920 252098 146976
rect 252154 146920 252159 146976
rect 248952 146918 252159 146920
rect 252093 146915 252159 146918
rect 306741 146842 306807 146845
rect 306741 146840 310040 146842
rect 306741 146784 306746 146840
rect 306802 146784 310040 146840
rect 306741 146782 310040 146784
rect 306741 146779 306807 146782
rect 214005 146704 217242 146706
rect 214005 146648 214010 146704
rect 214066 146648 217242 146704
rect 214005 146646 217242 146648
rect 214005 146643 214071 146646
rect 251357 146570 251423 146573
rect 248952 146568 251423 146570
rect 213913 146434 213979 146437
rect 213913 146432 216874 146434
rect 213913 146376 213918 146432
rect 213974 146376 216874 146432
rect 213913 146374 216874 146376
rect 213913 146371 213979 146374
rect 216814 146298 216874 146374
rect 217366 146298 217426 146540
rect 248952 146512 251362 146568
rect 251418 146512 251423 146568
rect 248952 146510 251423 146512
rect 251357 146507 251423 146510
rect 416773 146570 416839 146573
rect 416773 146568 420164 146570
rect 416773 146512 416778 146568
rect 416834 146512 420164 146568
rect 416773 146510 420164 146512
rect 416773 146507 416839 146510
rect 307661 146434 307727 146437
rect 307661 146432 310040 146434
rect 307661 146376 307666 146432
rect 307722 146376 310040 146432
rect 307661 146374 310040 146376
rect 307661 146371 307727 146374
rect 494102 146301 494162 146404
rect 324313 146298 324379 146301
rect 216814 146238 217426 146298
rect 321908 146296 324379 146298
rect 321908 146240 324318 146296
rect 324374 146240 324379 146296
rect 321908 146238 324379 146240
rect 494102 146296 494211 146301
rect 494102 146240 494150 146296
rect 494206 146240 494211 146296
rect 494102 146238 494211 146240
rect 324313 146235 324379 146238
rect 494145 146235 494211 146238
rect 254526 146026 254532 146028
rect 248952 145966 254532 146026
rect 254526 145964 254532 145966
rect 254596 145964 254602 146028
rect 307661 145890 307727 145893
rect 307661 145888 310040 145890
rect 213913 145346 213979 145349
rect 217182 145346 217242 145860
rect 307661 145832 307666 145888
rect 307722 145832 310040 145888
rect 307661 145830 310040 145832
rect 307661 145827 307727 145830
rect 252461 145618 252527 145621
rect 248952 145616 252527 145618
rect 248952 145560 252466 145616
rect 252522 145560 252527 145616
rect 248952 145558 252527 145560
rect 252461 145555 252527 145558
rect 257429 145618 257495 145621
rect 306966 145618 306972 145620
rect 257429 145616 306972 145618
rect 257429 145560 257434 145616
rect 257490 145560 306972 145616
rect 257429 145558 306972 145560
rect 257429 145555 257495 145558
rect 306966 145556 306972 145558
rect 307036 145556 307042 145620
rect 307569 145482 307635 145485
rect 324589 145482 324655 145485
rect 307569 145480 310040 145482
rect 307569 145424 307574 145480
rect 307630 145424 310040 145480
rect 307569 145422 310040 145424
rect 321908 145480 324655 145482
rect 321908 145424 324594 145480
rect 324650 145424 324655 145480
rect 321908 145422 324655 145424
rect 307569 145419 307635 145422
rect 324589 145419 324655 145422
rect 496813 145346 496879 145349
rect 213913 145344 217242 145346
rect 213913 145288 213918 145344
rect 213974 145288 217242 145344
rect 213913 145286 217242 145288
rect 494316 145344 496879 145346
rect 494316 145288 496818 145344
rect 496874 145288 496879 145344
rect 494316 145286 496879 145288
rect 213913 145283 213979 145286
rect 496813 145283 496879 145286
rect 214741 144938 214807 144941
rect 217182 144938 217242 145180
rect 252369 145074 252435 145077
rect 248952 145072 252435 145074
rect 248952 145016 252374 145072
rect 252430 145016 252435 145072
rect 248952 145014 252435 145016
rect 252369 145011 252435 145014
rect 307702 145012 307708 145076
rect 307772 145074 307778 145076
rect 307772 145014 310040 145074
rect 307772 145012 307778 145014
rect 214741 144936 217242 144938
rect 214741 144880 214746 144936
rect 214802 144880 217242 144936
rect 214741 144878 217242 144880
rect 214741 144875 214807 144878
rect 324313 144802 324379 144805
rect 321908 144800 324379 144802
rect 321908 144744 324318 144800
rect 324374 144744 324379 144800
rect 321908 144742 324379 144744
rect 324313 144739 324379 144742
rect 416773 144802 416839 144805
rect 416773 144800 420164 144802
rect 416773 144744 416778 144800
rect 416834 144744 420164 144800
rect 416773 144742 420164 144744
rect 416773 144739 416839 144742
rect 307661 144666 307727 144669
rect 307661 144664 310040 144666
rect 248860 144562 249442 144622
rect 307661 144608 307666 144664
rect 307722 144608 310040 144664
rect 307661 144606 310040 144608
rect 307661 144603 307727 144606
rect 214005 143986 214071 143989
rect 217182 143986 217242 144500
rect 249382 144394 249442 144562
rect 259494 144394 259500 144396
rect 249382 144334 259500 144394
rect 259494 144332 259500 144334
rect 259564 144332 259570 144396
rect 306925 144258 306991 144261
rect 496813 144258 496879 144261
rect 306925 144256 310040 144258
rect 306925 144200 306930 144256
rect 306986 144200 310040 144256
rect 306925 144198 310040 144200
rect 494316 144256 496879 144258
rect 494316 144200 496818 144256
rect 496874 144200 496879 144256
rect 494316 144198 496879 144200
rect 306925 144195 306991 144198
rect 496813 144195 496879 144198
rect 252461 144122 252527 144125
rect 248952 144120 252527 144122
rect 248952 144064 252466 144120
rect 252522 144064 252527 144120
rect 248952 144062 252527 144064
rect 252461 144059 252527 144062
rect 214005 143984 217242 143986
rect 214005 143928 214010 143984
rect 214066 143928 217242 143984
rect 214005 143926 217242 143928
rect 303153 143986 303219 143989
rect 307702 143986 307708 143988
rect 303153 143984 307708 143986
rect 303153 143928 303158 143984
rect 303214 143928 307708 143984
rect 303153 143926 307708 143928
rect 214005 143923 214071 143926
rect 303153 143923 303219 143926
rect 307702 143924 307708 143926
rect 307772 143924 307778 143988
rect 327206 143986 327212 143988
rect 321908 143926 327212 143986
rect 327206 143924 327212 143926
rect 327276 143924 327282 143988
rect 307569 143850 307635 143853
rect 307569 143848 310040 143850
rect 213913 143578 213979 143581
rect 217366 143578 217426 143820
rect 307569 143792 307574 143848
rect 307630 143792 310040 143848
rect 307569 143790 310040 143792
rect 307569 143787 307635 143790
rect 252369 143714 252435 143717
rect 248952 143712 252435 143714
rect 248952 143656 252374 143712
rect 252430 143656 252435 143712
rect 248952 143654 252435 143656
rect 252369 143651 252435 143654
rect 213913 143576 217426 143578
rect 213913 143520 213918 143576
rect 213974 143520 217426 143576
rect 213913 143518 217426 143520
rect 213913 143515 213979 143518
rect 307661 143442 307727 143445
rect 307661 143440 310040 143442
rect 307661 143384 307666 143440
rect 307722 143384 310040 143440
rect 307661 143382 310040 143384
rect 307661 143379 307727 143382
rect 214005 142762 214071 142765
rect 217182 142762 217242 143276
rect 252461 143170 252527 143173
rect 324405 143170 324471 143173
rect 248952 143168 252527 143170
rect 248952 143112 252466 143168
rect 252522 143112 252527 143168
rect 248952 143110 252527 143112
rect 321908 143168 324471 143170
rect 321908 143112 324410 143168
rect 324466 143112 324471 143168
rect 321908 143110 324471 143112
rect 252461 143107 252527 143110
rect 324405 143107 324471 143110
rect 416865 143170 416931 143173
rect 496813 143170 496879 143173
rect 416865 143168 420164 143170
rect 416865 143112 416870 143168
rect 416926 143112 420164 143168
rect 416865 143110 420164 143112
rect 494316 143168 496879 143170
rect 494316 143112 496818 143168
rect 496874 143112 496879 143168
rect 494316 143110 496879 143112
rect 416865 143107 416931 143110
rect 496813 143107 496879 143110
rect 306557 143034 306623 143037
rect 306557 143032 310040 143034
rect 306557 142976 306562 143032
rect 306618 142976 310040 143032
rect 306557 142974 310040 142976
rect 306557 142971 306623 142974
rect 252369 142762 252435 142765
rect 214005 142760 217242 142762
rect 214005 142704 214010 142760
rect 214066 142704 217242 142760
rect 214005 142702 217242 142704
rect 248952 142760 252435 142762
rect 248952 142704 252374 142760
rect 252430 142704 252435 142760
rect 248952 142702 252435 142704
rect 214005 142699 214071 142702
rect 252369 142699 252435 142702
rect 213913 142354 213979 142357
rect 217182 142354 217242 142596
rect 307109 142490 307175 142493
rect 324313 142490 324379 142493
rect 307109 142488 310040 142490
rect 307109 142432 307114 142488
rect 307170 142432 310040 142488
rect 307109 142430 310040 142432
rect 321908 142488 324379 142490
rect 321908 142432 324318 142488
rect 324374 142432 324379 142488
rect 321908 142430 324379 142432
rect 307109 142427 307175 142430
rect 324313 142427 324379 142430
rect 213913 142352 217242 142354
rect 213913 142296 213918 142352
rect 213974 142296 217242 142352
rect 213913 142294 217242 142296
rect 213913 142291 213979 142294
rect 263726 142218 263732 142220
rect 248952 142158 263732 142218
rect 263726 142156 263732 142158
rect 263796 142156 263802 142220
rect 306557 142082 306623 142085
rect 306557 142080 310040 142082
rect 306557 142024 306562 142080
rect 306618 142024 310040 142080
rect 306557 142022 310040 142024
rect 306557 142019 306623 142022
rect 496813 141946 496879 141949
rect 494316 141944 496879 141946
rect 214005 141402 214071 141405
rect 217182 141402 217242 141916
rect 494316 141888 496818 141944
rect 496874 141888 496879 141944
rect 494316 141886 496879 141888
rect 496813 141883 496879 141886
rect 253473 141810 253539 141813
rect 248952 141808 253539 141810
rect 248952 141752 253478 141808
rect 253534 141752 253539 141808
rect 248952 141750 253539 141752
rect 253473 141747 253539 141750
rect 307569 141674 307635 141677
rect 324313 141674 324379 141677
rect 307569 141672 310040 141674
rect 307569 141616 307574 141672
rect 307630 141616 310040 141672
rect 307569 141614 310040 141616
rect 321908 141672 324379 141674
rect 321908 141616 324318 141672
rect 324374 141616 324379 141672
rect 321908 141614 324379 141616
rect 307569 141611 307635 141614
rect 324313 141611 324379 141614
rect 214005 141400 217242 141402
rect 214005 141344 214010 141400
rect 214066 141344 217242 141400
rect 416773 141402 416839 141405
rect 416773 141400 420164 141402
rect 214005 141342 217242 141344
rect 214005 141339 214071 141342
rect 248860 141298 249442 141358
rect 416773 141344 416778 141400
rect 416834 141344 420164 141400
rect 416773 141342 420164 141344
rect 416773 141339 416839 141342
rect 213913 140858 213979 140861
rect 217182 140858 217242 141236
rect 249382 141130 249442 141298
rect 307477 141266 307543 141269
rect 494237 141266 494303 141269
rect 307477 141264 310040 141266
rect 307477 141208 307482 141264
rect 307538 141208 310040 141264
rect 307477 141206 310040 141208
rect 494237 141264 494346 141266
rect 494237 141208 494242 141264
rect 494298 141208 494346 141264
rect 307477 141203 307543 141206
rect 494237 141203 494346 141208
rect 259678 141130 259684 141132
rect 249382 141070 259684 141130
rect 259678 141068 259684 141070
rect 259748 141068 259754 141132
rect 253473 140994 253539 140997
rect 258390 140994 258396 140996
rect 253473 140992 258396 140994
rect 253473 140936 253478 140992
rect 253534 140936 258396 140992
rect 253473 140934 258396 140936
rect 253473 140931 253539 140934
rect 258390 140932 258396 140934
rect 258460 140932 258466 140996
rect 253197 140858 253263 140861
rect 213913 140856 217242 140858
rect 213913 140800 213918 140856
rect 213974 140800 217242 140856
rect 213913 140798 217242 140800
rect 248952 140856 253263 140858
rect 248952 140800 253202 140856
rect 253258 140800 253263 140856
rect 248952 140798 253263 140800
rect 213913 140795 213979 140798
rect 253197 140795 253263 140798
rect 307661 140858 307727 140861
rect 324405 140858 324471 140861
rect 307661 140856 310040 140858
rect 307661 140800 307666 140856
rect 307722 140800 310040 140856
rect 307661 140798 310040 140800
rect 321908 140856 324471 140858
rect 321908 140800 324410 140856
rect 324466 140800 324471 140856
rect 494286 140858 494346 141203
rect 495341 140858 495407 140861
rect 494286 140856 495407 140858
rect 494286 140828 495346 140856
rect 321908 140798 324471 140800
rect 494316 140800 495346 140828
rect 495402 140800 495407 140856
rect 494316 140798 495407 140800
rect 307661 140795 307727 140798
rect 324405 140795 324471 140798
rect 495341 140795 495407 140798
rect 213913 140042 213979 140045
rect 217182 140042 217242 140556
rect 255446 140450 255452 140452
rect 248952 140390 255452 140450
rect 255446 140388 255452 140390
rect 255516 140388 255522 140452
rect 307569 140450 307635 140453
rect 307569 140448 310040 140450
rect 307569 140392 307574 140448
rect 307630 140392 310040 140448
rect 307569 140390 310040 140392
rect 307569 140387 307635 140390
rect 326654 140178 326660 140180
rect 321908 140118 326660 140178
rect 326654 140116 326660 140118
rect 326724 140116 326730 140180
rect 213913 140040 217242 140042
rect 213913 139984 213918 140040
rect 213974 139984 217242 140040
rect 213913 139982 217242 139984
rect 307661 140042 307727 140045
rect 307661 140040 310040 140042
rect 307661 139984 307666 140040
rect 307722 139984 310040 140040
rect 307661 139982 310040 139984
rect 213913 139979 213979 139982
rect 307661 139979 307727 139982
rect 252461 139906 252527 139909
rect 248952 139904 252527 139906
rect 214649 139634 214715 139637
rect 217182 139634 217242 139876
rect 248952 139848 252466 139904
rect 252522 139848 252527 139904
rect 248952 139846 252527 139848
rect 252461 139843 252527 139846
rect 416773 139770 416839 139773
rect 496813 139770 496879 139773
rect 416773 139768 420164 139770
rect 416773 139712 416778 139768
rect 416834 139712 420164 139768
rect 416773 139710 420164 139712
rect 494316 139768 496879 139770
rect 494316 139712 496818 139768
rect 496874 139712 496879 139768
rect 494316 139710 496879 139712
rect 416773 139707 416839 139710
rect 496813 139707 496879 139710
rect 214649 139632 217242 139634
rect 214649 139576 214654 139632
rect 214710 139576 217242 139632
rect 214649 139574 217242 139576
rect 307293 139634 307359 139637
rect 307293 139632 310040 139634
rect 307293 139576 307298 139632
rect 307354 139576 310040 139632
rect 307293 139574 310040 139576
rect 214649 139571 214715 139574
rect 307293 139571 307359 139574
rect 249793 139498 249859 139501
rect 248952 139496 249859 139498
rect 248952 139440 249798 139496
rect 249854 139440 249859 139496
rect 248952 139438 249859 139440
rect 249793 139435 249859 139438
rect 327022 139362 327028 139364
rect 321908 139302 327028 139362
rect 327022 139300 327028 139302
rect 327092 139300 327098 139364
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect 213913 138818 213979 138821
rect 217182 138818 217242 139196
rect 306557 139090 306623 139093
rect 306557 139088 310040 139090
rect 306557 139032 306562 139088
rect 306618 139032 310040 139088
rect 306557 139030 310040 139032
rect 306557 139027 306623 139030
rect 248860 138850 249442 138910
rect 213913 138816 217242 138818
rect 213913 138760 213918 138816
rect 213974 138760 217242 138816
rect 213913 138758 217242 138760
rect 213913 138755 213979 138758
rect 249382 138682 249442 138850
rect 262254 138682 262260 138684
rect 214649 138138 214715 138141
rect 217182 138138 217242 138652
rect 249382 138622 262260 138682
rect 262254 138620 262260 138622
rect 262324 138620 262330 138684
rect 307293 138682 307359 138685
rect 496813 138682 496879 138685
rect 307293 138680 310040 138682
rect 307293 138624 307298 138680
rect 307354 138624 310040 138680
rect 307293 138622 310040 138624
rect 494316 138680 496879 138682
rect 494316 138624 496818 138680
rect 496874 138624 496879 138680
rect 494316 138622 496879 138624
rect 307293 138619 307359 138622
rect 496813 138619 496879 138622
rect 252461 138546 252527 138549
rect 324313 138546 324379 138549
rect 248952 138544 252527 138546
rect 248952 138488 252466 138544
rect 252522 138488 252527 138544
rect 248952 138486 252527 138488
rect 321908 138544 324379 138546
rect 321908 138488 324318 138544
rect 324374 138488 324379 138544
rect 321908 138486 324379 138488
rect 252461 138483 252527 138486
rect 324313 138483 324379 138486
rect 307661 138274 307727 138277
rect 307661 138272 310040 138274
rect 307661 138216 307666 138272
rect 307722 138216 310040 138272
rect 307661 138214 310040 138216
rect 307661 138211 307727 138214
rect 214649 138136 217242 138138
rect 214649 138080 214654 138136
rect 214710 138080 217242 138136
rect 214649 138078 217242 138080
rect 214649 138075 214715 138078
rect 416773 138002 416839 138005
rect 416773 138000 420164 138002
rect 214005 137458 214071 137461
rect 217182 137458 217242 137972
rect 248860 137898 249442 137958
rect 416773 137944 416778 138000
rect 416834 137944 420164 138000
rect 416773 137942 420164 137944
rect 416773 137939 416839 137942
rect 249382 137730 249442 137898
rect 307661 137866 307727 137869
rect 324313 137866 324379 137869
rect 307661 137864 310040 137866
rect 307661 137808 307666 137864
rect 307722 137808 310040 137864
rect 307661 137806 310040 137808
rect 321908 137864 324379 137866
rect 321908 137808 324318 137864
rect 324374 137808 324379 137864
rect 321908 137806 324379 137808
rect 307661 137803 307727 137806
rect 324313 137803 324379 137806
rect 249382 137670 253490 137730
rect 248860 137490 249442 137550
rect 214005 137456 217242 137458
rect 214005 137400 214010 137456
rect 214066 137400 217242 137456
rect 214005 137398 217242 137400
rect 214005 137395 214071 137398
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 213913 136778 213979 136781
rect 217182 136778 217242 137292
rect 248860 136946 249258 137006
rect 213913 136776 217242 136778
rect 213913 136720 213918 136776
rect 213974 136720 217242 136776
rect 213913 136718 217242 136720
rect 249198 136778 249258 136946
rect 249382 136914 249442 137490
rect 253430 137050 253490 137670
rect 496813 137458 496879 137461
rect 494316 137456 496879 137458
rect 309504 137354 310132 137414
rect 494316 137400 496818 137456
rect 496874 137400 496879 137456
rect 494316 137398 496879 137400
rect 496813 137395 496879 137398
rect 253606 137124 253612 137188
rect 253676 137186 253682 137188
rect 309504 137186 309564 137354
rect 253676 137126 309564 137186
rect 253676 137124 253682 137126
rect 263542 137050 263548 137052
rect 253430 136990 263548 137050
rect 263542 136988 263548 136990
rect 263612 136988 263618 137052
rect 307201 137050 307267 137053
rect 324405 137050 324471 137053
rect 307201 137048 310040 137050
rect 307201 136992 307206 137048
rect 307262 136992 310040 137048
rect 307201 136990 310040 136992
rect 321908 137048 324471 137050
rect 321908 136992 324410 137048
rect 324466 136992 324471 137048
rect 321908 136990 324471 136992
rect 307201 136987 307267 136990
rect 324405 136987 324471 136990
rect 269062 136914 269068 136916
rect 249382 136854 269068 136914
rect 269062 136852 269068 136854
rect 269132 136852 269138 136916
rect 252461 136778 252527 136781
rect 249198 136776 252527 136778
rect 249198 136720 252466 136776
rect 252522 136720 252527 136776
rect 249198 136718 252527 136720
rect 213913 136715 213979 136718
rect 252461 136715 252527 136718
rect 252461 136642 252527 136645
rect 248952 136640 252527 136642
rect 213913 136098 213979 136101
rect 217182 136098 217242 136612
rect 248952 136584 252466 136640
rect 252522 136584 252527 136640
rect 248952 136582 252527 136584
rect 252461 136579 252527 136582
rect 306557 136642 306623 136645
rect 306557 136640 310040 136642
rect 306557 136584 306562 136640
rect 306618 136584 310040 136640
rect 306557 136582 310040 136584
rect 306557 136579 306623 136582
rect 324313 136370 324379 136373
rect 321908 136368 324379 136370
rect 321908 136312 324318 136368
rect 324374 136312 324379 136368
rect 321908 136310 324379 136312
rect 324313 136307 324379 136310
rect 416773 136370 416839 136373
rect 496813 136370 496879 136373
rect 416773 136368 420164 136370
rect 416773 136312 416778 136368
rect 416834 136312 420164 136368
rect 416773 136310 420164 136312
rect 494316 136368 496879 136370
rect 494316 136312 496818 136368
rect 496874 136312 496879 136368
rect 494316 136310 496879 136312
rect 416773 136307 416839 136310
rect 496813 136307 496879 136310
rect 252277 136234 252343 136237
rect 248952 136232 252343 136234
rect 248952 136176 252282 136232
rect 252338 136176 252343 136232
rect 248952 136174 252343 136176
rect 252277 136171 252343 136174
rect 307569 136234 307635 136237
rect 307569 136232 310040 136234
rect 307569 136176 307574 136232
rect 307630 136176 310040 136232
rect 307569 136174 310040 136176
rect 307569 136171 307635 136174
rect 213913 136096 217242 136098
rect 213913 136040 213918 136096
rect 213974 136040 217242 136096
rect 213913 136038 217242 136040
rect 213913 136035 213979 136038
rect 169150 135492 169156 135556
rect 169220 135554 169226 135556
rect 217182 135554 217242 135932
rect 252369 135690 252435 135693
rect 248952 135688 252435 135690
rect 248952 135632 252374 135688
rect 252430 135632 252435 135688
rect 248952 135630 252435 135632
rect 252369 135627 252435 135630
rect 307661 135690 307727 135693
rect 307661 135688 310040 135690
rect 307661 135632 307666 135688
rect 307722 135632 310040 135688
rect 307661 135630 310040 135632
rect 307661 135627 307727 135630
rect 324405 135554 324471 135557
rect 169220 135494 217242 135554
rect 321908 135552 324471 135554
rect 321908 135496 324410 135552
rect 324466 135496 324471 135552
rect 321908 135494 324471 135496
rect 169220 135492 169226 135494
rect 324405 135491 324471 135494
rect 170254 135356 170260 135420
rect 170324 135418 170330 135420
rect 170324 135358 217242 135418
rect 170324 135356 170330 135358
rect 217182 135252 217242 135358
rect 252185 135282 252251 135285
rect 248952 135280 252251 135282
rect 248952 135224 252190 135280
rect 252246 135224 252251 135280
rect 248952 135222 252251 135224
rect 252185 135219 252251 135222
rect 307293 135282 307359 135285
rect 496905 135282 496971 135285
rect 307293 135280 310040 135282
rect 307293 135224 307298 135280
rect 307354 135224 310040 135280
rect 307293 135222 310040 135224
rect 494316 135280 496971 135282
rect 494316 135224 496910 135280
rect 496966 135224 496971 135280
rect 494316 135222 496971 135224
rect 307293 135219 307359 135222
rect 496905 135219 496971 135222
rect 306557 134874 306623 134877
rect 306557 134872 310040 134874
rect 306557 134816 306562 134872
rect 306618 134816 310040 134872
rect 306557 134814 310040 134816
rect 306557 134811 306623 134814
rect 252461 134738 252527 134741
rect 248952 134736 252527 134738
rect 248952 134680 252466 134736
rect 252522 134680 252527 134736
rect 248952 134678 252527 134680
rect 252461 134675 252527 134678
rect 214005 134330 214071 134333
rect 217182 134330 217242 134572
rect 309504 134362 310132 134422
rect 252369 134330 252435 134333
rect 214005 134328 217242 134330
rect 214005 134272 214010 134328
rect 214066 134272 217242 134328
rect 214005 134270 217242 134272
rect 248952 134328 252435 134330
rect 248952 134272 252374 134328
rect 252430 134272 252435 134328
rect 248952 134270 252435 134272
rect 214005 134267 214071 134270
rect 252369 134267 252435 134270
rect 250294 134132 250300 134196
rect 250364 134194 250370 134196
rect 309504 134194 309564 134362
rect 250364 134134 309564 134194
rect 321878 134194 321938 134708
rect 417325 134602 417391 134605
rect 419257 134602 419323 134605
rect 417325 134600 420164 134602
rect 417325 134544 417330 134600
rect 417386 134544 419262 134600
rect 419318 134544 420164 134600
rect 417325 134542 420164 134544
rect 417325 134539 417391 134542
rect 419257 134539 419323 134542
rect 323485 134194 323551 134197
rect 321878 134192 323551 134194
rect 321878 134136 323490 134192
rect 323546 134136 323551 134192
rect 321878 134134 323551 134136
rect 250364 134132 250370 134134
rect 323485 134131 323551 134134
rect 213913 134058 213979 134061
rect 307017 134058 307083 134061
rect 328494 134058 328500 134060
rect 213913 134056 217242 134058
rect 213913 134000 213918 134056
rect 213974 134000 217242 134056
rect 213913 133998 217242 134000
rect 213913 133995 213979 133998
rect 217182 133892 217242 133998
rect 307017 134056 310040 134058
rect 307017 134000 307022 134056
rect 307078 134000 310040 134056
rect 307017 133998 310040 134000
rect 321908 133998 328500 134058
rect 307017 133995 307083 133998
rect 328494 133996 328500 133998
rect 328564 133996 328570 134060
rect 323485 133922 323551 133925
rect 332542 133922 332548 133924
rect 323485 133920 332548 133922
rect 323485 133864 323490 133920
rect 323546 133864 332548 133920
rect 323485 133862 332548 133864
rect 323485 133859 323551 133862
rect 332542 133860 332548 133862
rect 332612 133860 332618 133924
rect 494286 133922 494346 134164
rect 502374 133922 502380 133924
rect 494286 133862 502380 133922
rect 502374 133860 502380 133862
rect 502444 133860 502450 133924
rect 252461 133786 252527 133789
rect 321737 133786 321803 133789
rect 248952 133784 252527 133786
rect 248952 133728 252466 133784
rect 252522 133728 252527 133784
rect 248952 133726 252527 133728
rect 252461 133723 252527 133726
rect 321694 133784 321803 133786
rect 321694 133728 321742 133784
rect 321798 133728 321803 133784
rect 321694 133723 321803 133728
rect 306557 133650 306623 133653
rect 306557 133648 310040 133650
rect 306557 133592 306562 133648
rect 306618 133592 310040 133648
rect 306557 133590 310040 133592
rect 306557 133587 306623 133590
rect 252277 133378 252343 133381
rect 248952 133376 252343 133378
rect 213913 132970 213979 132973
rect 217182 132970 217242 133348
rect 248952 133320 252282 133376
rect 252338 133320 252343 133376
rect 248952 133318 252343 133320
rect 252277 133315 252343 133318
rect 306925 133242 306991 133245
rect 306925 133240 310040 133242
rect 306925 133184 306930 133240
rect 306986 133184 310040 133240
rect 321694 133212 321754 133723
rect 306925 133182 310040 133184
rect 306925 133179 306991 133182
rect 213913 132968 217242 132970
rect 213913 132912 213918 132968
rect 213974 132912 217242 132968
rect 213913 132910 217242 132912
rect 419441 132970 419507 132973
rect 496813 132970 496879 132973
rect 419441 132968 420164 132970
rect 419441 132912 419446 132968
rect 419502 132912 420164 132968
rect 419441 132910 420164 132912
rect 494316 132968 496879 132970
rect 494316 132912 496818 132968
rect 496874 132912 496879 132968
rect 494316 132910 496879 132912
rect 213913 132907 213979 132910
rect 419441 132907 419507 132910
rect 496813 132907 496879 132910
rect 213913 132834 213979 132837
rect 252369 132834 252435 132837
rect 213913 132832 217242 132834
rect 213913 132776 213918 132832
rect 213974 132776 217242 132832
rect 213913 132774 217242 132776
rect 248952 132832 252435 132834
rect 248952 132776 252374 132832
rect 252430 132776 252435 132832
rect 248952 132774 252435 132776
rect 213913 132771 213979 132774
rect 217182 132668 217242 132774
rect 252369 132771 252435 132774
rect 307293 132698 307359 132701
rect 307293 132696 310040 132698
rect 307293 132640 307298 132696
rect 307354 132640 310040 132696
rect 307293 132638 310040 132640
rect 307293 132635 307359 132638
rect 252461 132426 252527 132429
rect 325877 132426 325943 132429
rect 248952 132424 252527 132426
rect 248952 132368 252466 132424
rect 252522 132368 252527 132424
rect 248952 132366 252527 132368
rect 321908 132424 325943 132426
rect 321908 132368 325882 132424
rect 325938 132368 325943 132424
rect 321908 132366 325943 132368
rect 252461 132363 252527 132366
rect 325877 132363 325943 132366
rect 307477 132290 307543 132293
rect 307477 132288 310040 132290
rect 307477 132232 307482 132288
rect 307538 132232 310040 132288
rect 307477 132230 310040 132232
rect 307477 132227 307543 132230
rect 321502 132092 321508 132156
rect 321572 132092 321578 132156
rect 494329 132154 494395 132157
rect 494286 132152 494395 132154
rect 494286 132096 494334 132152
rect 494390 132096 494395 132152
rect 213913 131474 213979 131477
rect 217182 131474 217242 131988
rect 252277 131882 252343 131885
rect 248952 131880 252343 131882
rect 248952 131824 252282 131880
rect 252338 131824 252343 131880
rect 248952 131822 252343 131824
rect 252277 131819 252343 131822
rect 307569 131882 307635 131885
rect 307569 131880 310040 131882
rect 307569 131824 307574 131880
rect 307630 131824 310040 131880
rect 307569 131822 310040 131824
rect 307569 131819 307635 131822
rect 321510 131716 321570 132092
rect 494286 132091 494395 132096
rect 494286 131852 494346 132091
rect 252369 131474 252435 131477
rect 213913 131472 217242 131474
rect 213913 131416 213918 131472
rect 213974 131416 217242 131472
rect 213913 131414 217242 131416
rect 248952 131472 252435 131474
rect 248952 131416 252374 131472
rect 252430 131416 252435 131472
rect 248952 131414 252435 131416
rect 213913 131411 213979 131414
rect 252369 131411 252435 131414
rect 307661 131474 307727 131477
rect 307661 131472 310040 131474
rect 307661 131416 307666 131472
rect 307722 131416 310040 131472
rect 307661 131414 310040 131416
rect 307661 131411 307727 131414
rect 417509 131338 417575 131341
rect 419717 131338 419783 131341
rect 417509 131336 420164 131338
rect 170438 131140 170444 131204
rect 170508 131202 170514 131204
rect 170508 131142 216874 131202
rect 170508 131140 170514 131142
rect 216814 131066 216874 131142
rect 217366 131066 217426 131308
rect 417509 131280 417514 131336
rect 417570 131280 419722 131336
rect 419778 131280 420164 131336
rect 417509 131278 420164 131280
rect 417509 131275 417575 131278
rect 419717 131275 419783 131278
rect 216814 131006 217426 131066
rect 306557 131066 306623 131069
rect 306557 131064 310040 131066
rect 306557 131008 306562 131064
rect 306618 131008 310040 131064
rect 306557 131006 310040 131008
rect 306557 131003 306623 131006
rect 252461 130930 252527 130933
rect 324313 130930 324379 130933
rect 248952 130928 252527 130930
rect 248952 130872 252466 130928
rect 252522 130872 252527 130928
rect 248952 130870 252527 130872
rect 321908 130928 324379 130930
rect 321908 130872 324318 130928
rect 324374 130872 324379 130928
rect 321908 130870 324379 130872
rect 252461 130867 252527 130870
rect 324313 130867 324379 130870
rect 495617 130794 495683 130797
rect 494316 130792 495683 130794
rect 494316 130736 495622 130792
rect 495678 130736 495683 130792
rect 494316 130734 495683 130736
rect 495617 130731 495683 130734
rect 306925 130658 306991 130661
rect 306925 130656 310040 130658
rect 214005 130114 214071 130117
rect 217182 130114 217242 130628
rect 306925 130600 306930 130656
rect 306986 130600 310040 130656
rect 306925 130598 310040 130600
rect 306925 130595 306991 130598
rect 252369 130522 252435 130525
rect 248952 130520 252435 130522
rect 248952 130464 252374 130520
rect 252430 130464 252435 130520
rect 248952 130462 252435 130464
rect 252369 130459 252435 130462
rect 309550 130146 310132 130206
rect 252461 130114 252527 130117
rect 214005 130112 217242 130114
rect 214005 130056 214010 130112
rect 214066 130056 217242 130112
rect 214005 130054 217242 130056
rect 248952 130112 252527 130114
rect 248952 130056 252466 130112
rect 252522 130056 252527 130112
rect 248952 130054 252527 130056
rect 214005 130051 214071 130054
rect 252461 130051 252527 130054
rect 260046 130052 260052 130116
rect 260116 130114 260122 130116
rect 309550 130114 309610 130146
rect 324405 130114 324471 130117
rect 260116 130054 309610 130114
rect 321908 130112 324471 130114
rect 321908 130056 324410 130112
rect 324466 130056 324471 130112
rect 321908 130054 324471 130056
rect 260116 130052 260122 130054
rect 324405 130051 324471 130054
rect 213913 129842 213979 129845
rect 213913 129840 216874 129842
rect 213913 129784 213918 129840
rect 213974 129784 216874 129840
rect 213913 129782 216874 129784
rect 213913 129779 213979 129782
rect 216814 129706 216874 129782
rect 217366 129706 217426 129948
rect 307477 129842 307543 129845
rect 307477 129840 310040 129842
rect 307477 129784 307482 129840
rect 307538 129784 310040 129840
rect 307477 129782 310040 129784
rect 307477 129779 307543 129782
rect 321553 129706 321619 129709
rect 496813 129706 496879 129709
rect 216814 129646 217426 129706
rect 321510 129704 321619 129706
rect 321510 129648 321558 129704
rect 321614 129648 321619 129704
rect 321510 129643 321619 129648
rect 494316 129704 496879 129706
rect 494316 129648 496818 129704
rect 496874 129648 496879 129704
rect 494316 129646 496879 129648
rect 496813 129643 496879 129646
rect 252461 129570 252527 129573
rect 248952 129568 252527 129570
rect 248952 129512 252466 129568
rect 252522 129512 252527 129568
rect 248952 129510 252527 129512
rect 252461 129507 252527 129510
rect 321510 129404 321570 129643
rect 419625 129570 419691 129573
rect 419625 129568 420164 129570
rect 419625 129512 419630 129568
rect 419686 129512 420164 129568
rect 419625 129510 420164 129512
rect 419625 129507 419691 129510
rect 67449 129298 67515 129301
rect 68142 129298 68816 129304
rect 67449 129296 68816 129298
rect 67449 129240 67454 129296
rect 67510 129244 68816 129296
rect 306925 129298 306991 129301
rect 306925 129296 310040 129298
rect 67510 129240 68202 129244
rect 67449 129238 68202 129240
rect 67449 129235 67515 129238
rect 213913 128890 213979 128893
rect 217182 128890 217242 129268
rect 306925 129240 306930 129296
rect 306986 129240 310040 129296
rect 306925 129238 310040 129240
rect 306925 129235 306991 129238
rect 252277 129162 252343 129165
rect 248952 129160 252343 129162
rect 248952 129104 252282 129160
rect 252338 129104 252343 129160
rect 248952 129102 252343 129104
rect 252277 129099 252343 129102
rect 494094 128964 494100 129028
rect 494164 128964 494170 129028
rect 213913 128888 217242 128890
rect 213913 128832 213918 128888
rect 213974 128832 217242 128888
rect 213913 128830 217242 128832
rect 307661 128890 307727 128893
rect 307661 128888 310040 128890
rect 307661 128832 307666 128888
rect 307722 128832 310040 128888
rect 307661 128830 310040 128832
rect 213913 128827 213979 128830
rect 307661 128827 307727 128830
rect 168966 128556 168972 128620
rect 169036 128618 169042 128620
rect 169036 128558 200130 128618
rect 169036 128556 169042 128558
rect 200070 128482 200130 128558
rect 217366 128482 217426 128724
rect 252369 128618 252435 128621
rect 324313 128618 324379 128621
rect 248952 128616 252435 128618
rect 248952 128560 252374 128616
rect 252430 128560 252435 128616
rect 248952 128558 252435 128560
rect 321908 128616 324379 128618
rect 321908 128560 324318 128616
rect 324374 128560 324379 128616
rect 321908 128558 324379 128560
rect 252369 128555 252435 128558
rect 324313 128555 324379 128558
rect 200070 128422 217426 128482
rect 307569 128482 307635 128485
rect 307569 128480 310040 128482
rect 307569 128424 307574 128480
rect 307630 128424 310040 128480
rect 494102 128452 494162 128964
rect 307569 128422 310040 128424
rect 307569 128419 307635 128422
rect 252277 128210 252343 128213
rect 248952 128208 252343 128210
rect 248952 128152 252282 128208
rect 252338 128152 252343 128208
rect 248952 128150 252343 128152
rect 252277 128147 252343 128150
rect 65517 128074 65583 128077
rect 68142 128074 68816 128080
rect 65517 128072 68816 128074
rect 65517 128016 65522 128072
rect 65578 128020 68816 128072
rect 307569 128074 307635 128077
rect 307569 128072 310040 128074
rect 65578 128016 68202 128020
rect 65517 128014 68202 128016
rect 65517 128011 65583 128014
rect 214005 127530 214071 127533
rect 217182 127530 217242 128044
rect 307569 128016 307574 128072
rect 307630 128016 310040 128072
rect 307569 128014 310040 128016
rect 307569 128011 307635 128014
rect 418705 127938 418771 127941
rect 419349 127938 419415 127941
rect 418705 127936 420164 127938
rect 418705 127880 418710 127936
rect 418766 127880 419354 127936
rect 419410 127880 420164 127936
rect 418705 127878 420164 127880
rect 418705 127875 418771 127878
rect 419349 127875 419415 127878
rect 324313 127802 324379 127805
rect 321908 127800 324379 127802
rect 321908 127744 324318 127800
rect 324374 127744 324379 127800
rect 321908 127742 324379 127744
rect 324313 127739 324379 127742
rect 252461 127666 252527 127669
rect 248952 127664 252527 127666
rect 248952 127608 252466 127664
rect 252522 127608 252527 127664
rect 248952 127606 252527 127608
rect 252461 127603 252527 127606
rect 307150 127604 307156 127668
rect 307220 127666 307226 127668
rect 307220 127606 310040 127666
rect 307220 127604 307226 127606
rect 214005 127528 217242 127530
rect 214005 127472 214010 127528
rect 214066 127472 217242 127528
rect 214005 127470 217242 127472
rect 214005 127467 214071 127470
rect 496813 127394 496879 127397
rect 494316 127392 496879 127394
rect 213913 127122 213979 127125
rect 217182 127122 217242 127364
rect 494316 127336 496818 127392
rect 496874 127336 496879 127392
rect 494316 127334 496879 127336
rect 496813 127331 496879 127334
rect 252369 127258 252435 127261
rect 248952 127256 252435 127258
rect 248952 127200 252374 127256
rect 252430 127200 252435 127256
rect 248952 127198 252435 127200
rect 252369 127195 252435 127198
rect 307661 127258 307727 127261
rect 307661 127256 310040 127258
rect 307661 127200 307666 127256
rect 307722 127200 310040 127256
rect 307661 127198 310040 127200
rect 307661 127195 307727 127198
rect 324405 127122 324471 127125
rect 213913 127120 217242 127122
rect 213913 127064 213918 127120
rect 213974 127064 217242 127120
rect 213913 127062 217242 127064
rect 321908 127120 324471 127122
rect 321908 127064 324410 127120
rect 324466 127064 324471 127120
rect 321908 127062 324471 127064
rect 213913 127059 213979 127062
rect 324405 127059 324471 127062
rect 307477 126850 307543 126853
rect 307477 126848 310040 126850
rect 307477 126792 307482 126848
rect 307538 126792 310040 126848
rect 307477 126790 310040 126792
rect 307477 126787 307543 126790
rect 252461 126714 252527 126717
rect 248952 126712 252527 126714
rect 67633 126306 67699 126309
rect 68142 126306 68816 126312
rect 67633 126304 68816 126306
rect 67633 126248 67638 126304
rect 67694 126252 68816 126304
rect 67694 126248 68202 126252
rect 67633 126246 68202 126248
rect 67633 126243 67699 126246
rect 214005 126170 214071 126173
rect 217182 126170 217242 126684
rect 248952 126656 252466 126712
rect 252522 126656 252527 126712
rect 248952 126654 252527 126656
rect 252461 126651 252527 126654
rect 307569 126442 307635 126445
rect 307569 126440 310040 126442
rect 307569 126384 307574 126440
rect 307630 126384 310040 126440
rect 307569 126382 310040 126384
rect 307569 126379 307635 126382
rect 252461 126306 252527 126309
rect 324497 126306 324563 126309
rect 496813 126306 496879 126309
rect 248952 126304 252527 126306
rect 248952 126248 252466 126304
rect 252522 126248 252527 126304
rect 248952 126246 252527 126248
rect 321908 126304 324563 126306
rect 321908 126248 324502 126304
rect 324558 126248 324563 126304
rect 321908 126246 324563 126248
rect 494316 126304 496879 126306
rect 494316 126248 496818 126304
rect 496874 126248 496879 126304
rect 494316 126246 496879 126248
rect 252461 126243 252527 126246
rect 324497 126243 324563 126246
rect 496813 126243 496879 126246
rect 214005 126168 217242 126170
rect 214005 126112 214010 126168
rect 214066 126112 217242 126168
rect 214005 126110 217242 126112
rect 418797 126170 418863 126173
rect 418797 126168 420164 126170
rect 418797 126112 418802 126168
rect 418858 126112 420164 126168
rect 418797 126110 420164 126112
rect 214005 126107 214071 126110
rect 418797 126107 418863 126110
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 213913 125762 213979 125765
rect 217182 125762 217242 126004
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 307661 125898 307727 125901
rect 307661 125896 310040 125898
rect 307661 125840 307666 125896
rect 307722 125840 310040 125896
rect 583520 125884 584960 125974
rect 307661 125838 310040 125840
rect 307661 125835 307727 125838
rect 251173 125762 251239 125765
rect 213913 125760 217242 125762
rect 213913 125704 213918 125760
rect 213974 125704 217242 125760
rect 213913 125702 217242 125704
rect 248952 125760 251239 125762
rect 248952 125704 251178 125760
rect 251234 125704 251239 125760
rect 248952 125702 251239 125704
rect 213913 125699 213979 125702
rect 251173 125699 251239 125702
rect 307477 125490 307543 125493
rect 324313 125490 324379 125493
rect 307477 125488 310040 125490
rect 307477 125432 307482 125488
rect 307538 125432 310040 125488
rect 307477 125430 310040 125432
rect 321908 125488 324379 125490
rect 321908 125432 324318 125488
rect 324374 125432 324379 125488
rect 321908 125430 324379 125432
rect 307477 125427 307543 125430
rect 324313 125427 324379 125430
rect 252093 125354 252159 125357
rect 248952 125352 252159 125354
rect 66161 125218 66227 125221
rect 68142 125218 68816 125224
rect 66161 125216 68816 125218
rect 66161 125160 66166 125216
rect 66222 125164 68816 125216
rect 66222 125160 68202 125164
rect 66161 125158 68202 125160
rect 66161 125155 66227 125158
rect 214005 124810 214071 124813
rect 217182 124810 217242 125324
rect 248952 125296 252098 125352
rect 252154 125296 252159 125352
rect 248952 125294 252159 125296
rect 252093 125291 252159 125294
rect 496813 125218 496879 125221
rect 494316 125216 496879 125218
rect 494316 125160 496818 125216
rect 496874 125160 496879 125216
rect 494316 125158 496879 125160
rect 496813 125155 496879 125158
rect 307569 125082 307635 125085
rect 307569 125080 310040 125082
rect 307569 125024 307574 125080
rect 307630 125024 310040 125080
rect 307569 125022 310040 125024
rect 307569 125019 307635 125022
rect 252461 124810 252527 124813
rect 324405 124810 324471 124813
rect 214005 124808 217242 124810
rect 214005 124752 214010 124808
rect 214066 124752 217242 124808
rect 214005 124750 217242 124752
rect 248952 124808 252527 124810
rect 248952 124752 252466 124808
rect 252522 124752 252527 124808
rect 248952 124750 252527 124752
rect 321908 124808 324471 124810
rect 321908 124752 324410 124808
rect 324466 124752 324471 124808
rect 321908 124750 324471 124752
rect 214005 124747 214071 124750
rect 252461 124747 252527 124750
rect 324405 124747 324471 124750
rect 307661 124674 307727 124677
rect 307661 124672 310040 124674
rect 213913 124402 213979 124405
rect 217182 124402 217242 124644
rect 307661 124616 307666 124672
rect 307722 124616 310040 124672
rect 307661 124614 310040 124616
rect 307661 124611 307727 124614
rect 419533 124538 419599 124541
rect 419533 124536 420164 124538
rect 419533 124480 419538 124536
rect 419594 124480 420164 124536
rect 419533 124478 420164 124480
rect 419533 124475 419599 124478
rect 252369 124402 252435 124405
rect 213913 124400 217242 124402
rect 213913 124344 213918 124400
rect 213974 124344 217242 124400
rect 213913 124342 217242 124344
rect 248952 124400 252435 124402
rect 248952 124344 252374 124400
rect 252430 124344 252435 124400
rect 248952 124342 252435 124344
rect 213913 124339 213979 124342
rect 252369 124339 252435 124342
rect 307293 124266 307359 124269
rect 307293 124264 310040 124266
rect 307293 124208 307298 124264
rect 307354 124208 310040 124264
rect 307293 124206 310040 124208
rect 307293 124203 307359 124206
rect 496905 124130 496971 124133
rect 494316 124128 496971 124130
rect -960 123572 480 123812
rect 66069 123586 66135 123589
rect 68142 123586 68816 123592
rect 66069 123584 68816 123586
rect 66069 123528 66074 123584
rect 66130 123532 68816 123584
rect 214005 123586 214071 123589
rect 217182 123586 217242 124100
rect 494316 124072 496910 124128
rect 496966 124072 496971 124128
rect 494316 124070 496971 124072
rect 496905 124067 496971 124070
rect 252185 123994 252251 123997
rect 324313 123994 324379 123997
rect 248952 123992 252251 123994
rect 248952 123936 252190 123992
rect 252246 123936 252251 123992
rect 248952 123934 252251 123936
rect 321908 123992 324379 123994
rect 321908 123936 324318 123992
rect 324374 123936 324379 123992
rect 321908 123934 324379 123936
rect 252185 123931 252251 123934
rect 324313 123931 324379 123934
rect 307569 123858 307635 123861
rect 307569 123856 310040 123858
rect 307569 123800 307574 123856
rect 307630 123800 310040 123856
rect 307569 123798 310040 123800
rect 307569 123795 307635 123798
rect 214005 123584 217242 123586
rect 66130 123528 68202 123532
rect 66069 123526 68202 123528
rect 214005 123528 214010 123584
rect 214066 123528 217242 123584
rect 214005 123526 217242 123528
rect 66069 123523 66135 123526
rect 214005 123523 214071 123526
rect 252461 123450 252527 123453
rect 308489 123450 308555 123453
rect 248952 123448 252527 123450
rect 213913 123178 213979 123181
rect 217182 123178 217242 123420
rect 248952 123392 252466 123448
rect 252522 123392 252527 123448
rect 248952 123390 252527 123392
rect 252461 123387 252527 123390
rect 258030 123448 308555 123450
rect 258030 123392 308494 123448
rect 308550 123392 308555 123448
rect 258030 123390 308555 123392
rect 251950 123252 251956 123316
rect 252020 123314 252026 123316
rect 258030 123314 258090 123390
rect 308489 123387 308555 123390
rect 309550 123346 310132 123406
rect 252020 123254 258090 123314
rect 305913 123314 305979 123317
rect 309550 123314 309610 123346
rect 305913 123312 309610 123314
rect 305913 123256 305918 123312
rect 305974 123256 309610 123312
rect 305913 123254 309610 123256
rect 252020 123252 252026 123254
rect 305913 123251 305979 123254
rect 324405 123178 324471 123181
rect 213913 123176 217242 123178
rect 213913 123120 213918 123176
rect 213974 123120 217242 123176
rect 213913 123118 217242 123120
rect 321908 123176 324471 123178
rect 321908 123120 324410 123176
rect 324466 123120 324471 123176
rect 321908 123118 324471 123120
rect 213913 123115 213979 123118
rect 324405 123115 324471 123118
rect 252277 123042 252343 123045
rect 248952 123040 252343 123042
rect 248952 122984 252282 123040
rect 252338 122984 252343 123040
rect 248952 122982 252343 122984
rect 252277 122979 252343 122982
rect 307661 123042 307727 123045
rect 307661 123040 310040 123042
rect 307661 122984 307666 123040
rect 307722 122984 310040 123040
rect 307661 122982 310040 122984
rect 307661 122979 307727 122982
rect 496813 122906 496879 122909
rect 494316 122904 496879 122906
rect 494316 122848 496818 122904
rect 496874 122848 496879 122904
rect 494316 122846 496879 122848
rect 496813 122843 496879 122846
rect 416773 122770 416839 122773
rect 416773 122768 420164 122770
rect 67357 122634 67423 122637
rect 68142 122634 68816 122640
rect 67357 122632 68816 122634
rect 67357 122576 67362 122632
rect 67418 122580 68816 122632
rect 67418 122576 68202 122580
rect 67357 122574 68202 122576
rect 67357 122571 67423 122574
rect 214005 122226 214071 122229
rect 217182 122226 217242 122740
rect 416773 122712 416778 122768
rect 416834 122712 420164 122768
rect 416773 122710 420164 122712
rect 416773 122707 416839 122710
rect 252461 122498 252527 122501
rect 248952 122496 252527 122498
rect 248952 122440 252466 122496
rect 252522 122440 252527 122496
rect 248952 122438 252527 122440
rect 252461 122435 252527 122438
rect 307477 122498 307543 122501
rect 324313 122498 324379 122501
rect 307477 122496 310040 122498
rect 307477 122440 307482 122496
rect 307538 122440 310040 122496
rect 307477 122438 310040 122440
rect 321908 122496 324379 122498
rect 321908 122440 324318 122496
rect 324374 122440 324379 122496
rect 321908 122438 324379 122440
rect 307477 122435 307543 122438
rect 324313 122435 324379 122438
rect 214005 122224 217242 122226
rect 214005 122168 214010 122224
rect 214066 122168 217242 122224
rect 214005 122166 217242 122168
rect 214005 122163 214071 122166
rect 252369 122090 252435 122093
rect 248952 122088 252435 122090
rect 213913 121546 213979 121549
rect 217182 121546 217242 122060
rect 248952 122032 252374 122088
rect 252430 122032 252435 122088
rect 248952 122030 252435 122032
rect 252369 122027 252435 122030
rect 307661 122090 307727 122093
rect 307661 122088 310040 122090
rect 307661 122032 307666 122088
rect 307722 122032 310040 122088
rect 307661 122030 310040 122032
rect 307661 122027 307727 122030
rect 496813 121818 496879 121821
rect 494316 121816 496879 121818
rect 494316 121760 496818 121816
rect 496874 121760 496879 121816
rect 494316 121758 496879 121760
rect 496813 121755 496879 121758
rect 307569 121682 307635 121685
rect 324405 121682 324471 121685
rect 307569 121680 310040 121682
rect 307569 121624 307574 121680
rect 307630 121624 310040 121680
rect 307569 121622 310040 121624
rect 321908 121680 324471 121682
rect 321908 121624 324410 121680
rect 324466 121624 324471 121680
rect 321908 121622 324471 121624
rect 307569 121619 307635 121622
rect 324405 121619 324471 121622
rect 252277 121546 252343 121549
rect 213913 121544 217242 121546
rect 213913 121488 213918 121544
rect 213974 121488 217242 121544
rect 213913 121486 217242 121488
rect 248952 121544 252343 121546
rect 248952 121488 252282 121544
rect 252338 121488 252343 121544
rect 248952 121486 252343 121488
rect 213913 121483 213979 121486
rect 252277 121483 252343 121486
rect 65149 120866 65215 120869
rect 68142 120866 68816 120872
rect 65149 120864 68816 120866
rect 65149 120808 65154 120864
rect 65210 120812 68816 120864
rect 214005 120866 214071 120869
rect 217182 120866 217242 121380
rect 307477 121274 307543 121277
rect 307477 121272 310040 121274
rect 307477 121216 307482 121272
rect 307538 121216 310040 121272
rect 307477 121214 310040 121216
rect 307477 121211 307543 121214
rect 251909 121138 251975 121141
rect 248952 121136 251975 121138
rect 248952 121080 251914 121136
rect 251970 121080 251975 121136
rect 248952 121078 251975 121080
rect 251909 121075 251975 121078
rect 416773 121138 416839 121141
rect 416773 121136 420164 121138
rect 416773 121080 416778 121136
rect 416834 121080 420164 121136
rect 416773 121078 420164 121080
rect 416773 121075 416839 121078
rect 214005 120864 217242 120866
rect 65210 120808 68202 120812
rect 65149 120806 68202 120808
rect 214005 120808 214010 120864
rect 214066 120808 217242 120864
rect 214005 120806 217242 120808
rect 307661 120866 307727 120869
rect 324957 120866 325023 120869
rect 307661 120864 310040 120866
rect 307661 120808 307666 120864
rect 307722 120808 310040 120864
rect 307661 120806 310040 120808
rect 321908 120864 325023 120866
rect 321908 120808 324962 120864
rect 325018 120808 325023 120864
rect 321908 120806 325023 120808
rect 65149 120803 65215 120806
rect 214005 120803 214071 120806
rect 307661 120803 307727 120806
rect 324957 120803 325023 120806
rect 498377 120730 498443 120733
rect 494316 120728 498443 120730
rect 213913 120186 213979 120189
rect 217182 120186 217242 120700
rect 494316 120672 498382 120728
rect 498438 120672 498443 120728
rect 494316 120670 498443 120672
rect 498377 120667 498443 120670
rect 252461 120594 252527 120597
rect 248952 120592 252527 120594
rect 248952 120536 252466 120592
rect 252522 120536 252527 120592
rect 248952 120534 252527 120536
rect 252461 120531 252527 120534
rect 307569 120458 307635 120461
rect 307569 120456 310040 120458
rect 307569 120400 307574 120456
rect 307630 120400 310040 120456
rect 307569 120398 310040 120400
rect 307569 120395 307635 120398
rect 252461 120186 252527 120189
rect 324313 120186 324379 120189
rect 213913 120184 217242 120186
rect 213913 120128 213918 120184
rect 213974 120128 217242 120184
rect 213913 120126 217242 120128
rect 248952 120184 252527 120186
rect 248952 120128 252466 120184
rect 252522 120128 252527 120184
rect 248952 120126 252527 120128
rect 321908 120184 324379 120186
rect 321908 120128 324318 120184
rect 324374 120128 324379 120184
rect 321908 120126 324379 120128
rect 213913 120123 213979 120126
rect 252461 120123 252527 120126
rect 324313 120123 324379 120126
rect 307477 120050 307543 120053
rect 307477 120048 310040 120050
rect 214005 119642 214071 119645
rect 217182 119642 217242 120020
rect 307477 119992 307482 120048
rect 307538 119992 310040 120048
rect 307477 119990 310040 119992
rect 307477 119987 307543 119990
rect 252461 119642 252527 119645
rect 214005 119640 217242 119642
rect 214005 119584 214010 119640
rect 214066 119584 217242 119640
rect 214005 119582 217242 119584
rect 248952 119640 252527 119642
rect 248952 119584 252466 119640
rect 252522 119584 252527 119640
rect 248952 119582 252527 119584
rect 214005 119579 214071 119582
rect 252461 119579 252527 119582
rect 307569 119642 307635 119645
rect 495433 119642 495499 119645
rect 307569 119640 310040 119642
rect 307569 119584 307574 119640
rect 307630 119584 310040 119640
rect 307569 119582 310040 119584
rect 494316 119640 495499 119642
rect 494316 119584 495438 119640
rect 495494 119584 495499 119640
rect 494316 119582 495499 119584
rect 307569 119579 307635 119582
rect 495433 119579 495499 119582
rect 213453 119098 213519 119101
rect 217182 119098 217242 119476
rect 324313 119370 324379 119373
rect 321908 119368 324379 119370
rect 321908 119312 324318 119368
rect 324374 119312 324379 119368
rect 321908 119310 324379 119312
rect 324313 119307 324379 119310
rect 417417 119370 417483 119373
rect 417417 119368 420164 119370
rect 417417 119312 417422 119368
rect 417478 119312 420164 119368
rect 417417 119310 420164 119312
rect 417417 119307 417483 119310
rect 252461 119234 252527 119237
rect 248952 119232 252527 119234
rect 248952 119176 252466 119232
rect 252522 119176 252527 119232
rect 248952 119174 252527 119176
rect 252461 119171 252527 119174
rect 213453 119096 217242 119098
rect 213453 119040 213458 119096
rect 213514 119040 217242 119096
rect 213453 119038 217242 119040
rect 307661 119098 307727 119101
rect 307661 119096 310040 119098
rect 307661 119040 307666 119096
rect 307722 119040 310040 119096
rect 307661 119038 310040 119040
rect 213453 119035 213519 119038
rect 307661 119035 307727 119038
rect 213913 118962 213979 118965
rect 213913 118960 217242 118962
rect 213913 118904 213918 118960
rect 213974 118904 217242 118960
rect 213913 118902 217242 118904
rect 213913 118899 213979 118902
rect 217182 118796 217242 118902
rect 251725 118826 251791 118829
rect 248952 118824 251791 118826
rect 248952 118768 251730 118824
rect 251786 118768 251791 118824
rect 248952 118766 251791 118768
rect 251725 118763 251791 118766
rect 305729 118826 305795 118829
rect 307569 118826 307635 118829
rect 305729 118824 307635 118826
rect 305729 118768 305734 118824
rect 305790 118768 307574 118824
rect 307630 118768 307635 118824
rect 305729 118766 307635 118768
rect 305729 118763 305795 118766
rect 307569 118763 307635 118766
rect 306557 118690 306623 118693
rect 306557 118688 310040 118690
rect 306557 118632 306562 118688
rect 306618 118632 310040 118688
rect 306557 118630 310040 118632
rect 306557 118627 306623 118630
rect 324313 118554 324379 118557
rect 321908 118552 324379 118554
rect 321908 118496 324318 118552
rect 324374 118496 324379 118552
rect 321908 118494 324379 118496
rect 324313 118491 324379 118494
rect 496813 118418 496879 118421
rect 494316 118416 496879 118418
rect 494316 118360 496818 118416
rect 496874 118360 496879 118416
rect 494316 118358 496879 118360
rect 496813 118355 496879 118358
rect 252461 118282 252527 118285
rect 248952 118280 252527 118282
rect 248952 118224 252466 118280
rect 252522 118224 252527 118280
rect 248952 118222 252527 118224
rect 252461 118219 252527 118222
rect 309550 118178 310132 118238
rect 214005 117602 214071 117605
rect 217182 117602 217242 118116
rect 302734 118084 302740 118148
rect 302804 118146 302810 118148
rect 309550 118146 309610 118178
rect 302804 118086 309610 118146
rect 302804 118084 302810 118086
rect 252369 117874 252435 117877
rect 248952 117872 252435 117874
rect 248952 117816 252374 117872
rect 252430 117816 252435 117872
rect 248952 117814 252435 117816
rect 252369 117811 252435 117814
rect 307569 117874 307635 117877
rect 324405 117874 324471 117877
rect 307569 117872 310040 117874
rect 307569 117816 307574 117872
rect 307630 117816 310040 117872
rect 307569 117814 310040 117816
rect 321908 117872 324471 117874
rect 321908 117816 324410 117872
rect 324466 117816 324471 117872
rect 321908 117814 324471 117816
rect 307569 117811 307635 117814
rect 324405 117811 324471 117814
rect 416773 117738 416839 117741
rect 416773 117736 420164 117738
rect 416773 117680 416778 117736
rect 416834 117680 420164 117736
rect 416773 117678 420164 117680
rect 416773 117675 416839 117678
rect 214005 117600 217242 117602
rect 214005 117544 214010 117600
rect 214066 117544 217242 117600
rect 214005 117542 217242 117544
rect 214005 117539 214071 117542
rect 307661 117466 307727 117469
rect 307661 117464 310040 117466
rect 213913 117330 213979 117333
rect 213913 117328 216874 117330
rect 213913 117272 213918 117328
rect 213974 117272 216874 117328
rect 213913 117270 216874 117272
rect 213913 117267 213979 117270
rect 216814 117194 216874 117270
rect 217366 117194 217426 117436
rect 307661 117408 307666 117464
rect 307722 117408 310040 117464
rect 307661 117406 310040 117408
rect 307661 117403 307727 117406
rect 251817 117330 251883 117333
rect 496905 117330 496971 117333
rect 248952 117328 251883 117330
rect 248952 117272 251822 117328
rect 251878 117272 251883 117328
rect 248952 117270 251883 117272
rect 494316 117328 496971 117330
rect 494316 117272 496910 117328
rect 496966 117272 496971 117328
rect 494316 117270 496971 117272
rect 251817 117267 251883 117270
rect 496905 117267 496971 117270
rect 216814 117134 217426 117194
rect 307569 117058 307635 117061
rect 324313 117058 324379 117061
rect 307569 117056 310040 117058
rect 307569 117000 307574 117056
rect 307630 117000 310040 117056
rect 307569 116998 310040 117000
rect 321908 117056 324379 117058
rect 321908 117000 324318 117056
rect 324374 117000 324379 117056
rect 321908 116998 324379 117000
rect 307569 116995 307635 116998
rect 324313 116995 324379 116998
rect 252369 116922 252435 116925
rect 248952 116920 252435 116922
rect 248952 116864 252374 116920
rect 252430 116864 252435 116920
rect 248952 116862 252435 116864
rect 252369 116859 252435 116862
rect 214005 116242 214071 116245
rect 217182 116242 217242 116756
rect 306741 116650 306807 116653
rect 306741 116648 310040 116650
rect 306741 116592 306746 116648
rect 306802 116592 310040 116648
rect 306741 116590 310040 116592
rect 306741 116587 306807 116590
rect 252461 116378 252527 116381
rect 324405 116378 324471 116381
rect 248952 116376 252527 116378
rect 248952 116320 252466 116376
rect 252522 116320 252527 116376
rect 248952 116318 252527 116320
rect 321908 116376 324471 116378
rect 321908 116320 324410 116376
rect 324466 116320 324471 116376
rect 321908 116318 324471 116320
rect 252461 116315 252527 116318
rect 324405 116315 324471 116318
rect 214005 116240 217242 116242
rect 214005 116184 214010 116240
rect 214066 116184 217242 116240
rect 214005 116182 217242 116184
rect 307661 116242 307727 116245
rect 496813 116242 496879 116245
rect 307661 116240 310040 116242
rect 307661 116184 307666 116240
rect 307722 116184 310040 116240
rect 307661 116182 310040 116184
rect 494316 116240 496879 116242
rect 494316 116184 496818 116240
rect 496874 116184 496879 116240
rect 494316 116182 496879 116184
rect 214005 116179 214071 116182
rect 307661 116179 307727 116182
rect 496813 116179 496879 116182
rect 416773 116106 416839 116109
rect 416773 116104 420164 116106
rect 213913 115970 213979 115973
rect 213913 115968 216874 115970
rect 213913 115912 213918 115968
rect 213974 115912 216874 115968
rect 213913 115910 216874 115912
rect 213913 115907 213979 115910
rect 216814 115834 216874 115910
rect 217366 115834 217426 116076
rect 416773 116048 416778 116104
rect 416834 116048 420164 116104
rect 416773 116046 420164 116048
rect 416773 116043 416839 116046
rect 252277 115970 252343 115973
rect 248952 115968 252343 115970
rect 248952 115912 252282 115968
rect 252338 115912 252343 115968
rect 248952 115910 252343 115912
rect 252277 115907 252343 115910
rect 216814 115774 217426 115834
rect 307477 115698 307543 115701
rect 307477 115696 310040 115698
rect 307477 115640 307482 115696
rect 307538 115640 310040 115696
rect 307477 115638 310040 115640
rect 307477 115635 307543 115638
rect 324313 115562 324379 115565
rect 321908 115560 324379 115562
rect 321908 115504 324318 115560
rect 324374 115504 324379 115560
rect 321908 115502 324379 115504
rect 324313 115499 324379 115502
rect 252461 115426 252527 115429
rect 248952 115424 252527 115426
rect 213913 115018 213979 115021
rect 217182 115018 217242 115396
rect 248952 115368 252466 115424
rect 252522 115368 252527 115424
rect 248952 115366 252527 115368
rect 252461 115363 252527 115366
rect 307569 115290 307635 115293
rect 307569 115288 310040 115290
rect 307569 115232 307574 115288
rect 307630 115232 310040 115288
rect 307569 115230 310040 115232
rect 307569 115227 307635 115230
rect 497457 115154 497523 115157
rect 494316 115152 497523 115154
rect 494316 115096 497462 115152
rect 497518 115096 497523 115152
rect 494316 115094 497523 115096
rect 497457 115091 497523 115094
rect 252369 115018 252435 115021
rect 213913 115016 217242 115018
rect 213913 114960 213918 115016
rect 213974 114960 217242 115016
rect 213913 114958 217242 114960
rect 248952 115016 252435 115018
rect 248952 114960 252374 115016
rect 252430 114960 252435 115016
rect 248952 114958 252435 114960
rect 213913 114955 213979 114958
rect 252369 114955 252435 114958
rect 307661 114882 307727 114885
rect 307661 114880 310040 114882
rect 216673 114610 216739 114613
rect 217182 114610 217242 114852
rect 307661 114824 307666 114880
rect 307722 114824 310040 114880
rect 307661 114822 310040 114824
rect 307661 114819 307727 114822
rect 324405 114746 324471 114749
rect 321908 114744 324471 114746
rect 321908 114688 324410 114744
rect 324466 114688 324471 114744
rect 321908 114686 324471 114688
rect 324405 114683 324471 114686
rect 216673 114608 217242 114610
rect 216673 114552 216678 114608
rect 216734 114552 217242 114608
rect 216673 114550 217242 114552
rect 216673 114547 216739 114550
rect 251766 114474 251772 114476
rect 248952 114414 251772 114474
rect 251766 114412 251772 114414
rect 251836 114412 251842 114476
rect 307661 114474 307727 114477
rect 307661 114472 310040 114474
rect 307661 114416 307666 114472
rect 307722 114416 310040 114472
rect 307661 114414 310040 114416
rect 307661 114411 307727 114414
rect 416773 114338 416839 114341
rect 416773 114336 420164 114338
rect 416773 114280 416778 114336
rect 416834 114280 420164 114336
rect 416773 114278 420164 114280
rect 416773 114275 416839 114278
rect 214005 113658 214071 113661
rect 217182 113658 217242 114172
rect 252461 114066 252527 114069
rect 248952 114064 252527 114066
rect 248952 114008 252466 114064
rect 252522 114008 252527 114064
rect 248952 114006 252527 114008
rect 252461 114003 252527 114006
rect 307109 114066 307175 114069
rect 324313 114066 324379 114069
rect 307109 114064 310040 114066
rect 307109 114008 307114 114064
rect 307170 114008 310040 114064
rect 307109 114006 310040 114008
rect 321908 114064 324379 114066
rect 321908 114008 324318 114064
rect 324374 114008 324379 114064
rect 321908 114006 324379 114008
rect 307109 114003 307175 114006
rect 324313 114003 324379 114006
rect 496813 113930 496879 113933
rect 494316 113928 496879 113930
rect 494316 113872 496818 113928
rect 496874 113872 496879 113928
rect 494316 113870 496879 113872
rect 496813 113867 496879 113870
rect 214005 113656 217242 113658
rect 214005 113600 214010 113656
rect 214066 113600 217242 113656
rect 214005 113598 217242 113600
rect 307569 113658 307635 113661
rect 307569 113656 310040 113658
rect 307569 113600 307574 113656
rect 307630 113600 310040 113656
rect 307569 113598 310040 113600
rect 214005 113595 214071 113598
rect 307569 113595 307635 113598
rect 252369 113522 252435 113525
rect 248952 113520 252435 113522
rect 213913 113250 213979 113253
rect 217182 113250 217242 113492
rect 248952 113464 252374 113520
rect 252430 113464 252435 113520
rect 248952 113462 252435 113464
rect 252369 113459 252435 113462
rect 213913 113248 217242 113250
rect 213913 113192 213918 113248
rect 213974 113192 217242 113248
rect 213913 113190 217242 113192
rect 307661 113250 307727 113253
rect 324405 113250 324471 113253
rect 307661 113248 310040 113250
rect 307661 113192 307666 113248
rect 307722 113192 310040 113248
rect 307661 113190 310040 113192
rect 321908 113248 324471 113250
rect 321908 113192 324410 113248
rect 324466 113192 324471 113248
rect 321908 113190 324471 113192
rect 213913 113187 213979 113190
rect 307661 113187 307727 113190
rect 324405 113187 324471 113190
rect 252093 113114 252159 113117
rect 248952 113112 252159 113114
rect 248952 113056 252098 113112
rect 252154 113056 252159 113112
rect 248952 113054 252159 113056
rect 252093 113051 252159 113054
rect 496905 112842 496971 112845
rect 494316 112840 496971 112842
rect 214005 112298 214071 112301
rect 217182 112298 217242 112812
rect 494316 112784 496910 112840
rect 496966 112784 496971 112840
rect 494316 112782 496971 112784
rect 496905 112779 496971 112782
rect 580257 112842 580323 112845
rect 583520 112842 584960 112932
rect 580257 112840 584960 112842
rect 580257 112784 580262 112840
rect 580318 112784 584960 112840
rect 580257 112782 584960 112784
rect 580257 112779 580323 112782
rect 252461 112706 252527 112709
rect 248952 112704 252527 112706
rect 248952 112648 252466 112704
rect 252522 112648 252527 112704
rect 248952 112646 252527 112648
rect 252461 112643 252527 112646
rect 306925 112706 306991 112709
rect 416773 112706 416839 112709
rect 306925 112704 310040 112706
rect 306925 112648 306930 112704
rect 306986 112648 310040 112704
rect 306925 112646 310040 112648
rect 416773 112704 420164 112706
rect 416773 112648 416778 112704
rect 416834 112648 420164 112704
rect 583520 112692 584960 112782
rect 416773 112646 420164 112648
rect 306925 112643 306991 112646
rect 416773 112643 416839 112646
rect 324313 112434 324379 112437
rect 321908 112432 324379 112434
rect 321908 112376 324318 112432
rect 324374 112376 324379 112432
rect 321908 112374 324379 112376
rect 324313 112371 324379 112374
rect 214005 112296 217242 112298
rect 214005 112240 214010 112296
rect 214066 112240 217242 112296
rect 214005 112238 217242 112240
rect 309133 112298 309199 112301
rect 309133 112296 310040 112298
rect 309133 112240 309138 112296
rect 309194 112240 310040 112296
rect 309133 112238 310040 112240
rect 214005 112235 214071 112238
rect 309133 112235 309199 112238
rect 252461 112162 252527 112165
rect 248952 112160 252527 112162
rect 213913 111890 213979 111893
rect 217366 111890 217426 112132
rect 248952 112104 252466 112160
rect 252522 112104 252527 112160
rect 248952 112102 252527 112104
rect 252461 112099 252527 112102
rect 213913 111888 217426 111890
rect 213913 111832 213918 111888
rect 213974 111832 217426 111888
rect 213913 111830 217426 111832
rect 307661 111890 307727 111893
rect 307661 111888 310040 111890
rect 307661 111832 307666 111888
rect 307722 111832 310040 111888
rect 307661 111830 310040 111832
rect 213913 111827 213979 111830
rect 307661 111827 307727 111830
rect 167913 111754 167979 111757
rect 252277 111754 252343 111757
rect 324313 111754 324379 111757
rect 496813 111754 496879 111757
rect 164694 111752 167979 111754
rect 164694 111696 167918 111752
rect 167974 111696 167979 111752
rect 164694 111694 167979 111696
rect 248952 111752 252343 111754
rect 248952 111696 252282 111752
rect 252338 111696 252343 111752
rect 248952 111694 252343 111696
rect 321908 111752 324379 111754
rect 321908 111696 324318 111752
rect 324374 111696 324379 111752
rect 321908 111694 324379 111696
rect 494316 111752 496879 111754
rect 494316 111696 496818 111752
rect 496874 111696 496879 111752
rect 494316 111694 496879 111696
rect 167913 111691 167979 111694
rect 252277 111691 252343 111694
rect 324313 111691 324379 111694
rect 496813 111691 496879 111694
rect 307477 111482 307543 111485
rect 307477 111480 310040 111482
rect 214005 110938 214071 110941
rect 217182 110938 217242 111452
rect 307477 111424 307482 111480
rect 307538 111424 310040 111480
rect 307477 111422 310040 111424
rect 307477 111419 307543 111422
rect 252369 111210 252435 111213
rect 248952 111208 252435 111210
rect 248952 111152 252374 111208
rect 252430 111152 252435 111208
rect 248952 111150 252435 111152
rect 252369 111147 252435 111150
rect 307569 111074 307635 111077
rect 307569 111072 310040 111074
rect 307569 111016 307574 111072
rect 307630 111016 310040 111072
rect 307569 111014 310040 111016
rect 307569 111011 307635 111014
rect 324405 110938 324471 110941
rect 214005 110936 217242 110938
rect 214005 110880 214010 110936
rect 214066 110880 217242 110936
rect 214005 110878 217242 110880
rect 321908 110936 324471 110938
rect 321908 110880 324410 110936
rect 324466 110880 324471 110936
rect 321908 110878 324471 110880
rect 214005 110875 214071 110878
rect 324405 110875 324471 110878
rect 416773 110938 416839 110941
rect 416773 110936 420164 110938
rect 416773 110880 416778 110936
rect 416834 110880 420164 110936
rect 416773 110878 420164 110880
rect 416773 110875 416839 110878
rect 252461 110802 252527 110805
rect 248952 110800 252527 110802
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 213913 110530 213979 110533
rect 217366 110530 217426 110772
rect 248952 110744 252466 110800
rect 252522 110744 252527 110800
rect 248952 110742 252527 110744
rect 252461 110739 252527 110742
rect 307661 110666 307727 110669
rect 496813 110666 496879 110669
rect 307661 110664 310040 110666
rect 307661 110608 307666 110664
rect 307722 110608 310040 110664
rect 307661 110606 310040 110608
rect 494316 110664 496879 110666
rect 494316 110608 496818 110664
rect 496874 110608 496879 110664
rect 494316 110606 496879 110608
rect 307661 110603 307727 110606
rect 496813 110603 496879 110606
rect 213913 110528 217426 110530
rect 213913 110472 213918 110528
rect 213974 110472 217426 110528
rect 213913 110470 217426 110472
rect 213913 110467 213979 110470
rect 252461 110258 252527 110261
rect 248952 110256 252527 110258
rect 167729 110122 167795 110125
rect 164694 110120 167795 110122
rect 164694 110064 167734 110120
rect 167790 110064 167795 110120
rect 164694 110062 167795 110064
rect 167729 110059 167795 110062
rect 214005 109714 214071 109717
rect 217182 109714 217242 110228
rect 248952 110200 252466 110256
rect 252522 110200 252527 110256
rect 248952 110198 252527 110200
rect 252461 110195 252527 110198
rect 306741 110258 306807 110261
rect 306741 110256 310040 110258
rect 306741 110200 306746 110256
rect 306802 110200 310040 110256
rect 306741 110198 310040 110200
rect 306741 110195 306807 110198
rect 324497 110122 324563 110125
rect 321908 110120 324563 110122
rect 321908 110064 324502 110120
rect 324558 110064 324563 110120
rect 321908 110062 324563 110064
rect 324497 110059 324563 110062
rect 252369 109850 252435 109853
rect 248952 109848 252435 109850
rect 248952 109792 252374 109848
rect 252430 109792 252435 109848
rect 248952 109790 252435 109792
rect 252369 109787 252435 109790
rect 307661 109850 307727 109853
rect 307661 109848 310040 109850
rect 307661 109792 307666 109848
rect 307722 109792 310040 109848
rect 307661 109790 310040 109792
rect 307661 109787 307727 109790
rect 214005 109712 217242 109714
rect 214005 109656 214010 109712
rect 214066 109656 217242 109712
rect 214005 109654 217242 109656
rect 214005 109651 214071 109654
rect 213913 109170 213979 109173
rect 217182 109170 217242 109548
rect 324313 109442 324379 109445
rect 496813 109442 496879 109445
rect 321908 109440 324379 109442
rect 321908 109384 324318 109440
rect 324374 109384 324379 109440
rect 321908 109382 324379 109384
rect 494316 109440 496879 109442
rect 494316 109384 496818 109440
rect 496874 109384 496879 109440
rect 494316 109382 496879 109384
rect 324313 109379 324379 109382
rect 496813 109379 496879 109382
rect 252277 109306 252343 109309
rect 248952 109304 252343 109306
rect 248952 109248 252282 109304
rect 252338 109248 252343 109304
rect 248952 109246 252343 109248
rect 252277 109243 252343 109246
rect 305637 109306 305703 109309
rect 306741 109306 306807 109309
rect 305637 109304 306807 109306
rect 305637 109248 305642 109304
rect 305698 109248 306746 109304
rect 306802 109248 306807 109304
rect 305637 109246 306807 109248
rect 305637 109243 305703 109246
rect 306741 109243 306807 109246
rect 306925 109306 306991 109309
rect 416773 109306 416839 109309
rect 306925 109304 310040 109306
rect 306925 109248 306930 109304
rect 306986 109248 310040 109304
rect 306925 109246 310040 109248
rect 416773 109304 420164 109306
rect 416773 109248 416778 109304
rect 416834 109248 420164 109304
rect 416773 109246 420164 109248
rect 306925 109243 306991 109246
rect 416773 109243 416839 109246
rect 213913 109168 217242 109170
rect 213913 109112 213918 109168
rect 213974 109112 217242 109168
rect 213913 109110 217242 109112
rect 213913 109107 213979 109110
rect 252461 108898 252527 108901
rect 248952 108896 252527 108898
rect 168097 108762 168163 108765
rect 164694 108760 168163 108762
rect 164694 108704 168102 108760
rect 168158 108704 168163 108760
rect 164694 108702 168163 108704
rect 168097 108699 168163 108702
rect 214005 108354 214071 108357
rect 217182 108354 217242 108868
rect 248952 108840 252466 108896
rect 252522 108840 252527 108896
rect 248952 108838 252527 108840
rect 252461 108835 252527 108838
rect 307569 108898 307635 108901
rect 307569 108896 310040 108898
rect 307569 108840 307574 108896
rect 307630 108840 310040 108896
rect 307569 108838 310040 108840
rect 307569 108835 307635 108838
rect 324589 108626 324655 108629
rect 321908 108624 324655 108626
rect 321908 108568 324594 108624
rect 324650 108568 324655 108624
rect 321908 108566 324655 108568
rect 324589 108563 324655 108566
rect 309550 108386 310132 108446
rect 252185 108354 252251 108357
rect 214005 108352 217242 108354
rect 214005 108296 214010 108352
rect 214066 108296 217242 108352
rect 214005 108294 217242 108296
rect 248952 108352 252251 108354
rect 248952 108296 252190 108352
rect 252246 108296 252251 108352
rect 248952 108294 252251 108296
rect 214005 108291 214071 108294
rect 252185 108291 252251 108294
rect 305821 108354 305887 108357
rect 309550 108354 309610 108386
rect 496997 108354 497063 108357
rect 305821 108352 309610 108354
rect 305821 108296 305826 108352
rect 305882 108296 309610 108352
rect 305821 108294 309610 108296
rect 494316 108352 497063 108354
rect 494316 108296 497002 108352
rect 497058 108296 497063 108352
rect 494316 108294 497063 108296
rect 305821 108291 305887 108294
rect 496997 108291 497063 108294
rect 213913 107946 213979 107949
rect 217182 107946 217242 108188
rect 307661 108082 307727 108085
rect 307661 108080 310040 108082
rect 307661 108024 307666 108080
rect 307722 108024 310040 108080
rect 307661 108022 310040 108024
rect 307661 108019 307727 108022
rect 251725 107946 251791 107949
rect 213913 107944 217242 107946
rect 213913 107888 213918 107944
rect 213974 107888 217242 107944
rect 213913 107886 217242 107888
rect 248952 107944 251791 107946
rect 248952 107888 251730 107944
rect 251786 107888 251791 107944
rect 248952 107886 251791 107888
rect 213913 107883 213979 107886
rect 251725 107883 251791 107886
rect 324313 107810 324379 107813
rect 321908 107808 324379 107810
rect 321908 107752 324318 107808
rect 324374 107752 324379 107808
rect 321908 107750 324379 107752
rect 324313 107747 324379 107750
rect 307661 107674 307727 107677
rect 307661 107672 310040 107674
rect 307661 107616 307666 107672
rect 307722 107616 310040 107672
rect 307661 107614 310040 107616
rect 307661 107611 307727 107614
rect 252461 107538 252527 107541
rect 248952 107536 252527 107538
rect 214005 106994 214071 106997
rect 217182 106994 217242 107508
rect 248952 107480 252466 107536
rect 252522 107480 252527 107536
rect 248952 107478 252527 107480
rect 252461 107475 252527 107478
rect 416773 107538 416839 107541
rect 416773 107536 420164 107538
rect 416773 107480 416778 107536
rect 416834 107480 420164 107536
rect 416773 107478 420164 107480
rect 416773 107475 416839 107478
rect 307569 107266 307635 107269
rect 496813 107266 496879 107269
rect 307569 107264 310040 107266
rect 307569 107208 307574 107264
rect 307630 107208 310040 107264
rect 307569 107206 310040 107208
rect 494316 107264 496879 107266
rect 494316 107208 496818 107264
rect 496874 107208 496879 107264
rect 494316 107206 496879 107208
rect 307569 107203 307635 107206
rect 496813 107203 496879 107206
rect 324313 107130 324379 107133
rect 321908 107128 324379 107130
rect 321908 107072 324318 107128
rect 324374 107072 324379 107128
rect 321908 107070 324379 107072
rect 324313 107067 324379 107070
rect 252093 106994 252159 106997
rect 214005 106992 217242 106994
rect 214005 106936 214010 106992
rect 214066 106936 217242 106992
rect 214005 106934 217242 106936
rect 248952 106992 252159 106994
rect 248952 106936 252098 106992
rect 252154 106936 252159 106992
rect 248952 106934 252159 106936
rect 214005 106931 214071 106934
rect 252093 106931 252159 106934
rect 307477 106858 307543 106861
rect 307477 106856 310040 106858
rect 213913 106586 213979 106589
rect 217182 106586 217242 106828
rect 307477 106800 307482 106856
rect 307538 106800 310040 106856
rect 307477 106798 310040 106800
rect 307477 106795 307543 106798
rect 251725 106586 251791 106589
rect 213913 106584 217242 106586
rect 213913 106528 213918 106584
rect 213974 106528 217242 106584
rect 213913 106526 217242 106528
rect 248952 106584 251791 106586
rect 248952 106528 251730 106584
rect 251786 106528 251791 106584
rect 248952 106526 251791 106528
rect 213913 106523 213979 106526
rect 251725 106523 251791 106526
rect 307661 106450 307727 106453
rect 307661 106448 310040 106450
rect 307661 106392 307666 106448
rect 307722 106392 310040 106448
rect 307661 106390 310040 106392
rect 307661 106387 307727 106390
rect 322933 106314 322999 106317
rect 321908 106312 322999 106314
rect 321908 106256 322938 106312
rect 322994 106256 322999 106312
rect 321908 106254 322999 106256
rect 322933 106251 322999 106254
rect 496905 106178 496971 106181
rect 494316 106176 496971 106178
rect 214005 105770 214071 105773
rect 217182 105770 217242 106148
rect 494316 106120 496910 106176
rect 496966 106120 496971 106176
rect 494316 106118 496971 106120
rect 496905 106115 496971 106118
rect 252461 106042 252527 106045
rect 248952 106040 252527 106042
rect 248952 105984 252466 106040
rect 252522 105984 252527 106040
rect 248952 105982 252527 105984
rect 252461 105979 252527 105982
rect 306925 105906 306991 105909
rect 416773 105906 416839 105909
rect 306925 105904 310040 105906
rect 306925 105848 306930 105904
rect 306986 105848 310040 105904
rect 306925 105846 310040 105848
rect 416773 105904 420164 105906
rect 416773 105848 416778 105904
rect 416834 105848 420164 105904
rect 416773 105846 420164 105848
rect 306925 105843 306991 105846
rect 416773 105843 416839 105846
rect 214005 105768 217242 105770
rect 214005 105712 214010 105768
rect 214066 105712 217242 105768
rect 214005 105710 217242 105712
rect 214005 105707 214071 105710
rect 252369 105634 252435 105637
rect 248952 105632 252435 105634
rect 214598 105164 214604 105228
rect 214668 105226 214674 105228
rect 217182 105226 217242 105604
rect 248952 105576 252374 105632
rect 252430 105576 252435 105632
rect 248952 105574 252435 105576
rect 252369 105571 252435 105574
rect 307477 105498 307543 105501
rect 307477 105496 310040 105498
rect 307477 105440 307482 105496
rect 307538 105440 310040 105496
rect 307477 105438 310040 105440
rect 307477 105435 307543 105438
rect 214668 105166 217242 105226
rect 214668 105164 214674 105166
rect 321878 105093 321938 105468
rect 213913 105090 213979 105093
rect 252277 105090 252343 105093
rect 213913 105088 217242 105090
rect 213913 105032 213918 105088
rect 213974 105032 217242 105088
rect 213913 105030 217242 105032
rect 248952 105088 252343 105090
rect 248952 105032 252282 105088
rect 252338 105032 252343 105088
rect 248952 105030 252343 105032
rect 213913 105027 213979 105030
rect 217182 104924 217242 105030
rect 252277 105027 252343 105030
rect 307661 105090 307727 105093
rect 307661 105088 310040 105090
rect 307661 105032 307666 105088
rect 307722 105032 310040 105088
rect 307661 105030 310040 105032
rect 321829 105088 321938 105093
rect 321829 105032 321834 105088
rect 321890 105032 321938 105088
rect 321829 105030 321938 105032
rect 307661 105027 307727 105030
rect 321829 105027 321895 105030
rect 494286 104821 494346 104924
rect 324405 104818 324471 104821
rect 321908 104816 324471 104818
rect 321908 104760 324410 104816
rect 324466 104760 324471 104816
rect 321908 104758 324471 104760
rect 324405 104755 324471 104758
rect 494237 104816 494346 104821
rect 494237 104760 494242 104816
rect 494298 104760 494346 104816
rect 494237 104758 494346 104760
rect 494237 104755 494303 104758
rect 252461 104682 252527 104685
rect 248952 104680 252527 104682
rect 248952 104624 252466 104680
rect 252522 104624 252527 104680
rect 248952 104622 252527 104624
rect 252461 104619 252527 104622
rect 306925 104682 306991 104685
rect 306925 104680 310040 104682
rect 306925 104624 306930 104680
rect 306986 104624 310040 104680
rect 306925 104622 310040 104624
rect 306925 104619 306991 104622
rect 307569 104274 307635 104277
rect 325601 104274 325667 104277
rect 307569 104272 310040 104274
rect 214414 103804 214420 103868
rect 214484 103866 214490 103868
rect 217182 103866 217242 104244
rect 307569 104216 307574 104272
rect 307630 104216 310040 104272
rect 307569 104214 310040 104216
rect 321878 104272 325667 104274
rect 321878 104216 325606 104272
rect 325662 104216 325667 104272
rect 321878 104214 325667 104216
rect 307569 104211 307635 104214
rect 252277 104138 252343 104141
rect 248952 104136 252343 104138
rect 248952 104080 252282 104136
rect 252338 104080 252343 104136
rect 248952 104078 252343 104080
rect 252277 104075 252343 104078
rect 321878 103972 321938 104214
rect 325601 104211 325667 104214
rect 416773 104138 416839 104141
rect 416773 104136 420164 104138
rect 416773 104080 416778 104136
rect 416834 104080 420164 104136
rect 416773 104078 420164 104080
rect 416773 104075 416839 104078
rect 214484 103806 217242 103866
rect 307661 103866 307727 103869
rect 495433 103866 495499 103869
rect 307661 103864 310040 103866
rect 307661 103808 307666 103864
rect 307722 103808 310040 103864
rect 307661 103806 310040 103808
rect 494316 103864 495499 103866
rect 494316 103808 495438 103864
rect 495494 103808 495499 103864
rect 494316 103806 495499 103808
rect 214484 103804 214490 103806
rect 307661 103803 307727 103806
rect 495433 103803 495499 103806
rect 213913 103730 213979 103733
rect 252369 103730 252435 103733
rect 213913 103728 217242 103730
rect 213913 103672 213918 103728
rect 213974 103672 217242 103728
rect 213913 103670 217242 103672
rect 248952 103728 252435 103730
rect 248952 103672 252374 103728
rect 252430 103672 252435 103728
rect 248952 103670 252435 103672
rect 213913 103667 213979 103670
rect 217182 103564 217242 103670
rect 252369 103667 252435 103670
rect 307569 103458 307635 103461
rect 307569 103456 310040 103458
rect 307569 103400 307574 103456
rect 307630 103400 310040 103456
rect 307569 103398 310040 103400
rect 307569 103395 307635 103398
rect 252461 103186 252527 103189
rect 248952 103184 252527 103186
rect 248952 103128 252466 103184
rect 252522 103128 252527 103184
rect 248952 103126 252527 103128
rect 252461 103123 252527 103126
rect 309504 102946 310132 103006
rect 213913 102506 213979 102509
rect 217182 102506 217242 102884
rect 305494 102852 305500 102916
rect 305564 102914 305570 102916
rect 309504 102914 309564 102946
rect 305564 102854 309564 102914
rect 305564 102852 305570 102854
rect 321694 102781 321754 103156
rect 252461 102778 252527 102781
rect 248952 102776 252527 102778
rect 248952 102720 252466 102776
rect 252522 102720 252527 102776
rect 248952 102718 252527 102720
rect 252461 102715 252527 102718
rect 321645 102776 321754 102781
rect 321645 102720 321650 102776
rect 321706 102720 321754 102776
rect 321645 102718 321754 102720
rect 321645 102715 321711 102718
rect 213913 102504 217242 102506
rect 213913 102448 213918 102504
rect 213974 102448 217242 102504
rect 213913 102446 217242 102448
rect 307661 102506 307727 102509
rect 416773 102506 416839 102509
rect 307661 102504 310040 102506
rect 307661 102448 307666 102504
rect 307722 102448 310040 102504
rect 416773 102504 420164 102506
rect 307661 102446 310040 102448
rect 213913 102443 213979 102446
rect 307661 102443 307727 102446
rect 65977 102370 66043 102373
rect 68142 102370 68816 102376
rect 65977 102368 68816 102370
rect 65977 102312 65982 102368
rect 66038 102316 68816 102368
rect 214833 102370 214899 102373
rect 214833 102368 217242 102370
rect 66038 102312 68202 102316
rect 65977 102310 68202 102312
rect 214833 102312 214838 102368
rect 214894 102312 217242 102368
rect 214833 102310 217242 102312
rect 65977 102307 66043 102310
rect 214833 102307 214899 102310
rect 217182 102204 217242 102310
rect 321694 102237 321754 102476
rect 416773 102448 416778 102504
rect 416834 102448 420164 102504
rect 416773 102446 420164 102448
rect 416773 102443 416839 102446
rect 252369 102234 252435 102237
rect 248952 102232 252435 102234
rect 248952 102176 252374 102232
rect 252430 102176 252435 102232
rect 248952 102174 252435 102176
rect 321694 102232 321803 102237
rect 493918 102236 493978 102748
rect 321694 102176 321742 102232
rect 321798 102176 321803 102232
rect 321694 102174 321803 102176
rect 252369 102171 252435 102174
rect 321737 102171 321803 102174
rect 493910 102172 493916 102236
rect 493980 102172 493986 102236
rect 307661 102098 307727 102101
rect 307661 102096 310040 102098
rect 307661 102040 307666 102096
rect 307722 102040 310040 102096
rect 307661 102038 310040 102040
rect 307661 102035 307727 102038
rect 251357 101826 251423 101829
rect 248952 101824 251423 101826
rect 248952 101768 251362 101824
rect 251418 101768 251423 101824
rect 248952 101766 251423 101768
rect 251357 101763 251423 101766
rect 307569 101690 307635 101693
rect 324313 101690 324379 101693
rect 497089 101690 497155 101693
rect 307569 101688 310040 101690
rect 307569 101632 307574 101688
rect 307630 101632 310040 101688
rect 307569 101630 310040 101632
rect 321908 101688 324379 101690
rect 321908 101632 324318 101688
rect 324374 101632 324379 101688
rect 321908 101630 324379 101632
rect 494316 101688 497155 101690
rect 494316 101632 497094 101688
rect 497150 101632 497155 101688
rect 494316 101630 497155 101632
rect 307569 101627 307635 101630
rect 324313 101627 324379 101630
rect 497089 101627 497155 101630
rect 214005 101282 214071 101285
rect 217182 101282 217242 101524
rect 252461 101418 252527 101421
rect 248952 101416 252527 101418
rect 248952 101360 252466 101416
rect 252522 101360 252527 101416
rect 248952 101358 252527 101360
rect 252461 101355 252527 101358
rect 214005 101280 217242 101282
rect 214005 101224 214010 101280
rect 214066 101224 217242 101280
rect 214005 101222 217242 101224
rect 306557 101282 306623 101285
rect 306557 101280 310040 101282
rect 306557 101224 306562 101280
rect 306618 101224 310040 101280
rect 306557 101222 310040 101224
rect 214005 101219 214071 101222
rect 306557 101219 306623 101222
rect 213913 101146 213979 101149
rect 213913 101144 217242 101146
rect 213913 101088 213918 101144
rect 213974 101088 217242 101144
rect 213913 101086 217242 101088
rect 213913 101083 213979 101086
rect 217182 100980 217242 101086
rect 251817 100874 251883 100877
rect 248952 100872 251883 100874
rect 248952 100816 251822 100872
rect 251878 100816 251883 100872
rect 248952 100814 251883 100816
rect 251817 100811 251883 100814
rect 306925 100874 306991 100877
rect 324497 100874 324563 100877
rect 306925 100872 310040 100874
rect 306925 100816 306930 100872
rect 306986 100816 310040 100872
rect 306925 100814 310040 100816
rect 321908 100872 324563 100874
rect 321908 100816 324502 100872
rect 324558 100816 324563 100872
rect 321908 100814 324563 100816
rect 306925 100811 306991 100814
rect 324497 100811 324563 100814
rect 416773 100874 416839 100877
rect 416773 100872 420164 100874
rect 416773 100816 416778 100872
rect 416834 100816 420164 100872
rect 416773 100814 420164 100816
rect 416773 100811 416839 100814
rect 66069 100738 66135 100741
rect 68142 100738 68816 100744
rect 66069 100736 68816 100738
rect 66069 100680 66074 100736
rect 66130 100684 68816 100736
rect 66130 100680 68202 100684
rect 66069 100678 68202 100680
rect 66069 100675 66135 100678
rect 493918 100469 493978 100572
rect 252461 100466 252527 100469
rect 248952 100464 252527 100466
rect 248952 100408 252466 100464
rect 252522 100408 252527 100464
rect 248952 100406 252527 100408
rect 252461 100403 252527 100406
rect 306557 100466 306623 100469
rect 306557 100464 310040 100466
rect 306557 100408 306562 100464
rect 306618 100408 310040 100464
rect 306557 100406 310040 100408
rect 493918 100464 494027 100469
rect 493918 100408 493966 100464
rect 494022 100408 494027 100464
rect 493918 100406 494027 100408
rect 306557 100403 306623 100406
rect 493961 100403 494027 100406
rect 166390 99996 166396 100060
rect 166460 100058 166466 100060
rect 214649 100058 214715 100061
rect 166460 100056 214715 100058
rect 166460 100000 214654 100056
rect 214710 100000 214715 100056
rect 166460 99998 214715 100000
rect 166460 99996 166466 99998
rect 214649 99995 214715 99998
rect 214005 99786 214071 99789
rect 217182 99786 217242 100300
rect 307569 100058 307635 100061
rect 307569 100056 310040 100058
rect 307569 100000 307574 100056
rect 307630 100000 310040 100056
rect 307569 99998 310040 100000
rect 307569 99995 307635 99998
rect 252369 99922 252435 99925
rect 248952 99920 252435 99922
rect 248952 99864 252374 99920
rect 252430 99864 252435 99920
rect 248952 99862 252435 99864
rect 252369 99859 252435 99862
rect 214005 99784 217242 99786
rect 214005 99728 214010 99784
rect 214066 99728 217242 99784
rect 214005 99726 217242 99728
rect 214005 99723 214071 99726
rect 321510 99653 321570 100164
rect 307661 99650 307727 99653
rect 307661 99648 310040 99650
rect 213913 99514 213979 99517
rect 213913 99512 216874 99514
rect 213913 99456 213918 99512
rect 213974 99456 216874 99512
rect 213913 99454 216874 99456
rect 213913 99451 213979 99454
rect 216814 99378 216874 99454
rect 217366 99378 217426 99620
rect 307661 99592 307666 99648
rect 307722 99592 310040 99648
rect 307661 99590 310040 99592
rect 321510 99648 321619 99653
rect 321510 99592 321558 99648
rect 321614 99592 321619 99648
rect 321510 99590 321619 99592
rect 307661 99587 307727 99590
rect 321553 99587 321619 99590
rect 252277 99514 252343 99517
rect 248952 99512 252343 99514
rect 248952 99456 252282 99512
rect 252338 99456 252343 99512
rect 248952 99454 252343 99456
rect 252277 99451 252343 99454
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 324313 99378 324379 99381
rect 216814 99318 217426 99378
rect 321908 99376 324379 99378
rect 321908 99320 324318 99376
rect 324374 99320 324379 99376
rect 321908 99318 324379 99320
rect 324313 99315 324379 99318
rect 360193 99378 360259 99381
rect 494278 99378 494284 99380
rect 360193 99376 494284 99378
rect 360193 99320 360198 99376
rect 360254 99320 494284 99376
rect 360193 99318 494284 99320
rect 360193 99315 360259 99318
rect 494278 99316 494284 99318
rect 494348 99316 494354 99380
rect 583520 99364 584960 99454
rect 307569 99106 307635 99109
rect 307569 99104 310040 99106
rect 307569 99048 307574 99104
rect 307630 99048 310040 99104
rect 307569 99046 310040 99048
rect 307569 99043 307635 99046
rect 252461 98970 252527 98973
rect 248952 98968 252527 98970
rect 214005 98426 214071 98429
rect 217182 98426 217242 98940
rect 248952 98912 252466 98968
rect 252522 98912 252527 98968
rect 248952 98910 252527 98912
rect 252461 98907 252527 98910
rect 306925 98698 306991 98701
rect 345013 98698 345079 98701
rect 360193 98698 360259 98701
rect 306925 98696 310040 98698
rect 306925 98640 306930 98696
rect 306986 98640 310040 98696
rect 306925 98638 310040 98640
rect 345013 98696 360259 98698
rect 345013 98640 345018 98696
rect 345074 98640 360198 98696
rect 360254 98640 360259 98696
rect 345013 98638 360259 98640
rect 306925 98635 306991 98638
rect 345013 98635 345079 98638
rect 360193 98635 360259 98638
rect 251909 98562 251975 98565
rect 324262 98562 324268 98564
rect 248952 98560 251975 98562
rect 248952 98504 251914 98560
rect 251970 98504 251975 98560
rect 248952 98502 251975 98504
rect 321908 98502 324268 98562
rect 251909 98499 251975 98502
rect 324262 98500 324268 98502
rect 324332 98500 324338 98564
rect 214005 98424 217242 98426
rect 214005 98368 214010 98424
rect 214066 98368 217242 98424
rect 214005 98366 217242 98368
rect 214005 98363 214071 98366
rect 307661 98290 307727 98293
rect 307661 98288 310040 98290
rect 213913 98018 213979 98021
rect 217366 98018 217426 98260
rect 307661 98232 307666 98288
rect 307722 98232 310040 98288
rect 307661 98230 310040 98232
rect 307661 98227 307727 98230
rect 252185 98018 252251 98021
rect 213913 98016 217426 98018
rect 213913 97960 213918 98016
rect 213974 97960 217426 98016
rect 213913 97958 217426 97960
rect 248952 98016 252251 98018
rect 248952 97960 252190 98016
rect 252246 97960 252251 98016
rect 248952 97958 252251 97960
rect 213913 97955 213979 97958
rect 252185 97955 252251 97958
rect 307477 97882 307543 97885
rect 324405 97882 324471 97885
rect 307477 97880 310040 97882
rect 307477 97824 307482 97880
rect 307538 97824 310040 97880
rect 307477 97822 310040 97824
rect 321908 97880 324471 97882
rect 321908 97824 324410 97880
rect 324466 97824 324471 97880
rect 321908 97822 324471 97824
rect 307477 97819 307543 97822
rect 324405 97819 324471 97822
rect -960 97610 480 97700
rect 2773 97610 2839 97613
rect 252461 97610 252527 97613
rect -960 97608 2839 97610
rect -960 97552 2778 97608
rect 2834 97552 2839 97608
rect 248952 97608 252527 97610
rect -960 97550 2839 97552
rect -960 97460 480 97550
rect 2773 97547 2839 97550
rect 214649 97066 214715 97069
rect 217182 97066 217242 97580
rect 248952 97552 252466 97608
rect 252522 97552 252527 97608
rect 248952 97550 252527 97552
rect 252461 97547 252527 97550
rect 309504 97370 310132 97430
rect 249190 97066 249196 97068
rect 214649 97064 217242 97066
rect 214649 97008 214654 97064
rect 214710 97008 217242 97064
rect 214649 97006 217242 97008
rect 248952 97006 249196 97066
rect 214649 97003 214715 97006
rect 249190 97004 249196 97006
rect 249260 97066 249266 97068
rect 251950 97066 251956 97068
rect 249260 97006 251956 97066
rect 249260 97004 249266 97006
rect 251950 97004 251956 97006
rect 252020 97004 252026 97068
rect 166206 96732 166212 96796
rect 166276 96794 166282 96796
rect 166276 96734 200130 96794
rect 166276 96732 166282 96734
rect 200070 96658 200130 96734
rect 217366 96658 217426 96900
rect 304206 96868 304212 96932
rect 304276 96930 304282 96932
rect 309504 96930 309564 97370
rect 324313 97066 324379 97069
rect 321908 97064 324379 97066
rect 304276 96870 309564 96930
rect 309734 96962 310132 97022
rect 321908 97008 324318 97064
rect 324374 97008 324379 97064
rect 321908 97006 324379 97008
rect 324313 97003 324379 97006
rect 304276 96868 304282 96870
rect 306966 96732 306972 96796
rect 307036 96794 307042 96796
rect 309734 96794 309794 96962
rect 307036 96734 309794 96794
rect 307036 96732 307042 96734
rect 252461 96658 252527 96661
rect 200070 96598 217426 96658
rect 248952 96656 252527 96658
rect 248952 96600 252466 96656
rect 252522 96600 252527 96656
rect 248952 96598 252527 96600
rect 252461 96595 252527 96598
rect 307661 96658 307727 96661
rect 307661 96656 310040 96658
rect 307661 96600 307666 96656
rect 307722 96600 310040 96656
rect 307661 96598 310040 96600
rect 307661 96595 307727 96598
rect 214741 95842 214807 95845
rect 217182 95842 217242 96356
rect 251173 96250 251239 96253
rect 248860 96248 251239 96250
rect 248860 96192 251178 96248
rect 251234 96192 251239 96248
rect 248860 96190 251239 96192
rect 251173 96187 251239 96190
rect 307661 96250 307727 96253
rect 307661 96248 310132 96250
rect 307661 96192 307666 96248
rect 307722 96192 310132 96248
rect 307661 96190 310132 96192
rect 307661 96187 307727 96190
rect 321510 95845 321570 96356
rect 335854 96324 335860 96388
rect 335924 96386 335930 96388
rect 343633 96386 343699 96389
rect 335924 96384 343699 96386
rect 335924 96328 343638 96384
rect 343694 96328 343699 96384
rect 335924 96326 343699 96328
rect 335924 96324 335930 96326
rect 343633 96323 343699 96326
rect 214741 95840 217242 95842
rect 214741 95784 214746 95840
rect 214802 95784 217242 95840
rect 214741 95782 217242 95784
rect 321461 95840 321570 95845
rect 321461 95784 321466 95840
rect 321522 95784 321570 95840
rect 321461 95782 321570 95784
rect 214741 95779 214807 95782
rect 321461 95779 321527 95782
rect 164877 95162 164943 95165
rect 166942 95162 166948 95164
rect 164877 95160 166948 95162
rect 164877 95104 164882 95160
rect 164938 95104 166948 95160
rect 164877 95102 166948 95104
rect 164877 95099 164943 95102
rect 166942 95100 166948 95102
rect 167012 95100 167018 95164
rect 381537 95162 381603 95165
rect 493910 95162 493916 95164
rect 381537 95160 493916 95162
rect 381537 95104 381542 95160
rect 381598 95104 493916 95160
rect 381537 95102 493916 95104
rect 381537 95099 381603 95102
rect 493910 95100 493916 95102
rect 493980 95100 493986 95164
rect 67449 94890 67515 94893
rect 214598 94890 214604 94892
rect 67449 94888 214604 94890
rect 67449 94832 67454 94888
rect 67510 94832 214604 94888
rect 67449 94830 214604 94832
rect 67449 94827 67515 94830
rect 214598 94828 214604 94830
rect 214668 94828 214674 94892
rect 85573 94756 85639 94757
rect 112345 94756 112411 94757
rect 125409 94756 125475 94757
rect 85528 94692 85534 94756
rect 85598 94754 85639 94756
rect 85598 94752 85690 94754
rect 85634 94696 85690 94752
rect 85598 94694 85690 94696
rect 85598 94692 85639 94694
rect 112320 94692 112326 94756
rect 112390 94754 112411 94756
rect 112390 94752 112482 94754
rect 112406 94696 112482 94752
rect 112390 94694 112482 94696
rect 112390 94692 112411 94694
rect 125376 94692 125382 94756
rect 125446 94754 125475 94756
rect 125446 94752 125538 94754
rect 125470 94696 125538 94752
rect 125446 94694 125538 94696
rect 125446 94692 125475 94694
rect 151302 94692 151308 94756
rect 151372 94754 151378 94756
rect 151624 94754 151630 94756
rect 151372 94694 151630 94754
rect 151372 94692 151378 94694
rect 151624 94692 151630 94694
rect 151694 94692 151700 94756
rect 85573 94691 85639 94692
rect 112345 94691 112411 94692
rect 125409 94691 125475 94692
rect 126646 93876 126652 93940
rect 126716 93938 126722 93940
rect 167637 93938 167703 93941
rect 126716 93936 167703 93938
rect 126716 93880 167642 93936
rect 167698 93880 167703 93936
rect 126716 93878 167703 93880
rect 126716 93876 126722 93878
rect 167637 93875 167703 93878
rect 57789 93802 57855 93805
rect 192569 93802 192635 93805
rect 57789 93800 192635 93802
rect 57789 93744 57794 93800
rect 57850 93744 192574 93800
rect 192630 93744 192635 93800
rect 57789 93742 192635 93744
rect 57789 93739 57855 93742
rect 192569 93739 192635 93742
rect 207657 93802 207723 93805
rect 324262 93802 324268 93804
rect 207657 93800 324268 93802
rect 207657 93744 207662 93800
rect 207718 93744 324268 93800
rect 207657 93742 324268 93744
rect 207657 93739 207723 93742
rect 324262 93740 324268 93742
rect 324332 93740 324338 93804
rect 118233 93668 118299 93669
rect 118182 93666 118188 93668
rect 118142 93606 118188 93666
rect 118252 93664 118299 93668
rect 169150 93666 169156 93668
rect 118294 93608 118299 93664
rect 118182 93604 118188 93606
rect 118252 93604 118299 93608
rect 118233 93603 118299 93604
rect 122790 93606 169156 93666
rect 98545 93532 98611 93533
rect 98494 93530 98500 93532
rect 98454 93470 98500 93530
rect 98564 93528 98611 93532
rect 98606 93472 98611 93528
rect 98494 93468 98500 93470
rect 98564 93468 98611 93472
rect 113214 93468 113220 93532
rect 113284 93530 113290 93532
rect 122790 93530 122850 93606
rect 169150 93604 169156 93606
rect 169220 93604 169226 93668
rect 129457 93532 129523 93533
rect 133137 93532 133203 93533
rect 151721 93532 151787 93533
rect 129406 93530 129412 93532
rect 113284 93470 122850 93530
rect 129366 93470 129412 93530
rect 129476 93528 129523 93532
rect 133086 93530 133092 93532
rect 129518 93472 129523 93528
rect 113284 93468 113290 93470
rect 129406 93468 129412 93470
rect 129476 93468 129523 93472
rect 133046 93470 133092 93530
rect 133156 93528 133203 93532
rect 151670 93530 151676 93532
rect 133198 93472 133203 93528
rect 133086 93468 133092 93470
rect 133156 93468 133203 93472
rect 151630 93470 151676 93530
rect 151740 93528 151787 93532
rect 151782 93472 151787 93528
rect 151670 93468 151676 93470
rect 151740 93468 151787 93472
rect 98545 93467 98611 93468
rect 129457 93467 129523 93468
rect 133137 93467 133203 93468
rect 151721 93467 151787 93468
rect 103329 93260 103395 93261
rect 110137 93260 110203 93261
rect 103278 93258 103284 93260
rect 103238 93198 103284 93258
rect 103348 93256 103395 93260
rect 110086 93258 110092 93260
rect 103390 93200 103395 93256
rect 103278 93196 103284 93198
rect 103348 93196 103395 93200
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 103329 93195 103395 93196
rect 110137 93195 110203 93196
rect 84326 92380 84332 92444
rect 84396 92442 84402 92444
rect 85113 92442 85179 92445
rect 86769 92444 86835 92445
rect 88977 92444 89043 92445
rect 107745 92444 107811 92445
rect 86718 92442 86724 92444
rect 84396 92440 85179 92442
rect 84396 92384 85118 92440
rect 85174 92384 85179 92440
rect 84396 92382 85179 92384
rect 86678 92382 86724 92442
rect 86788 92440 86835 92444
rect 88926 92442 88932 92444
rect 86830 92384 86835 92440
rect 84396 92380 84402 92382
rect 85113 92379 85179 92382
rect 86718 92380 86724 92382
rect 86788 92380 86835 92384
rect 88886 92382 88932 92442
rect 88996 92440 89043 92444
rect 107694 92442 107700 92444
rect 89038 92384 89043 92440
rect 88926 92380 88932 92382
rect 88996 92380 89043 92384
rect 107654 92382 107700 92442
rect 107764 92440 107811 92444
rect 107806 92384 107811 92440
rect 107694 92380 107700 92382
rect 107764 92380 107811 92384
rect 86769 92379 86835 92380
rect 88977 92379 89043 92380
rect 107745 92379 107811 92380
rect 114369 92442 114435 92445
rect 115473 92444 115539 92445
rect 114502 92442 114508 92444
rect 114369 92440 114508 92442
rect 114369 92384 114374 92440
rect 114430 92384 114508 92440
rect 114369 92382 114508 92384
rect 114369 92379 114435 92382
rect 114502 92380 114508 92382
rect 114572 92380 114578 92444
rect 115422 92442 115428 92444
rect 115382 92382 115428 92442
rect 115492 92440 115539 92444
rect 115534 92384 115539 92440
rect 115422 92380 115428 92382
rect 115492 92380 115539 92384
rect 120206 92380 120212 92444
rect 120276 92442 120282 92444
rect 120349 92442 120415 92445
rect 120276 92440 120415 92442
rect 120276 92384 120354 92440
rect 120410 92384 120415 92440
rect 120276 92382 120415 92384
rect 120276 92380 120282 92382
rect 115473 92379 115539 92380
rect 120349 92379 120415 92382
rect 121678 92380 121684 92444
rect 121748 92442 121754 92444
rect 122097 92442 122163 92445
rect 130745 92444 130811 92445
rect 130694 92442 130700 92444
rect 121748 92440 122163 92442
rect 121748 92384 122102 92440
rect 122158 92384 122163 92440
rect 121748 92382 122163 92384
rect 130654 92382 130700 92442
rect 130764 92440 130811 92444
rect 130806 92384 130811 92440
rect 121748 92380 121754 92382
rect 122097 92379 122163 92382
rect 130694 92380 130700 92382
rect 130764 92380 130811 92384
rect 134374 92380 134380 92444
rect 134444 92442 134450 92444
rect 135161 92442 135227 92445
rect 136081 92444 136147 92445
rect 136030 92442 136036 92444
rect 134444 92440 135227 92442
rect 134444 92384 135166 92440
rect 135222 92384 135227 92440
rect 134444 92382 135227 92384
rect 135990 92382 136036 92442
rect 136100 92440 136147 92444
rect 136142 92384 136147 92440
rect 134444 92380 134450 92382
rect 130745 92379 130811 92380
rect 135161 92379 135227 92382
rect 136030 92380 136036 92382
rect 136100 92380 136147 92384
rect 151486 92380 151492 92444
rect 151556 92442 151562 92444
rect 151629 92442 151695 92445
rect 151556 92440 151695 92442
rect 151556 92384 151634 92440
rect 151690 92384 151695 92440
rect 151556 92382 151695 92384
rect 151556 92380 151562 92382
rect 136081 92379 136147 92380
rect 151629 92379 151695 92382
rect 117998 92244 118004 92308
rect 118068 92306 118074 92308
rect 166390 92306 166396 92308
rect 118068 92246 166396 92306
rect 118068 92244 118074 92246
rect 166390 92244 166396 92246
rect 166460 92244 166466 92308
rect 90214 91700 90220 91764
rect 90284 91762 90290 91764
rect 90541 91762 90607 91765
rect 90284 91760 90607 91762
rect 90284 91704 90546 91760
rect 90602 91704 90607 91760
rect 90284 91702 90607 91704
rect 90284 91700 90290 91702
rect 90541 91699 90607 91702
rect 93894 91700 93900 91764
rect 93964 91762 93970 91764
rect 95049 91762 95115 91765
rect 126513 91764 126579 91765
rect 126462 91762 126468 91764
rect 93964 91760 95115 91762
rect 93964 91704 95054 91760
rect 95110 91704 95115 91760
rect 93964 91702 95115 91704
rect 126422 91702 126468 91762
rect 126532 91760 126579 91764
rect 126574 91704 126579 91760
rect 93964 91700 93970 91702
rect 95049 91699 95115 91702
rect 126462 91700 126468 91702
rect 126532 91700 126579 91704
rect 126513 91699 126579 91700
rect 110638 91564 110644 91628
rect 110708 91626 110714 91628
rect 198273 91626 198339 91629
rect 110708 91624 198339 91626
rect 110708 91568 198278 91624
rect 198334 91568 198339 91624
rect 110708 91566 198339 91568
rect 110708 91564 110714 91566
rect 198273 91563 198339 91566
rect 101857 91492 101923 91493
rect 122833 91492 122899 91493
rect 101806 91490 101812 91492
rect 101766 91430 101812 91490
rect 101876 91488 101923 91492
rect 101918 91432 101923 91488
rect 101806 91428 101812 91430
rect 101876 91428 101923 91432
rect 122782 91428 122788 91492
rect 122852 91490 122899 91492
rect 122852 91488 122944 91490
rect 122894 91432 122944 91488
rect 122852 91430 122944 91432
rect 122852 91428 122899 91430
rect 152038 91428 152044 91492
rect 152108 91490 152114 91492
rect 153009 91490 153075 91493
rect 152108 91488 153075 91490
rect 152108 91432 153014 91488
rect 153070 91432 153075 91488
rect 152108 91430 153075 91432
rect 152108 91428 152114 91430
rect 101857 91427 101923 91428
rect 122833 91427 122899 91428
rect 153009 91427 153075 91430
rect 96654 91292 96660 91356
rect 96724 91354 96730 91356
rect 97901 91354 97967 91357
rect 96724 91352 97967 91354
rect 96724 91296 97906 91352
rect 97962 91296 97967 91352
rect 96724 91294 97967 91296
rect 96724 91292 96730 91294
rect 97901 91291 97967 91294
rect 98126 91292 98132 91356
rect 98196 91354 98202 91356
rect 99189 91354 99255 91357
rect 98196 91352 99255 91354
rect 98196 91296 99194 91352
rect 99250 91296 99255 91352
rect 98196 91294 99255 91296
rect 98196 91292 98202 91294
rect 99189 91291 99255 91294
rect 100886 91292 100892 91356
rect 100956 91354 100962 91356
rect 102041 91354 102107 91357
rect 100956 91352 102107 91354
rect 100956 91296 102046 91352
rect 102102 91296 102107 91352
rect 100956 91294 102107 91296
rect 100956 91292 100962 91294
rect 102041 91291 102107 91294
rect 106774 91292 106780 91356
rect 106844 91354 106850 91356
rect 107285 91354 107351 91357
rect 106844 91352 107351 91354
rect 106844 91296 107290 91352
rect 107346 91296 107351 91352
rect 106844 91294 107351 91296
rect 106844 91292 106850 91294
rect 107285 91291 107351 91294
rect 109166 91292 109172 91356
rect 109236 91354 109242 91356
rect 110229 91354 110295 91357
rect 109236 91352 110295 91354
rect 109236 91296 110234 91352
rect 110290 91296 110295 91352
rect 109236 91294 110295 91296
rect 109236 91292 109242 91294
rect 110229 91291 110295 91294
rect 116710 91292 116716 91356
rect 116780 91354 116786 91356
rect 117129 91354 117195 91357
rect 116780 91352 117195 91354
rect 116780 91296 117134 91352
rect 117190 91296 117195 91352
rect 116780 91294 117195 91296
rect 116780 91292 116786 91294
rect 117129 91291 117195 91294
rect 119286 91292 119292 91356
rect 119356 91354 119362 91356
rect 119889 91354 119955 91357
rect 119356 91352 119955 91354
rect 119356 91296 119894 91352
rect 119950 91296 119955 91352
rect 119356 91294 119955 91296
rect 119356 91292 119362 91294
rect 119889 91291 119955 91294
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75361 91218 75427 91221
rect 88057 91220 88123 91221
rect 88006 91218 88012 91220
rect 74828 91216 75427 91218
rect 74828 91160 75366 91216
rect 75422 91160 75427 91216
rect 74828 91158 75427 91160
rect 87966 91158 88012 91218
rect 88076 91216 88123 91220
rect 88118 91160 88123 91216
rect 74828 91156 74834 91158
rect 75361 91155 75427 91158
rect 88006 91156 88012 91158
rect 88076 91156 88123 91160
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 92381 91218 92447 91221
rect 91388 91216 92447 91218
rect 91388 91160 92386 91216
rect 92442 91160 92447 91216
rect 91388 91158 92447 91160
rect 91388 91156 91394 91158
rect 88057 91155 88123 91156
rect 92381 91155 92447 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93761 91218 93827 91221
rect 92676 91216 93827 91218
rect 92676 91160 93766 91216
rect 93822 91160 93827 91216
rect 92676 91158 93827 91160
rect 92676 91156 92682 91158
rect 93761 91155 93827 91158
rect 94998 91156 95004 91220
rect 95068 91218 95074 91220
rect 95141 91218 95207 91221
rect 95068 91216 95207 91218
rect 95068 91160 95146 91216
rect 95202 91160 95207 91216
rect 95068 91158 95207 91160
rect 95068 91156 95074 91158
rect 95141 91155 95207 91158
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 96521 91155 96587 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97809 91218 97875 91221
rect 97276 91216 97875 91218
rect 97276 91160 97814 91216
rect 97870 91160 97875 91216
rect 97276 91158 97875 91160
rect 97276 91156 97282 91158
rect 97809 91155 97875 91158
rect 99046 91156 99052 91220
rect 99116 91218 99122 91220
rect 99281 91218 99347 91221
rect 99116 91216 99347 91218
rect 99116 91160 99286 91216
rect 99342 91160 99347 91216
rect 99116 91158 99347 91160
rect 99116 91156 99122 91158
rect 99281 91155 99347 91158
rect 99966 91156 99972 91220
rect 100036 91218 100042 91220
rect 100201 91218 100267 91221
rect 100569 91220 100635 91221
rect 100518 91218 100524 91220
rect 100036 91216 100267 91218
rect 100036 91160 100206 91216
rect 100262 91160 100267 91216
rect 100036 91158 100267 91160
rect 100478 91158 100524 91218
rect 100588 91216 100635 91220
rect 101949 91220 102015 91221
rect 101949 91218 101996 91220
rect 100630 91160 100635 91216
rect 100036 91156 100042 91158
rect 100201 91155 100267 91158
rect 100518 91156 100524 91158
rect 100588 91156 100635 91160
rect 101904 91216 101996 91218
rect 101904 91160 101954 91216
rect 101904 91158 101996 91160
rect 100569 91155 100635 91156
rect 101949 91156 101996 91158
rect 102060 91156 102066 91220
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 103421 91218 103487 91221
rect 102796 91216 103487 91218
rect 102796 91160 103426 91216
rect 103482 91160 103487 91216
rect 102796 91158 103487 91160
rect 102796 91156 102802 91158
rect 101949 91155 102015 91156
rect 103421 91155 103487 91158
rect 104198 91156 104204 91220
rect 104268 91218 104274 91220
rect 104433 91218 104499 91221
rect 104268 91216 104499 91218
rect 104268 91160 104438 91216
rect 104494 91160 104499 91216
rect 104268 91158 104499 91160
rect 104268 91156 104274 91158
rect 104433 91155 104499 91158
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104801 91218 104867 91221
rect 105537 91220 105603 91221
rect 105486 91218 105492 91220
rect 104636 91216 104867 91218
rect 104636 91160 104806 91216
rect 104862 91160 104867 91216
rect 104636 91158 104867 91160
rect 105446 91158 105492 91218
rect 105556 91216 105603 91220
rect 105598 91160 105603 91216
rect 104636 91156 104642 91158
rect 104801 91155 104867 91158
rect 105486 91156 105492 91158
rect 105556 91156 105603 91160
rect 105670 91156 105676 91220
rect 105740 91218 105746 91220
rect 106089 91218 106155 91221
rect 105740 91216 106155 91218
rect 105740 91160 106094 91216
rect 106150 91160 106155 91216
rect 105740 91158 106155 91160
rect 105740 91156 105746 91158
rect 105537 91155 105603 91156
rect 106089 91155 106155 91158
rect 106406 91156 106412 91220
rect 106476 91218 106482 91220
rect 107561 91218 107627 91221
rect 106476 91216 107627 91218
rect 106476 91160 107566 91216
rect 107622 91160 107627 91216
rect 106476 91158 107627 91160
rect 106476 91156 106482 91158
rect 107561 91155 107627 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108941 91218 109007 91221
rect 108132 91216 109007 91218
rect 108132 91160 108946 91216
rect 109002 91160 109007 91216
rect 108132 91158 109007 91160
rect 108132 91156 108138 91158
rect 108941 91155 109007 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110321 91218 110387 91221
rect 111241 91220 111307 91221
rect 111190 91218 111196 91220
rect 109604 91216 110387 91218
rect 109604 91160 110326 91216
rect 110382 91160 110387 91216
rect 109604 91158 110387 91160
rect 111150 91158 111196 91218
rect 111260 91216 111307 91220
rect 111302 91160 111307 91216
rect 109604 91156 109610 91158
rect 110321 91155 110387 91158
rect 111190 91156 111196 91158
rect 111260 91156 111307 91160
rect 111926 91156 111932 91220
rect 111996 91218 112002 91220
rect 112437 91218 112503 91221
rect 111996 91216 112503 91218
rect 111996 91160 112442 91216
rect 112498 91160 112503 91216
rect 111996 91158 112503 91160
rect 111996 91156 112002 91158
rect 111241 91155 111307 91156
rect 112437 91155 112503 91158
rect 114318 91156 114324 91220
rect 114388 91218 114394 91220
rect 114461 91218 114527 91221
rect 114921 91220 114987 91221
rect 115841 91220 115907 91221
rect 114870 91218 114876 91220
rect 114388 91216 114527 91218
rect 114388 91160 114466 91216
rect 114522 91160 114527 91216
rect 114388 91158 114527 91160
rect 114830 91158 114876 91218
rect 114940 91216 114987 91220
rect 115790 91218 115796 91220
rect 114982 91160 114987 91216
rect 114388 91156 114394 91158
rect 114461 91155 114527 91158
rect 114870 91156 114876 91158
rect 114940 91156 114987 91160
rect 115750 91158 115796 91218
rect 115860 91216 115907 91220
rect 115902 91160 115907 91216
rect 115790 91156 115796 91158
rect 115860 91156 115907 91160
rect 117078 91156 117084 91220
rect 117148 91218 117154 91220
rect 117221 91218 117287 91221
rect 117148 91216 117287 91218
rect 117148 91160 117226 91216
rect 117282 91160 117287 91216
rect 117148 91158 117287 91160
rect 117148 91156 117154 91158
rect 114921 91155 114987 91156
rect 115841 91155 115907 91156
rect 117221 91155 117287 91158
rect 119654 91156 119660 91220
rect 119724 91218 119730 91220
rect 119981 91218 120047 91221
rect 120625 91220 120691 91221
rect 120574 91218 120580 91220
rect 119724 91216 120047 91218
rect 119724 91160 119986 91216
rect 120042 91160 120047 91216
rect 119724 91158 120047 91160
rect 120534 91158 120580 91218
rect 120644 91216 120691 91220
rect 120686 91160 120691 91216
rect 119724 91156 119730 91158
rect 119981 91155 120047 91158
rect 120574 91156 120580 91158
rect 120644 91156 120691 91160
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122741 91218 122807 91221
rect 122116 91216 122807 91218
rect 122116 91160 122746 91216
rect 122802 91160 122807 91216
rect 122116 91158 122807 91160
rect 122116 91156 122122 91158
rect 120625 91155 120691 91156
rect 122741 91155 122807 91158
rect 123150 91156 123156 91220
rect 123220 91218 123226 91220
rect 123293 91218 123359 91221
rect 123220 91216 123359 91218
rect 123220 91160 123298 91216
rect 123354 91160 123359 91216
rect 123220 91158 123359 91160
rect 123220 91156 123226 91158
rect 123293 91155 123359 91158
rect 123937 91218 124003 91221
rect 124070 91218 124076 91220
rect 123937 91216 124076 91218
rect 123937 91160 123942 91216
rect 123998 91160 124076 91216
rect 123937 91158 124076 91160
rect 123937 91155 124003 91158
rect 124070 91156 124076 91158
rect 124140 91156 124146 91220
rect 124438 91156 124444 91220
rect 124508 91218 124514 91220
rect 124765 91218 124831 91221
rect 124508 91216 124831 91218
rect 124508 91160 124770 91216
rect 124826 91160 124831 91216
rect 124508 91158 124831 91160
rect 124508 91156 124514 91158
rect 124765 91155 124831 91158
rect 125726 91156 125732 91220
rect 125796 91218 125802 91220
rect 126881 91218 126947 91221
rect 127617 91220 127683 91221
rect 132401 91220 132467 91221
rect 127566 91218 127572 91220
rect 125796 91216 126947 91218
rect 125796 91160 126886 91216
rect 126942 91160 126947 91216
rect 125796 91158 126947 91160
rect 127526 91158 127572 91218
rect 127636 91216 127683 91220
rect 132350 91218 132356 91220
rect 127678 91160 127683 91216
rect 125796 91156 125802 91158
rect 126881 91155 126947 91158
rect 127566 91156 127572 91158
rect 127636 91156 127683 91160
rect 132310 91158 132356 91218
rect 132420 91216 132467 91220
rect 132462 91160 132467 91216
rect 132350 91156 132356 91158
rect 132420 91156 132467 91160
rect 151302 91156 151308 91220
rect 151372 91218 151378 91220
rect 151445 91218 151511 91221
rect 151372 91216 151511 91218
rect 151372 91160 151450 91216
rect 151506 91160 151511 91216
rect 151372 91158 151511 91160
rect 151372 91156 151378 91158
rect 127617 91155 127683 91156
rect 132401 91155 132467 91156
rect 151445 91155 151511 91158
rect 67633 91082 67699 91085
rect 214414 91082 214420 91084
rect 67633 91080 214420 91082
rect 67633 91024 67638 91080
rect 67694 91024 214420 91080
rect 67633 91022 214420 91024
rect 67633 91019 67699 91022
rect 214414 91020 214420 91022
rect 214484 91020 214490 91084
rect 66069 88226 66135 88229
rect 166206 88226 166212 88228
rect 66069 88224 166212 88226
rect 66069 88168 66074 88224
rect 66130 88168 166212 88224
rect 66069 88166 166212 88168
rect 66069 88163 66135 88166
rect 166206 88164 166212 88166
rect 166276 88164 166282 88228
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 112437 85506 112503 85509
rect 170254 85506 170260 85508
rect 112437 85504 170260 85506
rect 112437 85448 112442 85504
rect 112498 85448 170260 85504
rect 112437 85446 170260 85448
rect 112437 85443 112503 85446
rect 170254 85444 170260 85446
rect 170324 85444 170330 85508
rect -960 84690 480 84780
rect 173014 84764 173020 84828
rect 173084 84826 173090 84828
rect 261477 84826 261543 84829
rect 173084 84824 261543 84826
rect 173084 84768 261482 84824
rect 261538 84768 261543 84824
rect 173084 84766 261543 84768
rect 173084 84764 173090 84766
rect 261477 84763 261543 84766
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 187049 82242 187115 82245
rect 251357 82242 251423 82245
rect 334566 82242 334572 82244
rect 187049 82240 334572 82242
rect 187049 82184 187054 82240
rect 187110 82184 251362 82240
rect 251418 82184 334572 82240
rect 187049 82182 334572 82184
rect 187049 82179 187115 82182
rect 251357 82179 251423 82182
rect 334566 82180 334572 82182
rect 334636 82180 334642 82244
rect 188521 82106 188587 82109
rect 307150 82106 307156 82108
rect 188521 82104 307156 82106
rect 188521 82048 188526 82104
rect 188582 82048 307156 82104
rect 188521 82046 307156 82048
rect 188521 82043 188587 82046
rect 307150 82044 307156 82046
rect 307220 82044 307226 82108
rect 104801 81426 104867 81429
rect 170438 81426 170444 81428
rect 104801 81424 170444 81426
rect 104801 81368 104806 81424
rect 104862 81368 170444 81424
rect 104801 81366 170444 81368
rect 104801 81363 104867 81366
rect 170438 81364 170444 81366
rect 170508 81364 170514 81428
rect 191230 81364 191236 81428
rect 191300 81426 191306 81428
rect 316033 81426 316099 81429
rect 191300 81424 316099 81426
rect 191300 81368 316038 81424
rect 316094 81368 316099 81424
rect 191300 81366 316099 81368
rect 191300 81364 191306 81366
rect 316033 81363 316099 81366
rect 345054 81364 345060 81428
rect 345124 81426 345130 81428
rect 345749 81426 345815 81429
rect 345124 81424 345815 81426
rect 345124 81368 345754 81424
rect 345810 81368 345815 81424
rect 345124 81366 345815 81368
rect 345124 81364 345130 81366
rect 345749 81363 345815 81366
rect 177246 79324 177252 79388
rect 177316 79386 177322 79388
rect 260189 79386 260255 79389
rect 177316 79384 260255 79386
rect 177316 79328 260194 79384
rect 260250 79328 260255 79384
rect 177316 79326 260255 79328
rect 177316 79324 177322 79326
rect 260189 79323 260255 79326
rect 99281 78570 99347 78573
rect 168966 78570 168972 78572
rect 99281 78568 168972 78570
rect 99281 78512 99286 78568
rect 99342 78512 168972 78568
rect 99281 78510 168972 78512
rect 99281 78507 99347 78510
rect 168966 78508 168972 78510
rect 169036 78508 169042 78572
rect 304758 77828 304764 77892
rect 304828 77890 304834 77892
rect 338246 77890 338252 77892
rect 304828 77830 338252 77890
rect 304828 77828 304834 77830
rect 338246 77828 338252 77830
rect 338316 77890 338322 77892
rect 339125 77890 339191 77893
rect 338316 77888 339191 77890
rect 338316 77832 339130 77888
rect 339186 77832 339191 77888
rect 338316 77830 339191 77832
rect 338316 77828 338322 77830
rect 339125 77827 339191 77830
rect 273846 76604 273852 76668
rect 273916 76666 273922 76668
rect 276013 76666 276079 76669
rect 334801 76666 334867 76669
rect 273916 76664 334867 76666
rect 273916 76608 276018 76664
rect 276074 76608 334806 76664
rect 334862 76608 334867 76664
rect 273916 76606 334867 76608
rect 273916 76604 273922 76606
rect 276013 76603 276079 76606
rect 334801 76603 334867 76606
rect 11053 76530 11119 76533
rect 304206 76530 304212 76532
rect 11053 76528 304212 76530
rect 11053 76472 11058 76528
rect 11114 76472 304212 76528
rect 11053 76470 304212 76472
rect 11053 76467 11119 76470
rect 304206 76468 304212 76470
rect 304276 76468 304282 76532
rect 66662 75108 66668 75172
rect 66732 75170 66738 75172
rect 289077 75170 289143 75173
rect 66732 75168 289143 75170
rect 66732 75112 289082 75168
rect 289138 75112 289143 75168
rect 66732 75110 289143 75112
rect 66732 75108 66738 75110
rect 289077 75107 289143 75110
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 60590 62732 60596 62796
rect 60660 62794 60666 62796
rect 280797 62794 280863 62797
rect 60660 62792 280863 62794
rect 60660 62736 280802 62792
rect 280858 62736 280863 62792
rect 60660 62734 280863 62736
rect 60660 62732 60666 62734
rect 280797 62731 280863 62734
rect 260189 62114 260255 62117
rect 336038 62114 336044 62116
rect 260189 62112 336044 62114
rect 260189 62056 260194 62112
rect 260250 62056 336044 62112
rect 260189 62054 336044 62056
rect 260189 62051 260255 62054
rect 336038 62052 336044 62054
rect 336108 62052 336114 62116
rect 45553 61570 45619 61573
rect 260046 61570 260052 61572
rect 45553 61568 260052 61570
rect 45553 61512 45558 61568
rect 45614 61512 260052 61568
rect 45553 61510 260052 61512
rect 45553 61507 45619 61510
rect 260046 61508 260052 61510
rect 260116 61508 260122 61572
rect 271086 61508 271092 61572
rect 271156 61570 271162 61572
rect 271873 61570 271939 61573
rect 273161 61570 273227 61573
rect 271156 61568 273227 61570
rect 271156 61512 271878 61568
rect 271934 61512 273166 61568
rect 273222 61512 273227 61568
rect 271156 61510 273227 61512
rect 271156 61508 271162 61510
rect 271873 61507 271939 61510
rect 273161 61507 273227 61510
rect 61878 61372 61884 61436
rect 61948 61434 61954 61436
rect 285213 61434 285279 61437
rect 61948 61432 285279 61434
rect 61948 61376 285218 61432
rect 285274 61376 285279 61432
rect 61948 61374 285279 61376
rect 61948 61372 61954 61374
rect 285213 61371 285279 61374
rect 259453 60754 259519 60757
rect 260189 60754 260255 60757
rect 259453 60752 260255 60754
rect 259453 60696 259458 60752
rect 259514 60696 260194 60752
rect 260250 60696 260255 60752
rect 259453 60694 260255 60696
rect 259453 60691 259519 60694
rect 260189 60691 260255 60694
rect 59118 59876 59124 59940
rect 59188 59938 59194 59940
rect 332593 59938 332659 59941
rect 59188 59936 332659 59938
rect 59188 59880 332598 59936
rect 332654 59880 332659 59936
rect 59188 59878 332659 59880
rect 59188 59876 59194 59878
rect 332593 59875 332659 59878
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 59353 57218 59419 57221
rect 302734 57218 302740 57220
rect 59353 57216 302740 57218
rect 59353 57160 59358 57216
rect 59414 57160 302740 57216
rect 59353 57158 302740 57160
rect 59353 57155 59419 57158
rect 302734 57156 302740 57158
rect 302804 57156 302810 57220
rect 79317 51778 79383 51781
rect 306966 51778 306972 51780
rect 79317 51776 306972 51778
rect 79317 51720 79322 51776
rect 79378 51720 306972 51776
rect 79317 51718 306972 51720
rect 79317 51715 79383 51718
rect 306966 51716 306972 51718
rect 307036 51716 307042 51780
rect 340873 47564 340939 47565
rect 340822 47500 340828 47564
rect 340892 47562 340939 47564
rect 340892 47560 340984 47562
rect 340934 47504 340984 47560
rect 340892 47502 340984 47504
rect 340892 47500 340939 47502
rect 340873 47499 340939 47500
rect 284293 46882 284359 46885
rect 285213 46882 285279 46885
rect 338614 46882 338620 46884
rect 284293 46880 338620 46882
rect 284293 46824 284298 46880
rect 284354 46824 285218 46880
rect 285274 46824 338620 46880
rect 284293 46822 338620 46824
rect 284293 46819 284359 46822
rect 285213 46819 285279 46822
rect 338614 46820 338620 46822
rect 338684 46820 338690 46884
rect 347773 46882 347839 46885
rect 348417 46882 348483 46885
rect 496854 46882 496860 46884
rect 347773 46880 496860 46882
rect 347773 46824 347778 46880
rect 347834 46824 348422 46880
rect 348478 46824 496860 46880
rect 347773 46822 496860 46824
rect 347773 46819 347839 46822
rect 348417 46819 348483 46822
rect 496854 46820 496860 46822
rect 496924 46820 496930 46884
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 268326 44780 268332 44844
rect 268396 44842 268402 44844
rect 333973 44842 334039 44845
rect 495934 44842 495940 44844
rect 268396 44840 495940 44842
rect 268396 44784 333978 44840
rect 334034 44784 495940 44840
rect 268396 44782 495940 44784
rect 268396 44780 268402 44782
rect 333973 44779 334039 44782
rect 495934 44780 495940 44782
rect 496004 44780 496010 44844
rect 186814 43420 186820 43484
rect 186884 43482 186890 43484
rect 316125 43482 316191 43485
rect 317321 43482 317387 43485
rect 186884 43480 317387 43482
rect 186884 43424 316130 43480
rect 316186 43424 317326 43480
rect 317382 43424 317387 43480
rect 186884 43422 317387 43424
rect 186884 43420 186890 43422
rect 316125 43419 316191 43422
rect 317321 43419 317387 43422
rect 342345 41308 342411 41309
rect 342294 41306 342300 41308
rect 342254 41246 342300 41306
rect 342364 41304 342411 41308
rect 342406 41248 342411 41304
rect 342294 41244 342300 41246
rect 342364 41244 342411 41248
rect 342345 41243 342411 41244
rect 184054 40564 184060 40628
rect 184124 40626 184130 40628
rect 308489 40626 308555 40629
rect 184124 40624 308555 40626
rect 184124 40568 308494 40624
rect 308550 40568 308555 40624
rect 184124 40566 308555 40568
rect 184124 40564 184130 40566
rect 308489 40563 308555 40566
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 191046 29548 191052 29612
rect 191116 29610 191122 29612
rect 276657 29610 276723 29613
rect 278037 29610 278103 29613
rect 191116 29608 278103 29610
rect 191116 29552 276662 29608
rect 276718 29552 278042 29608
rect 278098 29552 278103 29608
rect 191116 29550 278103 29552
rect 191116 29548 191122 29550
rect 276657 29547 276723 29550
rect 278037 29547 278103 29550
rect 81433 26890 81499 26893
rect 250294 26890 250300 26892
rect 81433 26888 250300 26890
rect 81433 26832 81438 26888
rect 81494 26832 250300 26888
rect 81433 26830 250300 26832
rect 81433 26827 81499 26830
rect 250294 26828 250300 26830
rect 250364 26828 250370 26892
rect 192334 26148 192340 26212
rect 192404 26210 192410 26212
rect 330477 26210 330543 26213
rect 192404 26208 330543 26210
rect 192404 26152 330482 26208
rect 330538 26152 330543 26208
rect 192404 26150 330543 26152
rect 192404 26148 192410 26150
rect 330477 26147 330543 26150
rect 106273 25530 106339 25533
rect 253054 25530 253060 25532
rect 106273 25528 253060 25530
rect 106273 25472 106278 25528
rect 106334 25472 253060 25528
rect 106273 25470 253060 25472
rect 106273 25467 106339 25470
rect 253054 25468 253060 25470
rect 253124 25468 253130 25532
rect 329833 24986 329899 24989
rect 330477 24986 330543 24989
rect 329833 24984 330543 24986
rect 329833 24928 329838 24984
rect 329894 24928 330482 24984
rect 330538 24928 330543 24984
rect 329833 24926 330543 24928
rect 329833 24923 329899 24926
rect 330477 24923 330543 24926
rect 188286 20572 188292 20636
rect 188356 20634 188362 20636
rect 267733 20634 267799 20637
rect 268469 20634 268535 20637
rect 188356 20632 268535 20634
rect 188356 20576 267738 20632
rect 267794 20576 268474 20632
rect 268530 20576 268535 20632
rect 188356 20574 268535 20576
rect 188356 20572 188362 20574
rect 267733 20571 267799 20574
rect 268469 20571 268535 20574
rect 66110 19892 66116 19956
rect 66180 19954 66186 19956
rect 249241 19954 249307 19957
rect 66180 19952 249307 19954
rect 66180 19896 249246 19952
rect 249302 19896 249307 19952
rect 66180 19894 249307 19896
rect 66180 19892 66186 19894
rect 249241 19891 249307 19894
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 8201 16554 8267 16557
rect 248454 16554 248460 16556
rect 8201 16552 248460 16554
rect 8201 16496 8206 16552
rect 8262 16496 248460 16552
rect 8201 16494 248460 16496
rect 8201 16491 8267 16494
rect 248454 16492 248460 16494
rect 248524 16492 248530 16556
rect 44265 13018 44331 13021
rect 305494 13018 305500 13020
rect 44265 13016 305500 13018
rect 44265 12960 44270 13016
rect 44326 12960 305500 13016
rect 44265 12958 305500 12960
rect 44265 12955 44331 12958
rect 305494 12956 305500 12958
rect 305564 12956 305570 13020
rect 340822 11732 340828 11796
rect 340892 11794 340898 11796
rect 342161 11794 342227 11797
rect 340892 11792 342227 11794
rect 340892 11736 342166 11792
rect 342222 11736 342227 11792
rect 340892 11734 342227 11736
rect 340892 11732 340898 11734
rect 342161 11731 342227 11734
rect 62982 10916 62988 10980
rect 63052 10978 63058 10980
rect 242893 10978 242959 10981
rect 243537 10978 243603 10981
rect 63052 10976 243603 10978
rect 63052 10920 242898 10976
rect 242954 10920 243542 10976
rect 243598 10920 243603 10976
rect 63052 10918 243603 10920
rect 63052 10916 63058 10918
rect 242893 10915 242959 10918
rect 243537 10915 243603 10918
rect 339534 8196 339540 8260
rect 339604 8258 339610 8260
rect 339953 8258 340019 8261
rect 339604 8256 340019 8258
rect 339604 8200 339958 8256
rect 340014 8200 340019 8256
rect 339604 8198 340019 8200
rect 339604 8196 339610 8198
rect 339953 8195 340019 8198
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 193806 3980 193812 4044
rect 193876 4042 193882 4044
rect 240501 4042 240567 4045
rect 193876 4040 240567 4042
rect 193876 3984 240506 4040
rect 240562 3984 240567 4040
rect 193876 3982 240567 3984
rect 193876 3980 193882 3982
rect 240501 3979 240567 3982
rect 171961 3498 172027 3501
rect 178534 3498 178540 3500
rect 171961 3496 178540 3498
rect 171961 3440 171966 3496
rect 172022 3440 178540 3496
rect 171961 3438 178540 3440
rect 171961 3435 172027 3438
rect 178534 3436 178540 3438
rect 178604 3436 178610 3500
rect 304349 3498 304415 3501
rect 304758 3498 304764 3500
rect 304349 3496 304764 3498
rect 304349 3440 304354 3496
rect 304410 3440 304764 3496
rect 304349 3438 304764 3440
rect 304349 3435 304415 3438
rect 304758 3436 304764 3438
rect 304828 3436 304834 3500
rect 195094 3300 195100 3364
rect 195164 3362 195170 3364
rect 242985 3362 243051 3365
rect 195164 3360 243051 3362
rect 195164 3304 242990 3360
rect 243046 3304 243051 3360
rect 195164 3302 243051 3304
rect 195164 3300 195170 3302
rect 242985 3299 243051 3302
<< via3 >>
rect 81020 702612 81084 702676
rect 68876 702476 68940 702540
rect 89300 699756 89364 699820
rect 70900 681804 70964 681868
rect 84700 680580 84764 680644
rect 72924 680444 72988 680508
rect 77156 680444 77220 680508
rect 82492 680444 82556 680508
rect 86724 680444 86788 680508
rect 99052 680444 99116 680508
rect 104572 680444 104636 680508
rect 75132 680308 75196 680372
rect 78260 680308 78324 680372
rect 82676 680308 82740 680372
rect 88932 680308 88996 680372
rect 101996 680308 102060 680372
rect 70348 679824 70412 679828
rect 70348 679768 70398 679824
rect 70398 679768 70412 679824
rect 70348 679764 70412 679768
rect 100524 679764 100588 679828
rect 92244 679628 92308 679692
rect 95004 679628 95068 679692
rect 97764 679628 97828 679692
rect 104756 679628 104820 679692
rect 79180 679492 79244 679556
rect 83964 679492 84028 679556
rect 90956 679492 91020 679556
rect 93716 679492 93780 679556
rect 96476 679492 96540 679556
rect 103284 679492 103348 679556
rect 106780 679492 106844 679556
rect 71820 679416 71884 679420
rect 71820 679360 71834 679416
rect 71834 679360 71884 679416
rect 71820 679356 71884 679360
rect 73108 679356 73172 679420
rect 74764 679356 74828 679420
rect 75868 679356 75932 679420
rect 78444 679356 78508 679420
rect 78812 679416 78876 679420
rect 78812 679360 78862 679416
rect 78862 679360 78876 679416
rect 78812 679356 78876 679360
rect 80100 679416 80164 679420
rect 80100 679360 80150 679416
rect 80150 679360 80164 679416
rect 80100 679356 80164 679360
rect 82860 679356 82924 679420
rect 84516 679416 84580 679420
rect 84516 679360 84530 679416
rect 84530 679360 84580 679416
rect 84516 679356 84580 679360
rect 85804 679356 85868 679420
rect 87092 679416 87156 679420
rect 87092 679360 87142 679416
rect 87142 679360 87156 679416
rect 87092 679356 87156 679360
rect 87276 679356 87340 679420
rect 91508 679416 91572 679420
rect 91508 679360 91522 679416
rect 91522 679360 91572 679416
rect 91508 679356 91572 679360
rect 92612 679356 92676 679420
rect 94084 679356 94148 679420
rect 96292 679356 96356 679420
rect 97212 679356 97276 679420
rect 98500 679416 98564 679420
rect 98500 679360 98550 679416
rect 98550 679360 98564 679416
rect 98500 679356 98564 679360
rect 99972 679416 100036 679420
rect 99972 679360 100022 679416
rect 100022 679360 100036 679416
rect 99972 679356 100036 679360
rect 101260 679416 101324 679420
rect 101260 679360 101310 679416
rect 101310 679360 101324 679416
rect 101260 679356 101324 679360
rect 102732 679356 102796 679420
rect 105492 679356 105556 679420
rect 106964 679356 107028 679420
rect 118740 676228 118804 676292
rect 68876 673100 68940 673164
rect 115980 672964 116044 673028
rect 66668 672148 66732 672212
rect 68876 672148 68940 672212
rect 109540 671604 109604 671668
rect 44036 668068 44100 668132
rect 109356 667660 109420 667724
rect 61884 662628 61948 662692
rect 111196 661676 111260 661740
rect 68692 653924 68756 653988
rect 111932 653516 111996 653580
rect 68876 648620 68940 648684
rect 66116 645900 66180 645964
rect 115796 644404 115860 644468
rect 111748 643996 111812 644060
rect 57836 643180 57900 643244
rect 81020 639840 81084 639844
rect 81020 639784 81034 639840
rect 81034 639784 81084 639840
rect 81020 639780 81084 639784
rect 108252 639780 108316 639844
rect 96292 639644 96356 639708
rect 78444 638828 78508 638892
rect 82492 638828 82556 638892
rect 84516 638828 84580 638892
rect 92244 638828 92308 638892
rect 100524 638828 100588 638892
rect 103284 638828 103348 638892
rect 108988 638828 109052 638892
rect 89300 638692 89364 638756
rect 104940 637604 105004 637668
rect 109172 637604 109236 637668
rect 55076 629852 55140 629916
rect 121684 629852 121748 629916
rect 122972 627132 123036 627196
rect 50844 624412 50908 624476
rect 92612 593404 92676 593468
rect 94084 593268 94148 593332
rect 96476 590064 96540 590068
rect 96476 590008 96490 590064
rect 96490 590008 96540 590064
rect 96476 590004 96540 590008
rect 101260 589868 101324 589932
rect 124260 589324 124324 589388
rect 78812 589188 78876 589252
rect 82860 589188 82924 589252
rect 99972 589188 100036 589252
rect 91508 588508 91572 588572
rect 120028 588508 120092 588572
rect 87092 588236 87156 588300
rect 66116 587964 66180 588028
rect 80100 587828 80164 587892
rect 97212 587888 97276 587892
rect 97212 587832 97226 587888
rect 97226 587832 97276 587888
rect 97212 587828 97276 587832
rect 106964 587888 107028 587892
rect 106964 587832 106978 587888
rect 106978 587832 107028 587888
rect 106964 587828 107028 587832
rect 79180 587692 79244 587756
rect 106780 587420 106844 587484
rect 102732 587284 102796 587348
rect 98500 587148 98564 587212
rect 73108 586468 73172 586532
rect 75868 586468 75932 586532
rect 85804 586468 85868 586532
rect 102732 586468 102796 586532
rect 48084 585516 48148 585580
rect 74764 585516 74828 585580
rect 78260 585516 78324 585580
rect 101996 585516 102060 585580
rect 105492 585576 105556 585580
rect 105492 585520 105542 585576
rect 105542 585520 105556 585576
rect 77156 585380 77220 585444
rect 84700 585380 84764 585444
rect 105492 585516 105556 585520
rect 71820 585108 71884 585172
rect 78260 585168 78324 585172
rect 78260 585112 78274 585168
rect 78274 585112 78324 585168
rect 78260 585108 78324 585112
rect 87276 585108 87340 585172
rect 88932 585168 88996 585172
rect 88932 585112 88946 585168
rect 88946 585112 88996 585168
rect 88932 585108 88996 585112
rect 90956 585108 91020 585172
rect 97764 585108 97828 585172
rect 70900 584080 70964 584084
rect 70900 584024 70950 584080
rect 70950 584024 70964 584080
rect 70900 584020 70964 584024
rect 72924 584020 72988 584084
rect 99052 584080 99116 584084
rect 99052 584024 99102 584080
rect 99102 584024 99116 584080
rect 99052 584020 99116 584024
rect 104756 584020 104820 584084
rect 75132 583884 75196 583948
rect 104572 583884 104636 583948
rect 51764 583748 51828 583812
rect 53604 583808 53668 583812
rect 53604 583752 53618 583808
rect 53618 583752 53668 583808
rect 53604 583748 53668 583752
rect 83964 583808 84028 583812
rect 83964 583752 84014 583808
rect 84014 583752 84028 583808
rect 83964 583748 84028 583752
rect 86724 583748 86788 583812
rect 93716 583808 93780 583812
rect 93716 583752 93766 583808
rect 93766 583752 93780 583808
rect 93716 583748 93780 583752
rect 107516 582720 107580 582724
rect 107516 582664 107566 582720
rect 107566 582664 107580 582720
rect 107516 582660 107580 582664
rect 95004 582524 95068 582588
rect 128676 582524 128740 582588
rect 118004 582388 118068 582452
rect 58940 581980 59004 582044
rect 82676 581980 82740 582044
rect 125732 581844 125796 581908
rect 122052 581572 122116 581636
rect 70164 581224 70228 581228
rect 70164 581168 70214 581224
rect 70214 581168 70228 581224
rect 70164 581164 70228 581168
rect 122604 579668 122668 579732
rect 70348 579260 70412 579324
rect 107516 578716 107580 578780
rect 64644 578444 64708 578508
rect 70348 578444 70412 578508
rect 62988 578172 63052 578236
rect 117084 578172 117148 578236
rect 118740 578172 118804 578236
rect 118740 577492 118804 577556
rect 107516 576132 107580 576196
rect 115980 576132 116044 576196
rect 61700 575316 61764 575380
rect 114508 575044 114572 575108
rect 115980 574636 116044 574700
rect 60596 573956 60660 574020
rect 122972 572792 123036 572796
rect 122972 572736 122986 572792
rect 122986 572736 123036 572792
rect 122972 572732 123036 572736
rect 66668 572324 66732 572388
rect 66116 570964 66180 571028
rect 108804 570692 108868 570756
rect 108252 570420 108316 570484
rect 44036 568516 44100 568580
rect 113220 568516 113284 568580
rect 111196 564980 111260 565044
rect 58756 561852 58820 561916
rect 61884 561852 61948 561916
rect 107884 558452 107948 558516
rect 111564 558180 111628 558244
rect 121684 558180 121748 558244
rect 105492 556684 105556 556748
rect 107700 556412 107764 556476
rect 111932 556412 111996 556476
rect 68692 554644 68756 554708
rect 56548 553420 56612 553484
rect 122236 549884 122300 549948
rect 68876 549204 68940 549268
rect 111748 546892 111812 546956
rect 61332 546348 61396 546412
rect 65932 546136 65996 546140
rect 65932 546080 65982 546136
rect 65982 546080 65996 546136
rect 65932 546076 65996 546080
rect 115796 545124 115860 545188
rect 55076 544308 55140 544372
rect 57836 542948 57900 543012
rect 109172 542812 109236 542876
rect 65932 541724 65996 541788
rect 104940 539820 105004 539884
rect 50844 539412 50908 539476
rect 70348 538732 70412 538796
rect 125732 538732 125796 538796
rect 58940 537372 59004 537436
rect 70164 536692 70228 536756
rect 111564 536692 111628 536756
rect 114692 536284 114756 536348
rect 125548 535468 125612 535532
rect 50844 534108 50908 534172
rect 54892 533836 54956 533900
rect 56548 533836 56612 533900
rect 55076 533624 55140 533628
rect 55076 533568 55090 533624
rect 55090 533568 55140 533624
rect 55076 533564 55140 533568
rect 114508 533292 114572 533356
rect 125548 532204 125612 532268
rect 120028 532068 120092 532132
rect 128676 531932 128740 531996
rect 65932 525676 65996 525740
rect 65932 524452 65996 524516
rect 118924 498748 118988 498812
rect 122052 498204 122116 498268
rect 115980 497388 116044 497452
rect 110644 496028 110708 496092
rect 124260 495544 124324 495548
rect 124260 495488 124310 495544
rect 124310 495488 124324 495544
rect 124260 495484 124324 495488
rect 118004 494668 118068 494732
rect 113220 493308 113284 493372
rect 57836 492764 57900 492828
rect 53604 492628 53668 492692
rect 112300 492764 112364 492828
rect 118740 492492 118804 492556
rect 99236 491404 99300 491468
rect 111564 491132 111628 491196
rect 101260 490044 101324 490108
rect 48084 489772 48148 489836
rect 50292 488548 50356 488612
rect 51764 488548 51828 488612
rect 122604 488412 122668 488476
rect 99328 485964 99392 486028
rect 117084 485692 117148 485756
rect 70348 484604 70412 484668
rect 107516 484468 107580 484532
rect 123340 484468 123404 484532
rect 107516 483108 107580 483172
rect 107516 482972 107580 483036
rect 107516 481748 107580 481812
rect 64644 481476 64708 481540
rect 106780 481476 106844 481540
rect 105492 480116 105556 480180
rect 105492 479088 105556 479092
rect 105492 479032 105542 479088
rect 105542 479032 105556 479088
rect 105492 479028 105556 479032
rect 107884 478892 107948 478956
rect 62988 477592 63052 477596
rect 62988 477536 63038 477592
rect 63038 477536 63052 477592
rect 62988 477532 63052 477536
rect 61700 476308 61764 476372
rect 62988 476308 63052 476372
rect 59124 473452 59188 473516
rect 66668 473724 66732 473788
rect 60596 473316 60660 473380
rect 66116 471548 66180 471612
rect 114692 469236 114756 469300
rect 64092 467876 64156 467940
rect 107700 467876 107764 467940
rect 104020 465624 104084 465628
rect 104020 465568 104070 465624
rect 104070 465568 104084 465624
rect 104020 465564 104084 465568
rect 58756 463524 58820 463588
rect 58940 462224 59004 462228
rect 58940 462168 58990 462224
rect 58990 462168 59004 462224
rect 58940 462164 59004 462168
rect 58940 461484 59004 461548
rect 118740 459640 118804 459644
rect 118740 459584 118790 459640
rect 118790 459584 118804 459640
rect 118740 459580 118804 459584
rect 122236 456044 122300 456108
rect 132540 456044 132604 456108
rect 68876 453868 68940 453932
rect 118740 453248 118804 453252
rect 118740 453192 118790 453248
rect 118790 453192 118804 453248
rect 118740 453188 118804 453192
rect 128860 453188 128924 453252
rect 112300 452508 112364 452572
rect 61884 447264 61948 447268
rect 61884 447208 61898 447264
rect 61898 447208 61948 447264
rect 61884 447204 61948 447208
rect 61332 445980 61396 446044
rect 65380 445708 65444 445772
rect 51580 442444 51644 442508
rect 69796 442580 69860 442644
rect 99420 442444 99484 442508
rect 121684 441628 121748 441692
rect 99052 439860 99116 439924
rect 124260 439316 124324 439380
rect 54892 438908 54956 438972
rect 106780 438636 106844 438700
rect 59124 438092 59188 438156
rect 69060 438092 69124 438156
rect 50844 437412 50908 437476
rect 118924 437412 118988 437476
rect 70348 437276 70412 437340
rect 110644 437276 110708 437340
rect 55076 435916 55140 435980
rect 129780 407764 129844 407828
rect 338252 407084 338316 407148
rect 331260 406268 331324 406332
rect 180012 405724 180076 405788
rect 127020 404908 127084 404972
rect 342300 404364 342364 404428
rect 64092 401644 64156 401708
rect 120028 402188 120092 402252
rect 339540 401644 339604 401708
rect 125732 400828 125796 400892
rect 101260 400284 101324 400348
rect 345060 397428 345124 397492
rect 104020 396612 104084 396676
rect 118740 395388 118804 395452
rect 170260 395252 170324 395316
rect 68692 394708 68756 394772
rect 57836 393892 57900 393956
rect 118924 393892 118988 393956
rect 114508 391172 114572 391236
rect 50292 390764 50356 390828
rect 111564 390764 111628 390828
rect 166212 390628 166276 390692
rect 69612 389812 69676 389876
rect 61700 389268 61764 389332
rect 68876 389132 68940 389196
rect 122052 388316 122116 388380
rect 191236 388316 191300 388380
rect 53604 387908 53668 387972
rect 121868 387772 121932 387836
rect 122604 386956 122668 387020
rect 340828 385596 340892 385660
rect 61884 385052 61948 385116
rect 177252 385188 177316 385252
rect 62988 380972 63052 381036
rect 60596 380836 60660 380900
rect 68692 380700 68756 380764
rect 60596 379476 60660 379540
rect 349108 379476 349172 379540
rect 123340 378660 123404 378724
rect 69060 378524 69124 378588
rect 115428 377496 115492 377500
rect 115428 377440 115478 377496
rect 115478 377440 115492 377496
rect 115428 377436 115492 377440
rect 59124 376892 59188 376956
rect 66116 376892 66180 376956
rect 188292 374580 188356 374644
rect 324268 371316 324332 371380
rect 61884 367100 61948 367164
rect 60596 366964 60660 367028
rect 326660 365740 326724 365804
rect 58940 364380 59004 364444
rect 198596 364516 198660 364580
rect 332548 364380 332612 364444
rect 184060 363564 184124 363628
rect 196572 363156 196636 363220
rect 334020 363156 334084 363220
rect 328500 363020 328564 363084
rect 195100 362340 195164 362404
rect 199332 362204 199396 362268
rect 200620 361660 200684 361724
rect 121684 361524 121748 361588
rect 320220 360436 320284 360500
rect 118924 360164 118988 360228
rect 173020 359348 173084 359412
rect 321508 359076 321572 359140
rect 198780 358804 198844 358868
rect 320036 358804 320100 358868
rect 68876 356900 68940 356964
rect 69612 356628 69676 356692
rect 320036 356628 320100 356692
rect 494100 356628 494164 356692
rect 133828 353424 133892 353428
rect 133828 353368 133878 353424
rect 133878 353368 133892 353424
rect 133828 353364 133892 353368
rect 327028 353364 327092 353428
rect 66668 352548 66732 352612
rect 191052 351052 191116 351116
rect 178540 349692 178604 349756
rect 198780 349692 198844 349756
rect 186820 348468 186884 348532
rect 192340 348332 192404 348396
rect 66116 347712 66180 347716
rect 66116 347656 66166 347712
rect 66166 347656 66180 347712
rect 66116 347652 66180 347656
rect 118740 347652 118804 347716
rect 132540 347712 132604 347716
rect 132540 347656 132590 347712
rect 132590 347656 132604 347712
rect 132540 347652 132604 347656
rect 65380 347244 65444 347308
rect 200620 346292 200684 346356
rect 128860 342212 128924 342276
rect 122604 339628 122668 339692
rect 199332 339356 199396 339420
rect 125732 335276 125796 335340
rect 120028 335140 120092 335204
rect 127020 333916 127084 333980
rect 195100 333236 195164 333300
rect 69244 331196 69308 331260
rect 188476 331256 188540 331260
rect 188476 331200 188526 331256
rect 188526 331200 188540 331256
rect 188476 331196 188540 331200
rect 121868 327660 121932 327724
rect 69060 320724 69124 320788
rect 160692 318004 160756 318068
rect 129780 317324 129844 317388
rect 129780 316100 129844 316164
rect 193812 315284 193876 315348
rect 124260 314664 124324 314668
rect 124260 314608 124310 314664
rect 124310 314608 124324 314664
rect 124260 314604 124324 314608
rect 324268 311748 324332 311812
rect 152412 311068 152476 311132
rect 125732 308348 125796 308412
rect 195100 305628 195164 305692
rect 144132 302772 144196 302836
rect 70900 300868 70964 300932
rect 53604 298692 53668 298756
rect 196572 294476 196636 294540
rect 124812 292572 124876 292636
rect 69244 289444 69308 289508
rect 196572 284820 196636 284884
rect 70532 284004 70596 284068
rect 123340 279380 123404 279444
rect 57836 278896 57900 278900
rect 57836 278840 57850 278896
rect 57850 278840 57900 278896
rect 57836 278836 57900 278840
rect 125732 264012 125796 264076
rect 324268 258300 324332 258364
rect 70164 258028 70228 258092
rect 120580 253132 120644 253196
rect 61700 252724 61764 252788
rect 319300 252996 319364 253060
rect 195836 250820 195900 250884
rect 195836 250412 195900 250476
rect 197124 244020 197188 244084
rect 123340 243476 123404 243540
rect 70532 242388 70596 242452
rect 196020 242116 196084 242180
rect 120580 241436 120644 241500
rect 120028 241164 120092 241228
rect 200620 240756 200684 240820
rect 70532 240212 70596 240276
rect 330340 240076 330404 240140
rect 327212 239940 327276 240004
rect 196020 238716 196084 238780
rect 71084 238580 71148 238644
rect 188476 237900 188540 237964
rect 255268 236540 255332 236604
rect 160692 235860 160756 235924
rect 57836 234500 57900 234564
rect 133828 234364 133892 234428
rect 200620 234228 200684 234292
rect 318748 231644 318812 231708
rect 324268 230420 324332 230484
rect 70900 228924 70964 228988
rect 198596 228924 198660 228988
rect 198596 228244 198660 228308
rect 180012 227020 180076 227084
rect 252508 226884 252572 226948
rect 120028 224164 120092 224228
rect 271092 222804 271156 222868
rect 195836 218588 195900 218652
rect 335860 215868 335924 215932
rect 170260 211924 170324 211988
rect 197124 211788 197188 211852
rect 144132 210428 144196 210492
rect 268332 210428 268396 210492
rect 263548 210292 263612 210356
rect 273852 204852 273916 204916
rect 124812 200636 124876 200700
rect 263732 200636 263796 200700
rect 259500 199276 259564 199340
rect 69060 195196 69124 195260
rect 258580 192612 258644 192676
rect 258396 192476 258460 192540
rect 152412 191116 152476 191180
rect 503668 190980 503732 191044
rect 259684 189620 259748 189684
rect 266308 188260 266372 188324
rect 249380 186900 249444 186964
rect 262260 185540 262324 185604
rect 321324 184180 321388 184244
rect 166212 181460 166276 181524
rect 331444 181460 331508 181524
rect 260972 180100 261036 180164
rect 269068 179964 269132 180028
rect 255452 178876 255516 178940
rect 256740 178740 256804 178804
rect 262444 178604 262508 178668
rect 502380 178604 502444 178668
rect 166396 178060 166460 178124
rect 113220 177924 113284 177988
rect 100708 177652 100772 177716
rect 105676 177712 105740 177716
rect 105676 177656 105726 177712
rect 105726 177656 105740 177712
rect 105676 177652 105740 177656
rect 106964 177652 107028 177716
rect 110644 177712 110708 177716
rect 110644 177656 110694 177712
rect 110694 177656 110708 177712
rect 110644 177652 110708 177656
rect 116900 177712 116964 177716
rect 116900 177656 116950 177712
rect 116950 177656 116964 177712
rect 116900 177652 116964 177656
rect 119476 177652 119540 177716
rect 120764 177652 120828 177716
rect 123156 177652 123220 177716
rect 127020 177652 127084 177716
rect 129412 177712 129476 177716
rect 129412 177656 129462 177712
rect 129462 177656 129476 177712
rect 129412 177652 129476 177656
rect 130700 177652 130764 177716
rect 132356 177712 132420 177716
rect 132356 177656 132406 177712
rect 132406 177656 132420 177712
rect 132356 177652 132420 177656
rect 321692 177380 321756 177444
rect 104572 177108 104636 177172
rect 115796 177168 115860 177172
rect 115796 177112 115846 177168
rect 115846 177112 115860 177168
rect 109540 176972 109604 177036
rect 115796 177108 115860 177112
rect 125732 177108 125796 177172
rect 134380 177108 134444 177172
rect 97028 176700 97092 176764
rect 166212 176836 166276 176900
rect 108068 176760 108132 176764
rect 108068 176704 108118 176760
rect 108118 176704 108132 176760
rect 108068 176700 108132 176704
rect 112116 176700 112180 176764
rect 114324 176760 114388 176764
rect 114324 176704 114374 176760
rect 114374 176704 114388 176760
rect 114324 176700 114388 176704
rect 124444 176760 124508 176764
rect 124444 176704 124494 176760
rect 124494 176704 124508 176760
rect 124444 176700 124508 176704
rect 133092 176760 133156 176764
rect 133092 176704 133142 176760
rect 133142 176704 133156 176760
rect 133092 176700 133156 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 148180 176760 148244 176764
rect 148180 176704 148230 176760
rect 148230 176704 148244 176760
rect 148180 176700 148244 176704
rect 158852 176760 158916 176764
rect 158852 176704 158902 176760
rect 158902 176704 158916 176760
rect 158852 176700 158916 176704
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176428 128188 176492
rect 166948 175884 167012 175948
rect 249196 175884 249260 175948
rect 320220 175748 320284 175812
rect 306972 175612 307036 175676
rect 98316 175400 98380 175404
rect 98316 175344 98366 175400
rect 98366 175344 98380 175400
rect 98316 175340 98380 175344
rect 101996 175400 102060 175404
rect 101996 175344 102046 175400
rect 102046 175344 102060 175400
rect 101996 175340 102060 175344
rect 118372 175400 118436 175404
rect 118372 175344 118422 175400
rect 118422 175344 118436 175400
rect 118372 175340 118436 175344
rect 121868 175400 121932 175404
rect 121868 175344 121918 175400
rect 121918 175344 121932 175400
rect 121868 175340 121932 175344
rect 496860 174388 496924 174452
rect 249380 174252 249444 174316
rect 249196 173300 249260 173364
rect 334572 172484 334636 172548
rect 495940 172212 496004 172276
rect 331444 171124 331508 171188
rect 321324 170580 321388 170644
rect 336044 169764 336108 169828
rect 494284 169764 494348 169828
rect 258396 168404 258460 168468
rect 260972 167316 261036 167380
rect 349108 167044 349172 167108
rect 503668 166908 503732 166972
rect 321692 166772 321756 166836
rect 166396 163100 166460 163164
rect 262444 163100 262508 163164
rect 256740 161060 256804 161124
rect 252508 158748 252572 158812
rect 166212 157388 166276 157452
rect 338620 157388 338684 157452
rect 334020 156436 334084 156500
rect 330340 154804 330404 154868
rect 266308 153444 266372 153508
rect 251772 149636 251836 149700
rect 254532 148276 254596 148340
rect 255268 147868 255332 147932
rect 331260 147732 331324 147796
rect 254532 145964 254596 146028
rect 306972 145556 307036 145620
rect 307708 145012 307772 145076
rect 259500 144332 259564 144396
rect 307708 143924 307772 143988
rect 327212 143924 327276 143988
rect 263732 142156 263796 142220
rect 259684 141068 259748 141132
rect 258396 140932 258460 140996
rect 255452 140388 255516 140452
rect 326660 140116 326724 140180
rect 327028 139300 327092 139364
rect 262260 138620 262324 138684
rect 253612 137124 253676 137188
rect 263548 136988 263612 137052
rect 269068 136852 269132 136916
rect 169156 135492 169220 135556
rect 170260 135356 170324 135420
rect 250300 134132 250364 134196
rect 328500 133996 328564 134060
rect 332548 133860 332612 133924
rect 502380 133860 502444 133924
rect 321508 132092 321572 132156
rect 170444 131140 170508 131204
rect 260052 130052 260116 130116
rect 494100 128964 494164 129028
rect 168972 128556 169036 128620
rect 307156 127604 307220 127668
rect 251956 123252 252020 123316
rect 302740 118084 302804 118148
rect 251772 114412 251836 114476
rect 214604 105164 214668 105228
rect 214420 103804 214484 103868
rect 305500 102852 305564 102916
rect 493916 102172 493980 102236
rect 166396 99996 166460 100060
rect 494284 99316 494348 99380
rect 324268 98500 324332 98564
rect 249196 97004 249260 97068
rect 251956 97004 252020 97068
rect 166212 96732 166276 96796
rect 304212 96868 304276 96932
rect 306972 96732 307036 96796
rect 335860 96324 335924 96388
rect 166948 95100 167012 95164
rect 493916 95100 493980 95164
rect 214604 94828 214668 94892
rect 85534 94752 85598 94756
rect 85534 94696 85578 94752
rect 85578 94696 85598 94752
rect 85534 94692 85598 94696
rect 112326 94752 112390 94756
rect 112326 94696 112350 94752
rect 112350 94696 112390 94752
rect 112326 94692 112390 94696
rect 125382 94752 125446 94756
rect 125382 94696 125414 94752
rect 125414 94696 125446 94752
rect 125382 94692 125446 94696
rect 151308 94692 151372 94756
rect 151630 94692 151694 94756
rect 126652 93876 126716 93940
rect 324268 93740 324332 93804
rect 118188 93664 118252 93668
rect 118188 93608 118238 93664
rect 118238 93608 118252 93664
rect 118188 93604 118252 93608
rect 98500 93528 98564 93532
rect 98500 93472 98550 93528
rect 98550 93472 98564 93528
rect 98500 93468 98564 93472
rect 113220 93468 113284 93532
rect 169156 93604 169220 93668
rect 129412 93528 129476 93532
rect 129412 93472 129462 93528
rect 129462 93472 129476 93528
rect 129412 93468 129476 93472
rect 133092 93528 133156 93532
rect 133092 93472 133142 93528
rect 133142 93472 133156 93528
rect 133092 93468 133156 93472
rect 151676 93528 151740 93532
rect 151676 93472 151726 93528
rect 151726 93472 151740 93528
rect 151676 93468 151740 93472
rect 103284 93256 103348 93260
rect 103284 93200 103334 93256
rect 103334 93200 103348 93256
rect 103284 93196 103348 93200
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 84332 92380 84396 92444
rect 86724 92440 86788 92444
rect 86724 92384 86774 92440
rect 86774 92384 86788 92440
rect 86724 92380 86788 92384
rect 88932 92440 88996 92444
rect 88932 92384 88982 92440
rect 88982 92384 88996 92440
rect 88932 92380 88996 92384
rect 107700 92440 107764 92444
rect 107700 92384 107750 92440
rect 107750 92384 107764 92440
rect 107700 92380 107764 92384
rect 114508 92380 114572 92444
rect 115428 92440 115492 92444
rect 115428 92384 115478 92440
rect 115478 92384 115492 92440
rect 115428 92380 115492 92384
rect 120212 92380 120276 92444
rect 121684 92380 121748 92444
rect 130700 92440 130764 92444
rect 130700 92384 130750 92440
rect 130750 92384 130764 92440
rect 130700 92380 130764 92384
rect 134380 92380 134444 92444
rect 136036 92440 136100 92444
rect 136036 92384 136086 92440
rect 136086 92384 136100 92440
rect 136036 92380 136100 92384
rect 151492 92380 151556 92444
rect 118004 92244 118068 92308
rect 166396 92244 166460 92308
rect 90220 91700 90284 91764
rect 93900 91700 93964 91764
rect 126468 91760 126532 91764
rect 126468 91704 126518 91760
rect 126518 91704 126532 91760
rect 126468 91700 126532 91704
rect 110644 91564 110708 91628
rect 101812 91488 101876 91492
rect 101812 91432 101862 91488
rect 101862 91432 101876 91488
rect 101812 91428 101876 91432
rect 122788 91488 122852 91492
rect 122788 91432 122838 91488
rect 122838 91432 122852 91488
rect 122788 91428 122852 91432
rect 152044 91428 152108 91492
rect 96660 91292 96724 91356
rect 98132 91292 98196 91356
rect 100892 91292 100956 91356
rect 106780 91292 106844 91356
rect 109172 91292 109236 91356
rect 116716 91292 116780 91356
rect 119292 91292 119356 91356
rect 74764 91156 74828 91220
rect 88012 91216 88076 91220
rect 88012 91160 88062 91216
rect 88062 91160 88076 91216
rect 88012 91156 88076 91160
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91156 95068 91220
rect 96292 91156 96356 91220
rect 97212 91156 97276 91220
rect 99052 91156 99116 91220
rect 99972 91156 100036 91220
rect 100524 91216 100588 91220
rect 100524 91160 100574 91216
rect 100574 91160 100588 91216
rect 100524 91156 100588 91160
rect 101996 91216 102060 91220
rect 101996 91160 102010 91216
rect 102010 91160 102060 91216
rect 101996 91156 102060 91160
rect 102732 91156 102796 91220
rect 104204 91156 104268 91220
rect 104572 91156 104636 91220
rect 105492 91216 105556 91220
rect 105492 91160 105542 91216
rect 105542 91160 105556 91216
rect 105492 91156 105556 91160
rect 105676 91156 105740 91220
rect 106412 91156 106476 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 111196 91216 111260 91220
rect 111196 91160 111246 91216
rect 111246 91160 111260 91216
rect 111196 91156 111260 91160
rect 111932 91156 111996 91220
rect 114324 91156 114388 91220
rect 114876 91216 114940 91220
rect 114876 91160 114926 91216
rect 114926 91160 114940 91216
rect 114876 91156 114940 91160
rect 115796 91216 115860 91220
rect 115796 91160 115846 91216
rect 115846 91160 115860 91216
rect 115796 91156 115860 91160
rect 117084 91156 117148 91220
rect 119660 91156 119724 91220
rect 120580 91216 120644 91220
rect 120580 91160 120630 91216
rect 120630 91160 120644 91216
rect 120580 91156 120644 91160
rect 122052 91156 122116 91220
rect 123156 91156 123220 91220
rect 124076 91156 124140 91220
rect 124444 91156 124508 91220
rect 125732 91156 125796 91220
rect 127572 91216 127636 91220
rect 127572 91160 127622 91216
rect 127622 91160 127636 91216
rect 127572 91156 127636 91160
rect 132356 91216 132420 91220
rect 132356 91160 132406 91216
rect 132406 91160 132420 91216
rect 132356 91156 132420 91160
rect 151308 91156 151372 91220
rect 214420 91020 214484 91084
rect 166212 88164 166276 88228
rect 170260 85444 170324 85508
rect 173020 84764 173084 84828
rect 334572 82180 334636 82244
rect 307156 82044 307220 82108
rect 170444 81364 170508 81428
rect 191236 81364 191300 81428
rect 345060 81364 345124 81428
rect 177252 79324 177316 79388
rect 168972 78508 169036 78572
rect 304764 77828 304828 77892
rect 338252 77828 338316 77892
rect 273852 76604 273916 76668
rect 304212 76468 304276 76532
rect 66668 75108 66732 75172
rect 60596 62732 60660 62796
rect 336044 62052 336108 62116
rect 260052 61508 260116 61572
rect 271092 61508 271156 61572
rect 61884 61372 61948 61436
rect 59124 59876 59188 59940
rect 302740 57156 302804 57220
rect 306972 51716 307036 51780
rect 340828 47560 340892 47564
rect 340828 47504 340878 47560
rect 340878 47504 340892 47560
rect 340828 47500 340892 47504
rect 338620 46820 338684 46884
rect 496860 46820 496924 46884
rect 268332 44780 268396 44844
rect 495940 44780 496004 44844
rect 186820 43420 186884 43484
rect 342300 41304 342364 41308
rect 342300 41248 342350 41304
rect 342350 41248 342364 41304
rect 342300 41244 342364 41248
rect 184060 40564 184124 40628
rect 191052 29548 191116 29612
rect 250300 26828 250364 26892
rect 192340 26148 192404 26212
rect 253060 25468 253124 25532
rect 188292 20572 188356 20636
rect 66116 19892 66180 19956
rect 248460 16492 248524 16556
rect 305500 12956 305564 13020
rect 340828 11732 340892 11796
rect 62988 10916 63052 10980
rect 339540 8196 339604 8260
rect 193812 3980 193876 4044
rect 178540 3436 178604 3500
rect 304764 3436 304828 3500
rect 195100 3300 195164 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 44035 668132 44101 668133
rect 44035 668068 44036 668132
rect 44100 668068 44101 668132
rect 44035 668067 44101 668068
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 44038 568581 44098 668067
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 44035 568580 44101 568581
rect 44035 568516 44036 568580
rect 44100 568516 44101 568580
rect 44035 568515 44101 568516
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 550894 45854 586338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 57835 643244 57901 643245
rect 57835 643180 57836 643244
rect 57900 643180 57901 643244
rect 57835 643179 57901 643180
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55075 629916 55141 629917
rect 55075 629852 55076 629916
rect 55140 629852 55141 629916
rect 55075 629851 55141 629852
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 50843 624476 50909 624477
rect 50843 624412 50844 624476
rect 50908 624412 50909 624476
rect 50843 624411 50909 624412
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48083 585580 48149 585581
rect 48083 585516 48084 585580
rect 48148 585516 48149 585580
rect 48083 585515 48149 585516
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 48086 489837 48146 585515
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 50846 539477 50906 624411
rect 51763 583812 51829 583813
rect 51763 583748 51764 583812
rect 51828 583748 51829 583812
rect 51763 583747 51829 583748
rect 53603 583812 53669 583813
rect 53603 583748 53604 583812
rect 53668 583748 53669 583812
rect 53603 583747 53669 583748
rect 50843 539476 50909 539477
rect 50843 539412 50844 539476
rect 50908 539412 50909 539476
rect 50843 539411 50909 539412
rect 50846 538230 50906 539411
rect 50846 538170 51642 538230
rect 50843 534172 50909 534173
rect 50843 534108 50844 534172
rect 50908 534108 50909 534172
rect 50843 534107 50909 534108
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48083 489836 48149 489837
rect 48083 489772 48084 489836
rect 48148 489772 48149 489836
rect 48083 489771 48149 489772
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 482614 49574 518058
rect 50291 488612 50357 488613
rect 50291 488548 50292 488612
rect 50356 488548 50357 488612
rect 50291 488547 50357 488548
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 50294 390829 50354 488547
rect 50846 437477 50906 534107
rect 51582 442509 51642 538170
rect 51766 488613 51826 583747
rect 53606 492693 53666 583747
rect 55078 544373 55138 629851
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55075 544372 55141 544373
rect 55075 544308 55076 544372
rect 55140 544308 55141 544372
rect 55075 544307 55141 544308
rect 54891 533900 54957 533901
rect 54891 533836 54892 533900
rect 54956 533836 54957 533900
rect 54891 533835 54957 533836
rect 53603 492692 53669 492693
rect 53603 492628 53604 492692
rect 53668 492628 53669 492692
rect 53603 492627 53669 492628
rect 51763 488612 51829 488613
rect 51763 488548 51764 488612
rect 51828 488548 51829 488612
rect 51763 488547 51829 488548
rect 51579 442508 51645 442509
rect 51579 442444 51580 442508
rect 51644 442444 51645 442508
rect 51579 442443 51645 442444
rect 50843 437476 50909 437477
rect 50843 437412 50844 437476
rect 50908 437412 50909 437476
rect 50843 437411 50909 437412
rect 50291 390828 50357 390829
rect 50291 390764 50292 390828
rect 50356 390764 50357 390828
rect 50291 390763 50357 390764
rect 53606 387973 53666 492627
rect 54894 438973 54954 533835
rect 55075 533628 55141 533629
rect 55075 533564 55076 533628
rect 55140 533564 55141 533628
rect 55075 533563 55141 533564
rect 54891 438972 54957 438973
rect 54891 438908 54892 438972
rect 54956 438908 54957 438972
rect 54891 438907 54957 438908
rect 55078 435981 55138 533563
rect 55794 525454 56414 560898
rect 56547 553484 56613 553485
rect 56547 553420 56548 553484
rect 56612 553420 56613 553484
rect 56547 553419 56613 553420
rect 56550 533901 56610 553419
rect 57838 543013 57898 643179
rect 59514 637174 60134 672618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 61883 662692 61949 662693
rect 61883 662628 61884 662692
rect 61948 662628 61949 662692
rect 61883 662627 61949 662628
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 58939 582044 59005 582045
rect 58939 581980 58940 582044
rect 59004 581980 59005 582044
rect 58939 581979 59005 581980
rect 58755 561916 58821 561917
rect 58755 561852 58756 561916
rect 58820 561852 58821 561916
rect 58755 561851 58821 561852
rect 57835 543012 57901 543013
rect 57835 542948 57836 543012
rect 57900 542948 57901 543012
rect 57835 542947 57901 542948
rect 56547 533900 56613 533901
rect 56547 533836 56548 533900
rect 56612 533836 56613 533900
rect 56547 533835 56613 533836
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 57835 492828 57901 492829
rect 57835 492764 57836 492828
rect 57900 492764 57901 492828
rect 57835 492763 57901 492764
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55075 435980 55141 435981
rect 55075 435916 55076 435980
rect 55140 435916 55141 435980
rect 55075 435915 55141 435916
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 53603 387972 53669 387973
rect 53603 387908 53604 387972
rect 53668 387908 53669 387972
rect 53603 387907 53669 387908
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 53606 298757 53666 387907
rect 55794 381454 56414 416898
rect 57838 393957 57898 492763
rect 58758 463589 58818 561851
rect 58942 537437 59002 581979
rect 59514 565174 60134 600618
rect 61699 575380 61765 575381
rect 61699 575316 61700 575380
rect 61764 575316 61765 575380
rect 61699 575315 61765 575316
rect 60595 574020 60661 574021
rect 60595 573956 60596 574020
rect 60660 573956 60661 574020
rect 60595 573955 60661 573956
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 58939 537436 59005 537437
rect 58939 537372 58940 537436
rect 59004 537372 59005 537436
rect 58939 537371 59005 537372
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59123 473516 59189 473517
rect 59123 473452 59124 473516
rect 59188 473452 59189 473516
rect 59123 473451 59189 473452
rect 58755 463588 58821 463589
rect 58755 463524 58756 463588
rect 58820 463524 58821 463588
rect 58755 463523 58821 463524
rect 58939 462228 59005 462229
rect 58939 462164 58940 462228
rect 59004 462164 59005 462228
rect 58939 462163 59005 462164
rect 58942 461549 59002 462163
rect 58939 461548 59005 461549
rect 58939 461484 58940 461548
rect 59004 461484 59005 461548
rect 58939 461483 59005 461484
rect 57835 393956 57901 393957
rect 57835 393892 57836 393956
rect 57900 393892 57901 393956
rect 57835 393891 57901 393892
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 58942 364445 59002 461483
rect 59126 438157 59186 473451
rect 59514 457174 60134 492618
rect 60598 473381 60658 573955
rect 61331 546412 61397 546413
rect 61331 546348 61332 546412
rect 61396 546348 61397 546412
rect 61331 546347 61397 546348
rect 60595 473380 60661 473381
rect 60595 473316 60596 473380
rect 60660 473316 60661 473380
rect 60595 473315 60661 473316
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59123 438156 59189 438157
rect 59123 438092 59124 438156
rect 59188 438092 59189 438156
rect 59123 438091 59189 438092
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59123 376956 59189 376957
rect 59123 376892 59124 376956
rect 59188 376892 59189 376956
rect 59123 376891 59189 376892
rect 58939 364444 59005 364445
rect 58939 364380 58940 364444
rect 59004 364380 59005 364444
rect 58939 364379 59005 364380
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 53603 298756 53669 298757
rect 53603 298692 53604 298756
rect 53668 298692 53669 298756
rect 53603 298691 53669 298692
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 273454 56414 308898
rect 57835 278900 57901 278901
rect 57835 278836 57836 278900
rect 57900 278836 57901 278900
rect 57835 278835 57901 278836
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 57838 234565 57898 278835
rect 57835 234564 57901 234565
rect 57835 234500 57836 234564
rect 57900 234500 57901 234564
rect 57835 234499 57901 234500
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 59126 59941 59186 376891
rect 59514 349174 60134 384618
rect 60598 380901 60658 473315
rect 61334 446045 61394 546347
rect 61702 476373 61762 575315
rect 61886 561917 61946 662627
rect 63234 640894 63854 676338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 68875 702540 68941 702541
rect 68875 702476 68876 702540
rect 68940 702476 68941 702540
rect 68875 702475 68941 702476
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66667 672212 66733 672213
rect 66667 672148 66668 672212
rect 66732 672148 66733 672212
rect 66667 672147 66733 672148
rect 66115 645964 66181 645965
rect 66115 645900 66116 645964
rect 66180 645900 66181 645964
rect 66115 645899 66181 645900
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 62987 578236 63053 578237
rect 62987 578172 62988 578236
rect 63052 578172 63053 578236
rect 62987 578171 63053 578172
rect 61883 561916 61949 561917
rect 61883 561852 61884 561916
rect 61948 561852 61949 561916
rect 61883 561851 61949 561852
rect 62990 477597 63050 578171
rect 63234 568894 63854 604338
rect 66118 588029 66178 645899
rect 66115 588028 66181 588029
rect 66115 587964 66116 588028
rect 66180 587964 66181 588028
rect 66115 587963 66181 587964
rect 66118 586530 66178 587963
rect 65934 586470 66178 586530
rect 64643 578508 64709 578509
rect 64643 578444 64644 578508
rect 64708 578444 64709 578508
rect 64643 578443 64709 578444
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 62987 477596 63053 477597
rect 62987 477532 62988 477596
rect 63052 477532 63053 477596
rect 62987 477531 63053 477532
rect 61699 476372 61765 476373
rect 61699 476308 61700 476372
rect 61764 476308 61765 476372
rect 61699 476307 61765 476308
rect 62987 476372 63053 476373
rect 62987 476308 62988 476372
rect 63052 476308 63053 476372
rect 62987 476307 63053 476308
rect 61883 447268 61949 447269
rect 61883 447204 61884 447268
rect 61948 447204 61949 447268
rect 61883 447203 61949 447204
rect 61331 446044 61397 446045
rect 61331 445980 61332 446044
rect 61396 445980 61397 446044
rect 61331 445979 61397 445980
rect 61699 389332 61765 389333
rect 61699 389268 61700 389332
rect 61764 389268 61765 389332
rect 61699 389267 61765 389268
rect 60595 380900 60661 380901
rect 60595 380836 60596 380900
rect 60660 380836 60661 380900
rect 60595 380835 60661 380836
rect 60598 379541 60658 380835
rect 60595 379540 60661 379541
rect 60595 379476 60596 379540
rect 60660 379476 60661 379540
rect 60595 379475 60661 379476
rect 60595 367028 60661 367029
rect 60595 366964 60596 367028
rect 60660 366964 60661 367028
rect 60595 366963 60661 366964
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 60598 62797 60658 366963
rect 61702 252789 61762 389267
rect 61886 385117 61946 447203
rect 61883 385116 61949 385117
rect 61883 385052 61884 385116
rect 61948 385052 61949 385116
rect 61883 385051 61949 385052
rect 62990 381037 63050 476307
rect 63234 460894 63854 496338
rect 64646 481541 64706 578443
rect 65934 546141 65994 586470
rect 66670 572389 66730 672147
rect 66954 644614 67574 680058
rect 68878 673165 68938 702475
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 682000 74414 686898
rect 77514 691174 78134 706202
rect 81019 702676 81085 702677
rect 81019 702612 81020 702676
rect 81084 702612 81085 702676
rect 81019 702611 81085 702612
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 682000 78134 690618
rect 70899 681868 70965 681869
rect 70899 681804 70900 681868
rect 70964 681804 70965 681868
rect 70899 681803 70965 681804
rect 70347 679828 70413 679829
rect 70347 679764 70348 679828
rect 70412 679764 70413 679828
rect 70347 679763 70413 679764
rect 68875 673164 68941 673165
rect 68875 673100 68876 673164
rect 68940 673100 68941 673164
rect 68875 673099 68941 673100
rect 68878 672213 68938 673099
rect 68875 672212 68941 672213
rect 68875 672148 68876 672212
rect 68940 672148 68941 672212
rect 68875 672147 68941 672148
rect 70350 659670 70410 679763
rect 70166 659610 70410 659670
rect 68691 653988 68757 653989
rect 68691 653924 68692 653988
rect 68756 653924 68757 653988
rect 68691 653923 68757 653924
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66667 572388 66733 572389
rect 66667 572324 66668 572388
rect 66732 572324 66733 572388
rect 66667 572323 66733 572324
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66115 571028 66181 571029
rect 66115 570964 66116 571028
rect 66180 570964 66181 571028
rect 66115 570963 66181 570964
rect 65931 546140 65997 546141
rect 65931 546076 65932 546140
rect 65996 546076 65997 546140
rect 65931 546075 65997 546076
rect 65931 541788 65997 541789
rect 65931 541724 65932 541788
rect 65996 541724 65997 541788
rect 65931 541723 65997 541724
rect 65934 525741 65994 541723
rect 65931 525740 65997 525741
rect 65931 525676 65932 525740
rect 65996 525676 65997 525740
rect 65931 525675 65997 525676
rect 65934 524517 65994 525675
rect 65931 524516 65997 524517
rect 65931 524452 65932 524516
rect 65996 524452 65997 524516
rect 65931 524451 65997 524452
rect 64643 481540 64709 481541
rect 64643 481476 64644 481540
rect 64708 481476 64709 481540
rect 64643 481475 64709 481476
rect 66118 471613 66178 570963
rect 66670 473789 66730 572323
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 68694 554709 68754 653923
rect 70166 650010 70226 659610
rect 70166 649950 70410 650010
rect 68875 648684 68941 648685
rect 68875 648620 68876 648684
rect 68940 648620 68941 648684
rect 68875 648619 68941 648620
rect 68691 554708 68757 554709
rect 68691 554644 68692 554708
rect 68756 554644 68757 554708
rect 68691 554643 68757 554644
rect 68878 549269 68938 648619
rect 70163 581228 70229 581229
rect 70163 581164 70164 581228
rect 70228 581164 70229 581228
rect 70163 581163 70229 581164
rect 68875 549268 68941 549269
rect 68875 549204 68876 549268
rect 68940 549204 68941 549268
rect 68875 549203 68941 549204
rect 70166 536757 70226 581163
rect 70350 579325 70410 649950
rect 70902 584085 70962 681803
rect 72923 680508 72989 680509
rect 72923 680444 72924 680508
rect 72988 680444 72989 680508
rect 72923 680443 72989 680444
rect 77155 680508 77221 680509
rect 77155 680444 77156 680508
rect 77220 680444 77221 680508
rect 77155 680443 77221 680444
rect 71819 679420 71885 679421
rect 71819 679356 71820 679420
rect 71884 679356 71885 679420
rect 71819 679355 71885 679356
rect 71822 585173 71882 679355
rect 71819 585172 71885 585173
rect 71819 585108 71820 585172
rect 71884 585108 71885 585172
rect 71819 585107 71885 585108
rect 72926 584085 72986 680443
rect 75131 680372 75197 680373
rect 75131 680308 75132 680372
rect 75196 680308 75197 680372
rect 75131 680307 75197 680308
rect 73107 679420 73173 679421
rect 73107 679356 73108 679420
rect 73172 679356 73173 679420
rect 73107 679355 73173 679356
rect 74763 679420 74829 679421
rect 74763 679356 74764 679420
rect 74828 679356 74829 679420
rect 74763 679355 74829 679356
rect 73110 586533 73170 679355
rect 74208 651454 74528 651486
rect 74208 651218 74250 651454
rect 74486 651218 74528 651454
rect 74208 651134 74528 651218
rect 74208 650898 74250 651134
rect 74486 650898 74528 651134
rect 74208 650866 74528 650898
rect 73794 615454 74414 638000
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73107 586532 73173 586533
rect 73107 586468 73108 586532
rect 73172 586468 73173 586532
rect 73107 586467 73173 586468
rect 70899 584084 70965 584085
rect 70899 584020 70900 584084
rect 70964 584020 70965 584084
rect 70899 584019 70965 584020
rect 72923 584084 72989 584085
rect 72923 584020 72924 584084
rect 72988 584020 72989 584084
rect 72923 584019 72989 584020
rect 73794 584000 74414 614898
rect 74766 585581 74826 679355
rect 74763 585580 74829 585581
rect 74763 585516 74764 585580
rect 74828 585516 74829 585580
rect 74763 585515 74829 585516
rect 75134 583949 75194 680307
rect 75867 679420 75933 679421
rect 75867 679356 75868 679420
rect 75932 679356 75933 679420
rect 75867 679355 75933 679356
rect 75870 586533 75930 679355
rect 75867 586532 75933 586533
rect 75867 586468 75868 586532
rect 75932 586468 75933 586532
rect 75867 586467 75933 586468
rect 77158 585445 77218 680443
rect 78259 680372 78325 680373
rect 78259 680308 78260 680372
rect 78324 680308 78325 680372
rect 78259 680307 78325 680308
rect 77514 619174 78134 638000
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77155 585444 77221 585445
rect 77155 585380 77156 585444
rect 77220 585380 77221 585444
rect 77155 585379 77221 585380
rect 77514 584000 78134 618618
rect 78262 585581 78322 680307
rect 79179 679556 79245 679557
rect 79179 679492 79180 679556
rect 79244 679492 79245 679556
rect 79179 679491 79245 679492
rect 78443 679420 78509 679421
rect 78443 679356 78444 679420
rect 78508 679356 78509 679420
rect 78443 679355 78509 679356
rect 78811 679420 78877 679421
rect 78811 679356 78812 679420
rect 78876 679356 78877 679420
rect 78811 679355 78877 679356
rect 78446 638893 78506 679355
rect 78443 638892 78509 638893
rect 78443 638828 78444 638892
rect 78508 638828 78509 638892
rect 78443 638827 78509 638828
rect 78814 589253 78874 679355
rect 78811 589252 78877 589253
rect 78811 589188 78812 589252
rect 78876 589188 78877 589252
rect 78811 589187 78877 589188
rect 79182 587757 79242 679491
rect 80099 679420 80165 679421
rect 80099 679356 80100 679420
rect 80164 679356 80165 679420
rect 80099 679355 80165 679356
rect 80102 587893 80162 679355
rect 81022 639845 81082 702611
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 682000 81854 694338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 89299 699820 89365 699821
rect 89299 699756 89300 699820
rect 89364 699756 89365 699820
rect 89299 699755 89365 699756
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 682000 85574 698058
rect 84699 680644 84765 680645
rect 84699 680580 84700 680644
rect 84764 680580 84765 680644
rect 84699 680579 84765 680580
rect 82491 680508 82557 680509
rect 82491 680444 82492 680508
rect 82556 680444 82557 680508
rect 82491 680443 82557 680444
rect 81019 639844 81085 639845
rect 81019 639780 81020 639844
rect 81084 639780 81085 639844
rect 81019 639779 81085 639780
rect 82494 638893 82554 680443
rect 82675 680372 82741 680373
rect 82675 680308 82676 680372
rect 82740 680308 82741 680372
rect 82675 680307 82741 680308
rect 82491 638892 82557 638893
rect 82491 638828 82492 638892
rect 82556 638828 82557 638892
rect 82491 638827 82557 638828
rect 81234 622894 81854 638000
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 80099 587892 80165 587893
rect 80099 587828 80100 587892
rect 80164 587828 80165 587892
rect 80099 587827 80165 587828
rect 79179 587756 79245 587757
rect 79179 587692 79180 587756
rect 79244 587692 79245 587756
rect 79179 587691 79245 587692
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 78259 585580 78325 585581
rect 78259 585516 78260 585580
rect 78324 585516 78325 585580
rect 78259 585515 78325 585516
rect 78262 585173 78322 585515
rect 78259 585172 78325 585173
rect 78259 585108 78260 585172
rect 78324 585108 78325 585172
rect 78259 585107 78325 585108
rect 81234 584000 81854 586338
rect 75131 583948 75197 583949
rect 75131 583884 75132 583948
rect 75196 583884 75197 583948
rect 75131 583883 75197 583884
rect 82678 582045 82738 680307
rect 83963 679556 84029 679557
rect 83963 679492 83964 679556
rect 84028 679492 84029 679556
rect 83963 679491 84029 679492
rect 82859 679420 82925 679421
rect 82859 679356 82860 679420
rect 82924 679356 82925 679420
rect 82859 679355 82925 679356
rect 82862 589253 82922 679355
rect 82859 589252 82925 589253
rect 82859 589188 82860 589252
rect 82924 589188 82925 589252
rect 82859 589187 82925 589188
rect 83966 583813 84026 679491
rect 84515 679420 84581 679421
rect 84515 679356 84516 679420
rect 84580 679356 84581 679420
rect 84515 679355 84581 679356
rect 84518 638893 84578 679355
rect 84515 638892 84581 638893
rect 84515 638828 84516 638892
rect 84580 638828 84581 638892
rect 84515 638827 84581 638828
rect 84702 585445 84762 680579
rect 86723 680508 86789 680509
rect 86723 680444 86724 680508
rect 86788 680444 86789 680508
rect 86723 680443 86789 680444
rect 85803 679420 85869 679421
rect 85803 679356 85804 679420
rect 85868 679356 85869 679420
rect 85803 679355 85869 679356
rect 84954 626614 85574 638000
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84699 585444 84765 585445
rect 84699 585380 84700 585444
rect 84764 585380 84765 585444
rect 84699 585379 84765 585380
rect 84954 584000 85574 590058
rect 85806 586533 85866 679355
rect 85803 586532 85869 586533
rect 85803 586468 85804 586532
rect 85868 586468 85869 586532
rect 85803 586467 85869 586468
rect 86726 583813 86786 680443
rect 88931 680372 88997 680373
rect 88931 680308 88932 680372
rect 88996 680308 88997 680372
rect 88931 680307 88997 680308
rect 87091 679420 87157 679421
rect 87091 679356 87092 679420
rect 87156 679356 87157 679420
rect 87091 679355 87157 679356
rect 87275 679420 87341 679421
rect 87275 679356 87276 679420
rect 87340 679356 87341 679420
rect 87275 679355 87341 679356
rect 87094 588301 87154 679355
rect 87091 588300 87157 588301
rect 87091 588236 87092 588300
rect 87156 588236 87157 588300
rect 87091 588235 87157 588236
rect 87278 585173 87338 679355
rect 88934 585173 88994 680307
rect 89302 638757 89362 699755
rect 91794 682000 92414 705242
rect 95514 682000 96134 707162
rect 99234 682000 99854 709082
rect 102954 682000 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 682000 110414 686898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 99051 680508 99117 680509
rect 99051 680444 99052 680508
rect 99116 680444 99117 680508
rect 99051 680443 99117 680444
rect 104571 680508 104637 680509
rect 104571 680444 104572 680508
rect 104636 680444 104637 680508
rect 104571 680443 104637 680444
rect 92243 679692 92309 679693
rect 92243 679628 92244 679692
rect 92308 679628 92309 679692
rect 92243 679627 92309 679628
rect 95003 679692 95069 679693
rect 95003 679628 95004 679692
rect 95068 679628 95069 679692
rect 95003 679627 95069 679628
rect 97763 679692 97829 679693
rect 97763 679628 97764 679692
rect 97828 679628 97829 679692
rect 97763 679627 97829 679628
rect 90955 679556 91021 679557
rect 90955 679492 90956 679556
rect 91020 679492 91021 679556
rect 90955 679491 91021 679492
rect 89568 669454 89888 669486
rect 89568 669218 89610 669454
rect 89846 669218 89888 669454
rect 89568 669134 89888 669218
rect 89568 668898 89610 669134
rect 89846 668898 89888 669134
rect 89568 668866 89888 668898
rect 89299 638756 89365 638757
rect 89299 638692 89300 638756
rect 89364 638692 89365 638756
rect 89299 638691 89365 638692
rect 90958 585173 91018 679491
rect 91507 679420 91573 679421
rect 91507 679356 91508 679420
rect 91572 679356 91573 679420
rect 91507 679355 91573 679356
rect 91510 588573 91570 679355
rect 92246 638893 92306 679627
rect 93715 679556 93781 679557
rect 93715 679492 93716 679556
rect 93780 679492 93781 679556
rect 93715 679491 93781 679492
rect 92611 679420 92677 679421
rect 92611 679356 92612 679420
rect 92676 679356 92677 679420
rect 92611 679355 92677 679356
rect 92243 638892 92309 638893
rect 92243 638828 92244 638892
rect 92308 638828 92309 638892
rect 92243 638827 92309 638828
rect 91794 633454 92414 638000
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91507 588572 91573 588573
rect 91507 588508 91508 588572
rect 91572 588508 91573 588572
rect 91507 588507 91573 588508
rect 87275 585172 87341 585173
rect 87275 585108 87276 585172
rect 87340 585108 87341 585172
rect 87275 585107 87341 585108
rect 88931 585172 88997 585173
rect 88931 585108 88932 585172
rect 88996 585108 88997 585172
rect 88931 585107 88997 585108
rect 90955 585172 91021 585173
rect 90955 585108 90956 585172
rect 91020 585108 91021 585172
rect 90955 585107 91021 585108
rect 91794 584000 92414 596898
rect 92614 593469 92674 679355
rect 92611 593468 92677 593469
rect 92611 593404 92612 593468
rect 92676 593404 92677 593468
rect 92611 593403 92677 593404
rect 93718 583813 93778 679491
rect 94083 679420 94149 679421
rect 94083 679356 94084 679420
rect 94148 679356 94149 679420
rect 94083 679355 94149 679356
rect 94086 593333 94146 679355
rect 94083 593332 94149 593333
rect 94083 593268 94084 593332
rect 94148 593268 94149 593332
rect 94083 593267 94149 593268
rect 83963 583812 84029 583813
rect 83963 583748 83964 583812
rect 84028 583748 84029 583812
rect 83963 583747 84029 583748
rect 86723 583812 86789 583813
rect 86723 583748 86724 583812
rect 86788 583748 86789 583812
rect 86723 583747 86789 583748
rect 93715 583812 93781 583813
rect 93715 583748 93716 583812
rect 93780 583748 93781 583812
rect 93715 583747 93781 583748
rect 95006 582589 95066 679627
rect 96475 679556 96541 679557
rect 96475 679492 96476 679556
rect 96540 679492 96541 679556
rect 96475 679491 96541 679492
rect 96291 679420 96357 679421
rect 96291 679356 96292 679420
rect 96356 679356 96357 679420
rect 96291 679355 96357 679356
rect 96294 639709 96354 679355
rect 96291 639708 96357 639709
rect 96291 639644 96292 639708
rect 96356 639644 96357 639708
rect 96291 639643 96357 639644
rect 95514 637174 96134 638000
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 584000 96134 600618
rect 96478 590069 96538 679491
rect 97211 679420 97277 679421
rect 97211 679356 97212 679420
rect 97276 679356 97277 679420
rect 97211 679355 97277 679356
rect 96475 590068 96541 590069
rect 96475 590004 96476 590068
rect 96540 590004 96541 590068
rect 96475 590003 96541 590004
rect 97214 587893 97274 679355
rect 97211 587892 97277 587893
rect 97211 587828 97212 587892
rect 97276 587828 97277 587892
rect 97211 587827 97277 587828
rect 97766 585173 97826 679627
rect 98499 679420 98565 679421
rect 98499 679356 98500 679420
rect 98564 679356 98565 679420
rect 98499 679355 98565 679356
rect 98502 587213 98562 679355
rect 98499 587212 98565 587213
rect 98499 587148 98500 587212
rect 98564 587148 98565 587212
rect 98499 587147 98565 587148
rect 97763 585172 97829 585173
rect 97763 585108 97764 585172
rect 97828 585108 97829 585172
rect 97763 585107 97829 585108
rect 99054 584085 99114 680443
rect 101995 680372 102061 680373
rect 101995 680308 101996 680372
rect 102060 680308 102061 680372
rect 101995 680307 102061 680308
rect 100523 679828 100589 679829
rect 100523 679764 100524 679828
rect 100588 679764 100589 679828
rect 100523 679763 100589 679764
rect 99971 679420 100037 679421
rect 99971 679356 99972 679420
rect 100036 679356 100037 679420
rect 99971 679355 100037 679356
rect 99234 604894 99854 638000
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99051 584084 99117 584085
rect 99051 584020 99052 584084
rect 99116 584020 99117 584084
rect 99051 584019 99117 584020
rect 99234 584000 99854 604338
rect 99974 589253 100034 679355
rect 100526 638893 100586 679763
rect 101259 679420 101325 679421
rect 101259 679356 101260 679420
rect 101324 679356 101325 679420
rect 101259 679355 101325 679356
rect 100523 638892 100589 638893
rect 100523 638828 100524 638892
rect 100588 638828 100589 638892
rect 100523 638827 100589 638828
rect 101262 589933 101322 679355
rect 101259 589932 101325 589933
rect 101259 589868 101260 589932
rect 101324 589868 101325 589932
rect 101259 589867 101325 589868
rect 99971 589252 100037 589253
rect 99971 589188 99972 589252
rect 100036 589188 100037 589252
rect 99971 589187 100037 589188
rect 101998 585581 102058 680307
rect 103283 679556 103349 679557
rect 103283 679492 103284 679556
rect 103348 679492 103349 679556
rect 103283 679491 103349 679492
rect 102731 679420 102797 679421
rect 102731 679356 102732 679420
rect 102796 679356 102797 679420
rect 102731 679355 102797 679356
rect 102734 587349 102794 679355
rect 103286 638893 103346 679491
rect 103283 638892 103349 638893
rect 103283 638828 103284 638892
rect 103348 638828 103349 638892
rect 103283 638827 103349 638828
rect 102954 608614 103574 638000
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102731 587348 102797 587349
rect 102731 587284 102732 587348
rect 102796 587284 102797 587348
rect 102731 587283 102797 587284
rect 102734 586533 102794 587283
rect 102731 586532 102797 586533
rect 102731 586468 102732 586532
rect 102796 586468 102797 586532
rect 102731 586467 102797 586468
rect 101995 585580 102061 585581
rect 101995 585516 101996 585580
rect 102060 585516 102061 585580
rect 101995 585515 102061 585516
rect 102954 584000 103574 608058
rect 104574 583949 104634 680443
rect 104755 679692 104821 679693
rect 104755 679628 104756 679692
rect 104820 679628 104821 679692
rect 104755 679627 104821 679628
rect 104758 584085 104818 679627
rect 106779 679556 106845 679557
rect 106779 679492 106780 679556
rect 106844 679492 106845 679556
rect 106779 679491 106845 679492
rect 105491 679420 105557 679421
rect 105491 679356 105492 679420
rect 105556 679356 105557 679420
rect 105491 679355 105557 679356
rect 104928 651454 105248 651486
rect 104928 651218 104970 651454
rect 105206 651218 105248 651454
rect 104928 651134 105248 651218
rect 104928 650898 104970 651134
rect 105206 650898 105248 651134
rect 104928 650866 105248 650898
rect 104939 637668 105005 637669
rect 104939 637604 104940 637668
rect 105004 637604 105005 637668
rect 104939 637603 105005 637604
rect 104755 584084 104821 584085
rect 104755 584020 104756 584084
rect 104820 584020 104821 584084
rect 104755 584019 104821 584020
rect 104571 583948 104637 583949
rect 104571 583884 104572 583948
rect 104636 583884 104637 583948
rect 104571 583883 104637 583884
rect 95003 582588 95069 582589
rect 95003 582524 95004 582588
rect 95068 582524 95069 582588
rect 95003 582523 95069 582524
rect 82675 582044 82741 582045
rect 82675 581980 82676 582044
rect 82740 581980 82741 582044
rect 82675 581979 82741 581980
rect 76576 579454 76896 579486
rect 70347 579324 70413 579325
rect 70347 579260 70348 579324
rect 70412 579260 70413 579324
rect 70347 579259 70413 579260
rect 70350 578509 70410 579259
rect 76576 579218 76618 579454
rect 76854 579218 76896 579454
rect 76576 579134 76896 579218
rect 76576 578898 76618 579134
rect 76854 578898 76896 579134
rect 76576 578866 76896 578898
rect 87840 579454 88160 579486
rect 87840 579218 87882 579454
rect 88118 579218 88160 579454
rect 87840 579134 88160 579218
rect 87840 578898 87882 579134
rect 88118 578898 88160 579134
rect 87840 578866 88160 578898
rect 99104 579454 99424 579486
rect 99104 579218 99146 579454
rect 99382 579218 99424 579454
rect 99104 579134 99424 579218
rect 99104 578898 99146 579134
rect 99382 578898 99424 579134
rect 99104 578866 99424 578898
rect 70347 578508 70413 578509
rect 70347 578444 70348 578508
rect 70412 578444 70413 578508
rect 70347 578443 70413 578444
rect 82208 561454 82528 561486
rect 82208 561218 82250 561454
rect 82486 561218 82528 561454
rect 82208 561134 82528 561218
rect 82208 560898 82250 561134
rect 82486 560898 82528 561134
rect 82208 560866 82528 560898
rect 93472 561454 93792 561486
rect 93472 561218 93514 561454
rect 93750 561218 93792 561454
rect 93472 561134 93792 561218
rect 93472 560898 93514 561134
rect 93750 560898 93792 561134
rect 93472 560866 93792 560898
rect 76576 543454 76896 543486
rect 76576 543218 76618 543454
rect 76854 543218 76896 543454
rect 76576 543134 76896 543218
rect 76576 542898 76618 543134
rect 76854 542898 76896 543134
rect 76576 542866 76896 542898
rect 87840 543454 88160 543486
rect 87840 543218 87882 543454
rect 88118 543218 88160 543454
rect 87840 543134 88160 543218
rect 87840 542898 87882 543134
rect 88118 542898 88160 543134
rect 87840 542866 88160 542898
rect 99104 543454 99424 543486
rect 99104 543218 99146 543454
rect 99382 543218 99424 543454
rect 99104 543134 99424 543218
rect 99104 542898 99146 543134
rect 99382 542898 99424 543134
rect 99104 542866 99424 542898
rect 104942 539885 105002 637603
rect 105494 585581 105554 679355
rect 106782 587485 106842 679491
rect 106963 679420 107029 679421
rect 106963 679356 106964 679420
rect 107028 679356 107029 679420
rect 106963 679355 107029 679356
rect 106966 587893 107026 679355
rect 109539 671668 109605 671669
rect 109539 671604 109540 671668
rect 109604 671604 109605 671668
rect 109539 671603 109605 671604
rect 109355 667724 109421 667725
rect 109355 667660 109356 667724
rect 109420 667660 109421 667724
rect 109355 667659 109421 667660
rect 109358 667450 109418 667659
rect 108806 667390 109418 667450
rect 108806 654150 108866 667390
rect 109542 663810 109602 671603
rect 108622 654090 108866 654150
rect 108990 663750 109602 663810
rect 108990 654150 109050 663750
rect 111195 661740 111261 661741
rect 111195 661676 111196 661740
rect 111260 661676 111261 661740
rect 111195 661675 111261 661676
rect 108990 654090 109234 654150
rect 108622 650010 108682 654090
rect 108438 649950 108682 650010
rect 109174 650010 109234 654090
rect 109174 649950 109602 650010
rect 108438 647250 108498 649950
rect 108438 647190 108682 647250
rect 108251 639844 108317 639845
rect 108251 639780 108252 639844
rect 108316 639780 108317 639844
rect 108251 639779 108317 639780
rect 106963 587892 107029 587893
rect 106963 587828 106964 587892
rect 107028 587828 107029 587892
rect 106963 587827 107029 587828
rect 106779 587484 106845 587485
rect 106779 587420 106780 587484
rect 106844 587420 106845 587484
rect 106779 587419 106845 587420
rect 105491 585580 105557 585581
rect 105491 585516 105492 585580
rect 105556 585516 105557 585580
rect 105491 585515 105557 585516
rect 107515 582724 107581 582725
rect 107515 582660 107516 582724
rect 107580 582660 107581 582724
rect 107515 582659 107581 582660
rect 107518 578781 107578 582659
rect 107515 578780 107581 578781
rect 107515 578716 107516 578780
rect 107580 578716 107581 578780
rect 107515 578715 107581 578716
rect 107515 576196 107581 576197
rect 107515 576132 107516 576196
rect 107580 576132 107581 576196
rect 107515 576131 107581 576132
rect 105491 556748 105557 556749
rect 105491 556684 105492 556748
rect 105556 556684 105557 556748
rect 105491 556683 105557 556684
rect 104939 539884 105005 539885
rect 104939 539820 104940 539884
rect 105004 539820 105005 539884
rect 104939 539819 105005 539820
rect 70347 538796 70413 538797
rect 70347 538732 70348 538796
rect 70412 538732 70413 538796
rect 70347 538731 70413 538732
rect 70163 536756 70229 536757
rect 70163 536692 70164 536756
rect 70228 536692 70229 536756
rect 70163 536691 70229 536692
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66667 473788 66733 473789
rect 66667 473724 66668 473788
rect 66732 473724 66733 473788
rect 66667 473723 66733 473724
rect 66115 471612 66181 471613
rect 66115 471548 66116 471612
rect 66180 471548 66181 471612
rect 66115 471547 66181 471548
rect 64091 467940 64157 467941
rect 64091 467876 64092 467940
rect 64156 467876 64157 467940
rect 64091 467875 64157 467876
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 64094 401709 64154 467875
rect 65379 445772 65445 445773
rect 65379 445708 65380 445772
rect 65444 445708 65445 445772
rect 65379 445707 65445 445708
rect 64091 401708 64157 401709
rect 64091 401644 64092 401708
rect 64156 401644 64157 401708
rect 64091 401643 64157 401644
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 62987 381036 63053 381037
rect 62987 380972 62988 381036
rect 63052 380972 63053 381036
rect 62987 380971 63053 380972
rect 61883 367164 61949 367165
rect 61883 367100 61884 367164
rect 61948 367100 61949 367164
rect 61883 367099 61949 367100
rect 61699 252788 61765 252789
rect 61699 252724 61700 252788
rect 61764 252724 61765 252788
rect 61699 252723 61765 252724
rect 60595 62796 60661 62797
rect 60595 62732 60596 62796
rect 60660 62732 60661 62796
rect 60595 62731 60661 62732
rect 61886 61437 61946 367099
rect 61883 61436 61949 61437
rect 61883 61372 61884 61436
rect 61948 61372 61949 61436
rect 61883 61371 61949 61372
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59123 59940 59189 59941
rect 59123 59876 59124 59940
rect 59188 59876 59189 59940
rect 59123 59875 59189 59876
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 62990 10981 63050 380971
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 65382 347309 65442 445707
rect 66118 376957 66178 471547
rect 66954 464614 67574 500058
rect 70350 484669 70410 538731
rect 73794 507454 74414 538000
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 492000 74414 506898
rect 77514 511174 78134 538000
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 492000 78134 510618
rect 81234 514894 81854 538000
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 492000 81854 514338
rect 84954 518614 85574 538000
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 492000 85574 518058
rect 91794 525454 92414 538000
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 492000 92414 524898
rect 95514 529174 96134 538000
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 492000 96134 492618
rect 99234 532894 99854 538000
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 492000 99854 496338
rect 102954 536614 103574 538000
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 99235 491468 99301 491469
rect 99235 491404 99236 491468
rect 99300 491404 99301 491468
rect 99235 491403 99301 491404
rect 99238 486570 99298 491403
rect 101259 490108 101325 490109
rect 101259 490044 101260 490108
rect 101324 490044 101325 490108
rect 101259 490043 101325 490044
rect 99238 486510 99390 486570
rect 99330 486029 99390 486510
rect 99327 486028 99393 486029
rect 99327 485964 99328 486028
rect 99392 485964 99393 486028
rect 99327 485963 99393 485964
rect 70347 484668 70413 484669
rect 70347 484604 70348 484668
rect 70412 484604 70413 484668
rect 70347 484603 70413 484604
rect 75576 471454 75896 471486
rect 75576 471218 75618 471454
rect 75854 471218 75896 471454
rect 75576 471134 75896 471218
rect 75576 470898 75618 471134
rect 75854 470898 75896 471134
rect 75576 470866 75896 470898
rect 84840 471454 85160 471486
rect 84840 471218 84882 471454
rect 85118 471218 85160 471454
rect 84840 471134 85160 471218
rect 84840 470898 84882 471134
rect 85118 470898 85160 471134
rect 84840 470866 85160 470898
rect 94104 471454 94424 471486
rect 94104 471218 94146 471454
rect 94382 471218 94424 471454
rect 94104 471134 94424 471218
rect 94104 470898 94146 471134
rect 94382 470898 94424 471134
rect 94104 470866 94424 470898
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 68875 453932 68941 453933
rect 68875 453868 68876 453932
rect 68940 453868 68941 453932
rect 68875 453867 68941 453868
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 392614 67574 428058
rect 68691 394772 68757 394773
rect 68691 394708 68692 394772
rect 68756 394708 68757 394772
rect 68691 394707 68757 394708
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66115 376956 66181 376957
rect 66115 376892 66116 376956
rect 66180 376892 66181 376956
rect 66115 376891 66181 376892
rect 66954 356614 67574 392058
rect 68694 380765 68754 394707
rect 68878 389197 68938 453867
rect 80208 453454 80528 453486
rect 80208 453218 80250 453454
rect 80486 453218 80528 453454
rect 80208 453134 80528 453218
rect 80208 452898 80250 453134
rect 80486 452898 80528 453134
rect 80208 452866 80528 452898
rect 89472 453454 89792 453486
rect 89472 453218 89514 453454
rect 89750 453218 89792 453454
rect 89472 453134 89792 453218
rect 89472 452898 89514 453134
rect 89750 452898 89792 453134
rect 89472 452866 89792 452898
rect 69795 442644 69861 442645
rect 69795 442580 69796 442644
rect 69860 442580 69861 442644
rect 69795 442579 69861 442580
rect 69798 442370 69858 442579
rect 99419 442508 99485 442509
rect 99419 442444 99420 442508
rect 99484 442444 99485 442508
rect 99419 442443 99485 442444
rect 99422 442370 99482 442443
rect 69798 442310 70410 442370
rect 69059 438156 69125 438157
rect 69059 438092 69060 438156
rect 69124 438092 69125 438156
rect 69059 438091 69125 438092
rect 68875 389196 68941 389197
rect 68875 389132 68876 389196
rect 68940 389132 68941 389196
rect 68875 389131 68941 389132
rect 68691 380764 68757 380765
rect 68691 380700 68692 380764
rect 68756 380700 68757 380764
rect 68691 380699 68757 380700
rect 68878 356965 68938 389131
rect 69062 378589 69122 438091
rect 70350 437341 70410 442310
rect 99054 442310 99482 442370
rect 99054 439925 99114 442310
rect 99051 439924 99117 439925
rect 99051 439860 99052 439924
rect 99116 439860 99117 439924
rect 99051 439859 99117 439860
rect 70347 437340 70413 437341
rect 70347 437276 70348 437340
rect 70412 437276 70413 437340
rect 70347 437275 70413 437276
rect 73794 435454 74414 438000
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 69611 389876 69677 389877
rect 69611 389812 69612 389876
rect 69676 389812 69677 389876
rect 69611 389811 69677 389812
rect 69059 378588 69125 378589
rect 69059 378524 69060 378588
rect 69124 378524 69125 378588
rect 69059 378523 69125 378524
rect 68875 356964 68941 356965
rect 68875 356900 68876 356964
rect 68940 356900 68941 356964
rect 68875 356899 68941 356900
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 352612 66733 352613
rect 66667 352548 66668 352612
rect 66732 352548 66733 352612
rect 66667 352547 66733 352548
rect 66115 347716 66181 347717
rect 66115 347652 66116 347716
rect 66180 347652 66181 347716
rect 66115 347651 66181 347652
rect 65379 347308 65445 347309
rect 65379 347244 65380 347308
rect 65444 347244 65445 347308
rect 65379 347243 65445 347244
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 62987 10980 63053 10981
rect 62987 10916 62988 10980
rect 63052 10916 63053 10980
rect 62987 10915 63053 10916
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 28338
rect 66118 19957 66178 347651
rect 66670 75173 66730 352547
rect 66954 320614 67574 356058
rect 69062 320789 69122 378523
rect 69614 356693 69674 389811
rect 73794 388000 74414 398898
rect 77514 403174 78134 438000
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 388000 78134 402618
rect 81234 406894 81854 438000
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 388000 81854 406338
rect 84954 410614 85574 438000
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 388000 85574 410058
rect 91794 417454 92414 438000
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 388000 92414 416898
rect 95514 421174 96134 438000
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 388000 96134 420618
rect 99234 424894 99854 438000
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 388894 99854 424338
rect 101262 400349 101322 490043
rect 102954 464614 103574 500058
rect 105494 480181 105554 556683
rect 107518 484533 107578 576131
rect 108254 570485 108314 639779
rect 108622 637590 108682 647190
rect 109542 640350 109602 649950
rect 108990 640290 109602 640350
rect 108990 638893 109050 640290
rect 108987 638892 109053 638893
rect 108987 638828 108988 638892
rect 109052 638828 109053 638892
rect 108987 638827 109053 638828
rect 109171 637668 109237 637669
rect 109171 637604 109172 637668
rect 109236 637604 109237 637668
rect 109171 637603 109237 637604
rect 108622 637530 108866 637590
rect 108806 570757 108866 637530
rect 108803 570756 108869 570757
rect 108803 570692 108804 570756
rect 108868 570692 108869 570756
rect 108803 570691 108869 570692
rect 108251 570484 108317 570485
rect 108251 570420 108252 570484
rect 108316 570420 108317 570484
rect 108251 570419 108317 570420
rect 107883 558516 107949 558517
rect 107883 558452 107884 558516
rect 107948 558452 107949 558516
rect 107883 558451 107949 558452
rect 107699 556476 107765 556477
rect 107699 556412 107700 556476
rect 107764 556412 107765 556476
rect 107699 556411 107765 556412
rect 107515 484532 107581 484533
rect 107515 484468 107516 484532
rect 107580 484468 107581 484532
rect 107515 484467 107581 484468
rect 107518 483173 107578 484467
rect 107515 483172 107581 483173
rect 107515 483108 107516 483172
rect 107580 483108 107581 483172
rect 107515 483107 107581 483108
rect 107515 483036 107581 483037
rect 107515 482972 107516 483036
rect 107580 482972 107581 483036
rect 107515 482971 107581 482972
rect 107518 481813 107578 482971
rect 107515 481812 107581 481813
rect 107515 481748 107516 481812
rect 107580 481748 107581 481812
rect 107515 481747 107581 481748
rect 106779 481540 106845 481541
rect 106779 481476 106780 481540
rect 106844 481476 106845 481540
rect 106779 481475 106845 481476
rect 105491 480180 105557 480181
rect 105491 480116 105492 480180
rect 105556 480116 105557 480180
rect 105491 480115 105557 480116
rect 105494 479093 105554 480115
rect 105491 479092 105557 479093
rect 105491 479028 105492 479092
rect 105556 479028 105557 479092
rect 105491 479027 105557 479028
rect 104019 465628 104085 465629
rect 104019 465564 104020 465628
rect 104084 465564 104085 465628
rect 104019 465563 104085 465564
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 101259 400348 101325 400349
rect 101259 400284 101260 400348
rect 101324 400284 101325 400348
rect 101259 400283 101325 400284
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 388000 99854 388338
rect 102954 392614 103574 428058
rect 104022 396677 104082 465563
rect 106782 438701 106842 481475
rect 107702 467941 107762 556411
rect 107886 478957 107946 558451
rect 109174 542877 109234 637603
rect 109794 615454 110414 638000
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 111198 565045 111258 661675
rect 113514 655174 114134 690618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 115979 673028 116045 673029
rect 115979 672964 115980 673028
rect 116044 672964 116045 673028
rect 115979 672963 116045 672964
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 111931 653580 111997 653581
rect 111931 653516 111932 653580
rect 111996 653516 111997 653580
rect 111931 653515 111997 653516
rect 111747 644060 111813 644061
rect 111747 643996 111748 644060
rect 111812 643996 111813 644060
rect 111747 643995 111813 643996
rect 111195 565044 111261 565045
rect 111195 564980 111196 565044
rect 111260 564980 111261 565044
rect 111195 564979 111261 564980
rect 111563 558244 111629 558245
rect 111563 558180 111564 558244
rect 111628 558180 111629 558244
rect 111563 558179 111629 558180
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109171 542876 109237 542877
rect 109171 542812 109172 542876
rect 109236 542812 109237 542876
rect 109171 542811 109237 542812
rect 109794 507454 110414 542898
rect 111566 536757 111626 558179
rect 111750 546957 111810 643995
rect 111934 556477 111994 653515
rect 113514 619174 114134 654618
rect 115795 644468 115861 644469
rect 115795 644404 115796 644468
rect 115860 644404 115861 644468
rect 115795 644403 115861 644404
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113219 568580 113285 568581
rect 113219 568516 113220 568580
rect 113284 568516 113285 568580
rect 113219 568515 113285 568516
rect 111931 556476 111997 556477
rect 111931 556412 111932 556476
rect 111996 556412 111997 556476
rect 111931 556411 111997 556412
rect 111747 546956 111813 546957
rect 111747 546892 111748 546956
rect 111812 546892 111813 546956
rect 111747 546891 111813 546892
rect 111563 536756 111629 536757
rect 111563 536692 111564 536756
rect 111628 536692 111629 536756
rect 111563 536691 111629 536692
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 107883 478956 107949 478957
rect 107883 478892 107884 478956
rect 107948 478892 107949 478956
rect 107883 478891 107949 478892
rect 109794 471454 110414 506898
rect 110643 496092 110709 496093
rect 110643 496028 110644 496092
rect 110708 496028 110709 496092
rect 110643 496027 110709 496028
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 107699 467940 107765 467941
rect 107699 467876 107700 467940
rect 107764 467876 107765 467940
rect 107699 467875 107765 467876
rect 106779 438700 106845 438701
rect 106779 438636 106780 438700
rect 106844 438636 106845 438700
rect 106779 438635 106845 438636
rect 109794 435454 110414 470898
rect 110646 437341 110706 496027
rect 113222 493373 113282 568515
rect 113514 547174 114134 582618
rect 114507 575108 114573 575109
rect 114507 575044 114508 575108
rect 114572 575044 114573 575108
rect 114507 575043 114573 575044
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 114510 533357 114570 575043
rect 115798 545189 115858 644403
rect 115982 576197 116042 672963
rect 117234 658894 117854 694338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 118739 676292 118805 676293
rect 118739 676228 118740 676292
rect 118804 676228 118805 676292
rect 118739 676227 118805 676228
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117083 578236 117149 578237
rect 117083 578172 117084 578236
rect 117148 578172 117149 578236
rect 117083 578171 117149 578172
rect 115979 576196 116045 576197
rect 115979 576132 115980 576196
rect 116044 576132 116045 576196
rect 115979 576131 116045 576132
rect 115979 574700 116045 574701
rect 115979 574636 115980 574700
rect 116044 574636 116045 574700
rect 115979 574635 116045 574636
rect 115795 545188 115861 545189
rect 115795 545124 115796 545188
rect 115860 545124 115861 545188
rect 115795 545123 115861 545124
rect 114691 536348 114757 536349
rect 114691 536284 114692 536348
rect 114756 536284 114757 536348
rect 114691 536283 114757 536284
rect 114507 533356 114573 533357
rect 114507 533292 114508 533356
rect 114572 533292 114573 533356
rect 114507 533291 114573 533292
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113219 493372 113285 493373
rect 113219 493308 113220 493372
rect 113284 493308 113285 493372
rect 113219 493307 113285 493308
rect 112299 492828 112365 492829
rect 112299 492764 112300 492828
rect 112364 492764 112365 492828
rect 112299 492763 112365 492764
rect 111563 491196 111629 491197
rect 111563 491132 111564 491196
rect 111628 491132 111629 491196
rect 111563 491131 111629 491132
rect 110643 437340 110709 437341
rect 110643 437276 110644 437340
rect 110708 437276 110709 437340
rect 110643 437275 110709 437276
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 104019 396676 104085 396677
rect 104019 396612 104020 396676
rect 104084 396612 104085 396676
rect 104019 396611 104085 396612
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 388000 103574 392058
rect 109794 388000 110414 398898
rect 111566 390829 111626 491131
rect 112302 452573 112362 492763
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 112299 452572 112365 452573
rect 112299 452508 112300 452572
rect 112364 452508 112365 452572
rect 112299 452507 112365 452508
rect 113514 439174 114134 474618
rect 114694 469301 114754 536283
rect 115982 497453 116042 574635
rect 115979 497452 116045 497453
rect 115979 497388 115980 497452
rect 116044 497388 116045 497452
rect 115979 497387 116045 497388
rect 117086 485757 117146 578171
rect 117234 550894 117854 586338
rect 118003 582452 118069 582453
rect 118003 582388 118004 582452
rect 118068 582388 118069 582452
rect 118003 582387 118069 582388
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117083 485756 117149 485757
rect 117083 485692 117084 485756
rect 117148 485692 117149 485756
rect 117083 485691 117149 485692
rect 117234 478894 117854 514338
rect 118006 494733 118066 582387
rect 118742 578237 118802 676227
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 121683 629916 121749 629917
rect 121683 629852 121684 629916
rect 121748 629852 121749 629916
rect 121683 629851 121749 629852
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120027 588572 120093 588573
rect 120027 588508 120028 588572
rect 120092 588508 120093 588572
rect 120027 588507 120093 588508
rect 118739 578236 118805 578237
rect 118739 578172 118740 578236
rect 118804 578172 118805 578236
rect 118739 578171 118805 578172
rect 118739 577556 118805 577557
rect 118739 577492 118740 577556
rect 118804 577492 118805 577556
rect 118739 577491 118805 577492
rect 118003 494732 118069 494733
rect 118003 494668 118004 494732
rect 118068 494668 118069 494732
rect 118003 494667 118069 494668
rect 118742 492557 118802 577491
rect 120030 532133 120090 588507
rect 120954 554614 121574 590058
rect 121686 558245 121746 629851
rect 122971 627196 123037 627197
rect 122971 627132 122972 627196
rect 123036 627132 123037 627196
rect 122971 627131 123037 627132
rect 122051 581636 122117 581637
rect 122051 581572 122052 581636
rect 122116 581572 122117 581636
rect 122051 581571 122117 581572
rect 121683 558244 121749 558245
rect 121683 558180 121684 558244
rect 121748 558180 121749 558244
rect 121683 558179 121749 558180
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120027 532132 120093 532133
rect 120027 532068 120028 532132
rect 120092 532068 120093 532132
rect 120027 532067 120093 532068
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 118923 498812 118989 498813
rect 118923 498748 118924 498812
rect 118988 498748 118989 498812
rect 118923 498747 118989 498748
rect 118739 492556 118805 492557
rect 118739 492492 118740 492556
rect 118804 492492 118805 492556
rect 118739 492491 118805 492492
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 114691 469300 114757 469301
rect 114691 469236 114692 469300
rect 114756 469236 114757 469300
rect 114691 469235 114757 469236
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 111563 390828 111629 390829
rect 111563 390764 111564 390828
rect 111628 390764 111629 390828
rect 111563 390763 111629 390764
rect 113514 388000 114134 402618
rect 117234 442894 117854 478338
rect 118739 459644 118805 459645
rect 118739 459580 118740 459644
rect 118804 459580 118805 459644
rect 118739 459579 118805 459580
rect 118742 453253 118802 459579
rect 118739 453252 118805 453253
rect 118739 453188 118740 453252
rect 118804 453188 118805 453252
rect 118739 453187 118805 453188
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 118926 437477 118986 498747
rect 120954 482614 121574 518058
rect 122054 498269 122114 581571
rect 122603 579732 122669 579733
rect 122603 579668 122604 579732
rect 122668 579668 122669 579732
rect 122603 579667 122669 579668
rect 122235 549948 122301 549949
rect 122235 549884 122236 549948
rect 122300 549884 122301 549948
rect 122235 549883 122301 549884
rect 122051 498268 122117 498269
rect 122051 498204 122052 498268
rect 122116 498204 122117 498268
rect 122051 498203 122117 498204
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 118923 437476 118989 437477
rect 118923 437412 118924 437476
rect 118988 437412 118989 437476
rect 118923 437411 118989 437412
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 114507 391236 114573 391237
rect 114507 391172 114508 391236
rect 114572 391172 114573 391236
rect 114507 391171 114573 391172
rect 114510 383670 114570 391171
rect 117234 388000 117854 406338
rect 120954 410614 121574 446058
rect 121683 441692 121749 441693
rect 121683 441628 121684 441692
rect 121748 441628 121749 441692
rect 121683 441627 121749 441628
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120027 402252 120093 402253
rect 120027 402188 120028 402252
rect 120092 402188 120093 402252
rect 120027 402187 120093 402188
rect 118739 395452 118805 395453
rect 118739 395388 118740 395452
rect 118804 395388 118805 395452
rect 118739 395387 118805 395388
rect 114510 383610 115490 383670
rect 89568 381454 89888 381486
rect 89568 381218 89610 381454
rect 89846 381218 89888 381454
rect 89568 381134 89888 381218
rect 89568 380898 89610 381134
rect 89846 380898 89888 381134
rect 89568 380866 89888 380898
rect 115430 377501 115490 383610
rect 115427 377500 115493 377501
rect 115427 377436 115428 377500
rect 115492 377436 115493 377500
rect 115427 377435 115493 377436
rect 74208 363454 74528 363486
rect 74208 363218 74250 363454
rect 74486 363218 74528 363454
rect 74208 363134 74528 363218
rect 74208 362898 74250 363134
rect 74486 362898 74528 363134
rect 74208 362866 74528 362898
rect 104928 363454 105248 363486
rect 104928 363218 104970 363454
rect 105206 363218 105248 363454
rect 104928 363134 105248 363218
rect 104928 362898 104970 363134
rect 105206 362898 105248 363134
rect 104928 362866 105248 362898
rect 69611 356692 69677 356693
rect 69611 356628 69612 356692
rect 69676 356628 69677 356692
rect 69611 356627 69677 356628
rect 118742 347717 118802 395387
rect 118923 393956 118989 393957
rect 118923 393892 118924 393956
rect 118988 393892 118989 393956
rect 118923 393891 118989 393892
rect 118926 360229 118986 393891
rect 118923 360228 118989 360229
rect 118923 360164 118924 360228
rect 118988 360164 118989 360228
rect 118923 360163 118989 360164
rect 118739 347716 118805 347717
rect 118739 347652 118740 347716
rect 118804 347652 118805 347716
rect 118739 347651 118805 347652
rect 89568 345454 89888 345486
rect 89568 345218 89610 345454
rect 89846 345218 89888 345454
rect 89568 345134 89888 345218
rect 89568 344898 89610 345134
rect 89846 344898 89888 345134
rect 89568 344866 89888 344898
rect 69243 331260 69309 331261
rect 69243 331196 69244 331260
rect 69308 331196 69309 331260
rect 69243 331195 69309 331196
rect 69059 320788 69125 320789
rect 69059 320724 69060 320788
rect 69124 320724 69125 320788
rect 69059 320723 69125 320724
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 69246 289509 69306 331195
rect 73794 327454 74414 338000
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 70899 300932 70965 300933
rect 70899 300868 70900 300932
rect 70964 300868 70965 300932
rect 70899 300867 70965 300868
rect 69243 289508 69309 289509
rect 69243 289444 69244 289508
rect 69308 289444 69309 289508
rect 69243 289443 69309 289444
rect 70902 287070 70962 300867
rect 73794 294000 74414 326898
rect 77514 331174 78134 338000
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 294000 78134 294618
rect 81234 334894 81854 338000
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 294000 81854 298338
rect 84954 302614 85574 338000
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 294000 85574 302058
rect 91794 309454 92414 338000
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 294000 92414 308898
rect 95514 313174 96134 338000
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 294000 96134 312618
rect 99234 316894 99854 338000
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 294000 99854 316338
rect 102954 320614 103574 338000
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 294000 103574 320058
rect 109794 327454 110414 338000
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 294000 110414 326898
rect 113514 331174 114134 338000
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 294000 114134 294618
rect 117234 334894 117854 338000
rect 120030 335205 120090 402187
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 121686 361589 121746 441627
rect 122054 388381 122114 498203
rect 122238 456109 122298 549883
rect 122606 488477 122666 579667
rect 122974 572797 123034 627131
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 124259 589388 124325 589389
rect 124259 589324 124260 589388
rect 124324 589324 124325 589388
rect 124259 589323 124325 589324
rect 122971 572796 123037 572797
rect 122971 572732 122972 572796
rect 123036 572732 123037 572796
rect 122971 572731 123037 572732
rect 124262 495549 124322 589323
rect 125731 581908 125797 581909
rect 125731 581844 125732 581908
rect 125796 581844 125797 581908
rect 125731 581843 125797 581844
rect 125734 538797 125794 581843
rect 127794 561454 128414 596898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 128675 582588 128741 582589
rect 128675 582524 128676 582588
rect 128740 582524 128741 582588
rect 128675 582523 128741 582524
rect 128678 567210 128738 582523
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 125731 538796 125797 538797
rect 125731 538732 125732 538796
rect 125796 538732 125797 538796
rect 125731 538731 125797 538732
rect 125547 535532 125613 535533
rect 125547 535468 125548 535532
rect 125612 535468 125613 535532
rect 125547 535467 125613 535468
rect 125550 532269 125610 535467
rect 125547 532268 125613 532269
rect 125547 532204 125548 532268
rect 125612 532204 125613 532268
rect 125547 532203 125613 532204
rect 127794 525454 128414 560898
rect 128494 567150 128738 567210
rect 128494 557550 128554 567150
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 128494 557490 128738 557550
rect 128678 531997 128738 557490
rect 128675 531996 128741 531997
rect 128675 531932 128676 531996
rect 128740 531932 128741 531996
rect 128675 531931 128741 531932
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 124259 495548 124325 495549
rect 124259 495484 124260 495548
rect 124324 495484 124325 495548
rect 124259 495483 124325 495484
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 122603 488476 122669 488477
rect 122603 488412 122604 488476
rect 122668 488412 122669 488476
rect 122603 488411 122669 488412
rect 123339 484532 123405 484533
rect 123339 484468 123340 484532
rect 123404 484468 123405 484532
rect 123339 484467 123405 484468
rect 122235 456108 122301 456109
rect 122235 456044 122236 456108
rect 122300 456044 122301 456108
rect 122235 456043 122301 456044
rect 122051 388380 122117 388381
rect 122051 388316 122052 388380
rect 122116 388316 122117 388380
rect 122051 388315 122117 388316
rect 121867 387836 121933 387837
rect 121867 387772 121868 387836
rect 121932 387772 121933 387836
rect 121867 387771 121933 387772
rect 121683 361588 121749 361589
rect 121683 361524 121684 361588
rect 121748 361524 121749 361588
rect 121683 361523 121749 361524
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120027 335204 120093 335205
rect 120027 335140 120028 335204
rect 120092 335140 120093 335204
rect 120027 335139 120093 335140
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 294000 117854 298338
rect 120954 302614 121574 338058
rect 121870 327725 121930 387771
rect 122603 387020 122669 387021
rect 122603 386956 122604 387020
rect 122668 386956 122669 387020
rect 122603 386955 122669 386956
rect 122606 339693 122666 386955
rect 123342 378725 123402 484467
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 127794 453134 128414 453218
rect 128859 453252 128925 453253
rect 128859 453188 128860 453252
rect 128924 453188 128925 453252
rect 128859 453187 128925 453188
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 124259 439380 124325 439381
rect 124259 439316 124260 439380
rect 124324 439316 124325 439380
rect 124259 439315 124325 439316
rect 123339 378724 123405 378725
rect 123339 378660 123340 378724
rect 123404 378660 123405 378724
rect 123339 378659 123405 378660
rect 122603 339692 122669 339693
rect 122603 339628 122604 339692
rect 122668 339628 122669 339692
rect 122603 339627 122669 339628
rect 121867 327724 121933 327725
rect 121867 327660 121868 327724
rect 121932 327660 121933 327724
rect 121867 327659 121933 327660
rect 124262 314669 124322 439315
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127019 404972 127085 404973
rect 127019 404908 127020 404972
rect 127084 404908 127085 404972
rect 127019 404907 127085 404908
rect 125731 400892 125797 400893
rect 125731 400828 125732 400892
rect 125796 400828 125797 400892
rect 125731 400827 125797 400828
rect 125734 335341 125794 400827
rect 125731 335340 125797 335341
rect 125731 335276 125732 335340
rect 125796 335276 125797 335340
rect 125731 335275 125797 335276
rect 127022 333981 127082 404907
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127019 333980 127085 333981
rect 127019 333916 127020 333980
rect 127084 333916 127085 333980
rect 127019 333915 127085 333916
rect 124259 314668 124325 314669
rect 124259 314604 124260 314668
rect 124324 314604 124325 314668
rect 124259 314603 124325 314604
rect 127794 309454 128414 344898
rect 128862 342277 128922 453187
rect 131514 421174 132134 456618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 132539 456108 132605 456109
rect 132539 456044 132540 456108
rect 132604 456044 132605 456108
rect 132539 456043 132605 456044
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 129779 407828 129845 407829
rect 129779 407764 129780 407828
rect 129844 407764 129845 407828
rect 129779 407763 129845 407764
rect 128859 342276 128925 342277
rect 128859 342212 128860 342276
rect 128924 342212 128925 342276
rect 128859 342211 128925 342212
rect 129782 317389 129842 407763
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 129779 317388 129845 317389
rect 129779 317324 129780 317388
rect 129844 317324 129845 317388
rect 129779 317323 129845 317324
rect 129782 316165 129842 317323
rect 129779 316164 129845 316165
rect 129779 316100 129780 316164
rect 129844 316100 129845 316164
rect 129779 316099 129845 316100
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 125731 308412 125797 308413
rect 125731 308348 125732 308412
rect 125796 308348 125797 308412
rect 125731 308347 125797 308348
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 294000 121574 302058
rect 124811 292636 124877 292637
rect 124811 292572 124812 292636
rect 124876 292572 124877 292636
rect 124811 292571 124877 292572
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 70534 287010 70962 287070
rect 70534 284069 70594 287010
rect 66954 248614 67574 284058
rect 70531 284068 70597 284069
rect 70531 284004 70532 284068
rect 70596 284004 70597 284068
rect 70531 284003 70597 284004
rect 123339 279444 123405 279445
rect 123339 279380 123340 279444
rect 123404 279380 123405 279444
rect 123339 279379 123405 279380
rect 89568 273454 89888 273486
rect 89568 273218 89610 273454
rect 89846 273218 89888 273454
rect 89568 273134 89888 273218
rect 89568 272898 89610 273134
rect 89846 272898 89888 273134
rect 89568 272866 89888 272898
rect 70163 258092 70229 258093
rect 70163 258028 70164 258092
rect 70228 258028 70229 258092
rect 70163 258027 70229 258028
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 70166 238770 70226 258027
rect 74208 255454 74528 255486
rect 74208 255218 74250 255454
rect 74486 255218 74528 255454
rect 74208 255134 74528 255218
rect 74208 254898 74250 255134
rect 74486 254898 74528 255134
rect 74208 254866 74528 254898
rect 104928 255454 105248 255486
rect 104928 255218 104970 255454
rect 105206 255218 105248 255454
rect 104928 255134 105248 255218
rect 104928 254898 104970 255134
rect 105206 254898 105248 255134
rect 104928 254866 105248 254898
rect 120579 253196 120645 253197
rect 120579 253132 120580 253196
rect 120644 253132 120645 253196
rect 120579 253131 120645 253132
rect 70531 242452 70597 242453
rect 70531 242388 70532 242452
rect 70596 242450 70597 242452
rect 70596 242390 71146 242450
rect 70596 242388 70597 242390
rect 70531 242387 70597 242388
rect 70531 240276 70597 240277
rect 70531 240212 70532 240276
rect 70596 240212 70597 240276
rect 70531 240211 70597 240212
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176600 67574 212058
rect 69062 238710 70226 238770
rect 70534 238770 70594 240211
rect 70534 238710 70962 238770
rect 69062 195261 69122 238710
rect 70902 228989 70962 238710
rect 71086 238645 71146 242390
rect 120582 241501 120642 253131
rect 123342 243541 123402 279379
rect 123339 243540 123405 243541
rect 123339 243476 123340 243540
rect 123404 243476 123405 243540
rect 123339 243475 123405 243476
rect 120579 241500 120645 241501
rect 120579 241436 120580 241500
rect 120644 241436 120645 241500
rect 120579 241435 120645 241436
rect 120027 241228 120093 241229
rect 120027 241164 120028 241228
rect 120092 241164 120093 241228
rect 120027 241163 120093 241164
rect 71083 238644 71149 238645
rect 71083 238580 71084 238644
rect 71148 238580 71149 238644
rect 71083 238579 71149 238580
rect 70899 228988 70965 228989
rect 70899 228924 70900 228988
rect 70964 228924 70965 228988
rect 70899 228923 70965 228924
rect 73794 219454 74414 238000
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 69059 195260 69125 195261
rect 69059 195196 69060 195260
rect 69124 195196 69125 195260
rect 69059 195195 69125 195196
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 223174 78134 238000
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 238000
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 230614 85574 238000
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 238000
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 238000
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 238000
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 176764 97093 176765
rect 97027 176700 97028 176764
rect 97092 176700 97093 176764
rect 97027 176699 97093 176700
rect 97030 175130 97090 176699
rect 99234 176600 99854 208338
rect 102954 212614 103574 238000
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177716 100773 177717
rect 100707 177652 100708 177716
rect 100772 177652 100773 177716
rect 100707 177651 100773 177652
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 98315 175404 98381 175405
rect 98315 175340 98316 175404
rect 98380 175340 98381 175404
rect 98315 175339 98381 175340
rect 96960 175070 97090 175130
rect 98318 175130 98378 175339
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177651
rect 102954 176600 103574 212058
rect 109794 219454 110414 238000
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 105675 177716 105741 177717
rect 105675 177652 105676 177716
rect 105740 177652 105741 177716
rect 105675 177651 105741 177652
rect 106963 177716 107029 177717
rect 106963 177652 106964 177716
rect 107028 177652 107029 177716
rect 106963 177651 107029 177652
rect 104571 177172 104637 177173
rect 104571 177108 104572 177172
rect 104636 177108 104637 177172
rect 104571 177107 104637 177108
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 101995 175404 102061 175405
rect 101995 175340 101996 175404
rect 102060 175340 102061 175404
rect 101995 175339 102061 175340
rect 101998 175130 102058 175339
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 177107
rect 105678 175130 105738 177651
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 177651
rect 109539 177036 109605 177037
rect 109539 176972 109540 177036
rect 109604 176972 109605 177036
rect 109539 176971 109605 176972
rect 108067 176764 108133 176765
rect 108067 176700 108068 176764
rect 108132 176700 108133 176764
rect 108067 176699 108133 176700
rect 108070 175130 108130 176699
rect 109542 175130 109602 176971
rect 109794 176600 110414 182898
rect 113514 223174 114134 238000
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113219 177988 113285 177989
rect 113219 177924 113220 177988
rect 113284 177924 113285 177988
rect 113219 177923 113285 177924
rect 110643 177716 110709 177717
rect 110643 177652 110644 177716
rect 110708 177652 110709 177716
rect 110643 177651 110709 177652
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 177651
rect 112115 176764 112181 176765
rect 112115 176700 112116 176764
rect 112180 176700 112181 176764
rect 112115 176699 112181 176700
rect 112118 175130 112178 176699
rect 113222 175130 113282 177923
rect 113514 176600 114134 186618
rect 117234 226894 117854 238000
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 120030 224229 120090 241163
rect 120954 230614 121574 238000
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120027 224228 120093 224229
rect 120027 224164 120028 224228
rect 120092 224164 120093 224228
rect 120027 224163 120093 224164
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 116899 177716 116965 177717
rect 116899 177652 116900 177716
rect 116964 177652 116965 177716
rect 116899 177651 116965 177652
rect 115795 177172 115861 177173
rect 115795 177108 115796 177172
rect 115860 177108 115861 177172
rect 115795 177107 115861 177108
rect 114323 176764 114389 176765
rect 114323 176700 114324 176764
rect 114388 176700 114389 176764
rect 114323 176699 114389 176700
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 176699
rect 115798 175130 115858 177107
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 177651
rect 117234 176600 117854 190338
rect 120954 194614 121574 230058
rect 124814 200701 124874 292571
rect 125734 264077 125794 308347
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 125731 264076 125797 264077
rect 125731 264012 125732 264076
rect 125796 264012 125797 264076
rect 125731 264011 125797 264012
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 124811 200700 124877 200701
rect 124811 200636 124812 200700
rect 124876 200636 124877 200700
rect 124811 200635 124877 200636
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 119475 177716 119541 177717
rect 119475 177652 119476 177716
rect 119540 177652 119541 177716
rect 119475 177651 119541 177652
rect 120763 177716 120829 177717
rect 120763 177652 120764 177716
rect 120828 177652 120829 177716
rect 120763 177651 120829 177652
rect 118371 175404 118437 175405
rect 118371 175340 118372 175404
rect 118436 175340 118437 175404
rect 118371 175339 118437 175340
rect 118374 175130 118434 175339
rect 119478 175130 119538 177651
rect 120766 175130 120826 177651
rect 120954 176600 121574 194058
rect 123155 177716 123221 177717
rect 123155 177652 123156 177716
rect 123220 177652 123221 177716
rect 123155 177651 123221 177652
rect 127019 177716 127085 177717
rect 127019 177652 127020 177716
rect 127084 177652 127085 177716
rect 127019 177651 127085 177652
rect 121867 175404 121933 175405
rect 121867 175340 121868 175404
rect 121932 175340 121933 175404
rect 121867 175339 121933 175340
rect 121870 175130 121930 175339
rect 123158 175130 123218 177651
rect 125731 177172 125797 177173
rect 125731 177108 125732 177172
rect 125796 177108 125797 177172
rect 125731 177107 125797 177108
rect 124443 176764 124509 176765
rect 124443 176700 124444 176764
rect 124508 176700 124509 176764
rect 124443 176699 124509 176700
rect 124446 175130 124506 176699
rect 125734 175130 125794 177107
rect 127022 175130 127082 177651
rect 127794 176600 128414 200898
rect 131514 313174 132134 348618
rect 132542 347717 132602 456043
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 133827 353428 133893 353429
rect 133827 353364 133828 353428
rect 133892 353364 133893 353428
rect 133827 353363 133893 353364
rect 132539 347716 132605 347717
rect 132539 347652 132540 347716
rect 132604 347652 132605 347716
rect 132539 347651 132605 347652
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 133830 234429 133890 353363
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 133827 234428 133893 234429
rect 133827 234364 133828 234428
rect 133892 234364 133893 234428
rect 133827 234363 133893 234364
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 177716 129477 177717
rect 129411 177652 129412 177716
rect 129476 177652 129477 177716
rect 129411 177651 129477 177652
rect 130699 177716 130765 177717
rect 130699 177652 130700 177716
rect 130764 177652 130765 177716
rect 130699 177651 130765 177652
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177651
rect 130702 175130 130762 177651
rect 131514 176600 132134 204618
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177716 132421 177717
rect 132355 177652 132356 177716
rect 132420 177652 132421 177716
rect 132355 177651 132421 177652
rect 132358 175130 132418 177651
rect 134379 177172 134445 177173
rect 134379 177108 134380 177172
rect 134444 177108 134445 177172
rect 134379 177107 134445 177108
rect 133091 176764 133157 176765
rect 133091 176700 133092 176764
rect 133156 176700 133157 176764
rect 133091 176699 133157 176700
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 176699
rect 134382 175130 134442 177107
rect 135234 176600 135854 208338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 144131 302836 144197 302837
rect 144131 302772 144132 302836
rect 144196 302772 144197 302836
rect 144131 302771 144197 302772
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 144134 210493 144194 302771
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 144131 210492 144197 210493
rect 144131 210428 144132 210492
rect 144196 210428 144197 210492
rect 144131 210427 144197 210428
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 152411 311132 152477 311133
rect 152411 311068 152412 311132
rect 152476 311068 152477 311132
rect 152411 311067 152477 311068
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 152414 191181 152474 311067
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 152411 191180 152477 191181
rect 152411 191116 152412 191180
rect 152476 191116 152477 191180
rect 152411 191115 152477 191116
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 176764 148245 176765
rect 148179 176700 148180 176764
rect 148244 176700 148245 176764
rect 148179 176699 148245 176700
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 176699
rect 149514 176600 150134 186618
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 166211 390692 166277 390693
rect 166211 390628 166212 390692
rect 166276 390628 166277 390692
rect 166211 390627 166277 390628
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 160691 318068 160757 318069
rect 160691 318004 160692 318068
rect 160756 318004 160757 318068
rect 160691 318003 160757 318004
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 160694 235925 160754 318003
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 160691 235924 160757 235925
rect 160691 235860 160692 235924
rect 160756 235860 160757 235924
rect 160691 235859 160757 235860
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 166214 181525 166274 390627
rect 167514 385174 168134 420618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 170259 395316 170325 395317
rect 170259 395252 170260 395316
rect 170324 395252 170325 395316
rect 170259 395251 170325 395252
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 170262 211989 170322 395251
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 180011 405788 180077 405789
rect 180011 405724 180012 405788
rect 180076 405724 180077 405788
rect 180011 405723 180077 405724
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 173019 359412 173085 359413
rect 173019 359348 173020 359412
rect 173084 359348 173085 359412
rect 173019 359347 173085 359348
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 170259 211988 170325 211989
rect 170259 211924 170260 211988
rect 170324 211924 170325 211988
rect 170259 211923 170325 211924
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 166211 181524 166277 181525
rect 166211 181460 166212 181524
rect 166276 181460 166277 181524
rect 166211 181459 166277 181460
rect 166395 178124 166461 178125
rect 166395 178060 166396 178124
rect 166460 178060 166461 178124
rect 166395 178059 166461 178060
rect 166211 176900 166277 176901
rect 166211 176836 166212 176900
rect 166276 176836 166277 176900
rect 166211 176835 166277 176836
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 166214 157453 166274 176835
rect 166398 163165 166458 178059
rect 166947 175948 167013 175949
rect 166947 175884 166948 175948
rect 167012 175884 167013 175948
rect 166947 175883 167013 175884
rect 166395 163164 166461 163165
rect 166395 163100 166396 163164
rect 166460 163100 166461 163164
rect 166395 163099 166461 163100
rect 166211 157452 166277 157453
rect 166211 157388 166212 157452
rect 166276 157388 166277 157452
rect 166211 157387 166277 157388
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 166395 100060 166461 100061
rect 166395 99996 166396 100060
rect 166460 99996 166461 100060
rect 166395 99995 166461 99996
rect 166211 96796 166277 96797
rect 166211 96732 166212 96796
rect 166276 96732 166277 96796
rect 166211 96731 166277 96732
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 66667 75172 66733 75173
rect 66667 75108 66668 75172
rect 66732 75108 66733 75172
rect 66667 75107 66733 75108
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 66115 19956 66181 19957
rect 66115 19892 66116 19956
rect 66180 19892 66181 19956
rect 66115 19891 66181 19892
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 92445 84394 94830
rect 85536 94757 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 85533 94756 85599 94757
rect 85533 94692 85534 94756
rect 85598 94692 85599 94756
rect 85533 94691 85599 94692
rect 84331 92444 84397 92445
rect 84331 92380 84332 92444
rect 84396 92380 84397 92444
rect 84331 92379 84397 92380
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 86726 92445 86786 94830
rect 86723 92444 86789 92445
rect 86723 92380 86724 92444
rect 86788 92380 86789 92444
rect 86723 92379 86789 92380
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 92445 88994 94830
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 90222 91765 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 90219 91764 90285 91765
rect 90219 91700 90220 91764
rect 90284 91700 90285 91764
rect 90219 91699 90285 91700
rect 91326 91221 91386 94830
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91765 93962 94830
rect 93899 91764 93965 91765
rect 93899 91700 93900 91764
rect 93964 91700 93965 91764
rect 93899 91699 93965 91700
rect 95006 91221 95066 94830
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91357 96722 94830
rect 96659 91356 96725 91357
rect 96659 91292 96660 91356
rect 96724 91292 96725 91356
rect 96659 91291 96725 91292
rect 97214 91221 97274 94830
rect 98134 91357 98194 94830
rect 98502 93533 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 98499 93532 98565 93533
rect 98499 93468 98500 93532
rect 98564 93468 98565 93532
rect 98499 93467 98565 93468
rect 98131 91356 98197 91357
rect 98131 91292 98132 91356
rect 98196 91292 98197 91356
rect 98131 91291 98197 91292
rect 99054 91221 99114 94830
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 91221 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 100526 91221 100586 94830
rect 100894 91357 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 101992 94830 102058 94890
rect 101814 91493 101874 94830
rect 101811 91492 101877 91493
rect 101811 91428 101812 91492
rect 101876 91428 101877 91492
rect 101811 91427 101877 91428
rect 100891 91356 100957 91357
rect 100891 91292 100892 91356
rect 100956 91292 100957 91356
rect 100891 91291 100957 91292
rect 101998 91221 102058 94830
rect 102734 94830 103004 94890
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 103216 94830 103346 94890
rect 102734 91221 102794 94830
rect 103286 93261 103346 94830
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 103283 93260 103349 93261
rect 103283 93196 103284 93260
rect 103348 93196 103349 93260
rect 103283 93195 103349 93196
rect 99971 91220 100037 91221
rect 99971 91156 99972 91220
rect 100036 91156 100037 91220
rect 99971 91155 100037 91156
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91221 104266 94830
rect 104574 91221 104634 94830
rect 105494 91221 105554 94830
rect 105678 91221 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 106414 91221 106474 94830
rect 106782 91357 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 107702 92445 107762 94830
rect 107699 92444 107765 92445
rect 107699 92380 107700 92444
rect 107764 92380 107765 92444
rect 107699 92379 107765 92380
rect 106779 91356 106845 91357
rect 106779 91292 106780 91356
rect 106844 91292 106845 91356
rect 106779 91291 106845 91292
rect 108070 91221 108130 94830
rect 109174 91357 109234 94830
rect 109171 91356 109237 91357
rect 109171 91292 109172 91356
rect 109236 91292 109237 91356
rect 109171 91291 109237 91292
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105491 91220 105557 91221
rect 105491 91156 105492 91220
rect 105556 91156 105557 91220
rect 105491 91155 105557 91156
rect 105675 91220 105741 91221
rect 105675 91156 105676 91220
rect 105740 91156 105741 91220
rect 105675 91155 105741 91156
rect 106411 91220 106477 91221
rect 106411 91156 106412 91220
rect 106476 91156 106477 91220
rect 106411 91155 106477 91156
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91629 110706 94830
rect 110643 91628 110709 91629
rect 110643 91564 110644 91628
rect 110708 91564 110709 91628
rect 110643 91563 110709 91564
rect 111198 91221 111258 94830
rect 111934 91221 111994 94830
rect 112328 94757 112388 95200
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 113144 94830 113282 94890
rect 113688 94830 114202 94890
rect 114368 94830 114570 94890
rect 114776 94830 114938 94890
rect 112325 94756 112391 94757
rect 112325 94692 112326 94756
rect 112390 94692 112391 94756
rect 112325 94691 112391 94692
rect 113222 93533 113282 94830
rect 114142 93870 114202 94830
rect 114142 93810 114386 93870
rect 113219 93532 113285 93533
rect 113219 93468 113220 93532
rect 113284 93468 113285 93532
rect 113219 93467 113285 93468
rect 111195 91220 111261 91221
rect 111195 91156 111196 91220
rect 111260 91156 111261 91220
rect 111195 91155 111261 91156
rect 111931 91220 111997 91221
rect 111931 91156 111932 91220
rect 111996 91156 111997 91220
rect 111931 91155 111997 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 93810
rect 114510 92445 114570 94830
rect 114507 92444 114573 92445
rect 114507 92380 114508 92444
rect 114572 92380 114573 92444
rect 114507 92379 114573 92380
rect 114878 91221 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 92445 115490 94830
rect 115427 92444 115493 92445
rect 115427 92380 115428 92444
rect 115492 92380 115493 92444
rect 115427 92379 115493 92380
rect 115798 91221 115858 94830
rect 116718 91357 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 91356 116781 91357
rect 116715 91292 116716 91356
rect 116780 91292 116781 91356
rect 116715 91291 116781 91292
rect 117086 91221 117146 94830
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 114875 91220 114941 91221
rect 114875 91156 114876 91220
rect 114940 91156 114941 91220
rect 114875 91155 114941 91156
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 92309 118066 94830
rect 118190 93669 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 118187 93668 118253 93669
rect 118187 93604 118188 93668
rect 118252 93604 118253 93668
rect 118187 93603 118253 93604
rect 118003 92308 118069 92309
rect 118003 92244 118004 92308
rect 118068 92244 118069 92308
rect 118003 92243 118069 92244
rect 119294 91357 119354 94830
rect 119291 91356 119357 91357
rect 119291 91292 119292 91356
rect 119356 91292 119357 91356
rect 119291 91291 119357 91292
rect 119662 91221 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 120214 92445 120274 94830
rect 120211 92444 120277 92445
rect 120211 92380 120212 92444
rect 120276 92380 120277 92444
rect 120211 92379 120277 92380
rect 120582 91221 120642 94830
rect 119659 91220 119725 91221
rect 119659 91156 119660 91220
rect 119724 91156 119725 91220
rect 119659 91155 119725 91156
rect 120579 91220 120645 91221
rect 120579 91156 120580 91220
rect 120644 91156 120645 91220
rect 120579 91155 120645 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 121686 92445 121746 94830
rect 121683 92444 121749 92445
rect 121683 92380 121684 92444
rect 121748 92380 121749 92444
rect 121683 92379 121749 92380
rect 122054 91221 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 123158 91221 123218 94830
rect 124078 91221 124138 94830
rect 124446 91221 124506 94830
rect 125384 94757 125444 95200
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125381 94756 125447 94757
rect 125381 94692 125382 94756
rect 125446 94692 125447 94756
rect 125381 94691 125447 94692
rect 125734 91221 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 126470 91765 126530 94830
rect 126654 93941 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 126651 93940 126717 93941
rect 126651 93876 126652 93940
rect 126716 93876 126717 93940
rect 126651 93875 126717 93876
rect 126467 91764 126533 91765
rect 126467 91700 126468 91764
rect 126532 91700 126533 91764
rect 126467 91699 126533 91700
rect 127574 91221 127634 94830
rect 129414 93533 129474 94830
rect 129411 93532 129477 93533
rect 129411 93468 129412 93532
rect 129476 93468 129477 93532
rect 129411 93467 129477 93468
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 123155 91220 123221 91221
rect 123155 91156 123156 91220
rect 123220 91156 123221 91220
rect 123155 91155 123221 91156
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 124443 91220 124509 91221
rect 124443 91156 124444 91220
rect 124508 91156 124509 91220
rect 124443 91155 124509 91156
rect 125731 91220 125797 91221
rect 125731 91156 125732 91220
rect 125796 91156 125797 91220
rect 125731 91155 125797 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 130702 92445 130762 94830
rect 130699 92444 130765 92445
rect 130699 92380 130700 92444
rect 130764 92380 130765 92444
rect 130699 92379 130765 92380
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91221 132418 94830
rect 133136 94754 133196 95200
rect 133094 94694 133196 94754
rect 134360 94754 134420 95200
rect 135584 94754 135644 95200
rect 151496 94890 151556 95200
rect 151494 94830 151556 94890
rect 151307 94756 151373 94757
rect 134360 94694 134442 94754
rect 135584 94694 136098 94754
rect 133094 93533 133154 94694
rect 133091 93532 133157 93533
rect 133091 93468 133092 93532
rect 133156 93468 133157 93532
rect 133091 93467 133157 93468
rect 134382 92445 134442 94694
rect 134379 92444 134445 92445
rect 134379 92380 134380 92444
rect 134444 92380 134445 92444
rect 134379 92379 134445 92380
rect 132355 91220 132421 91221
rect 132355 91156 132356 91220
rect 132420 91156 132421 91220
rect 132355 91155 132421 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 92445 136098 94694
rect 151307 94692 151308 94756
rect 151372 94692 151373 94756
rect 151307 94691 151373 94692
rect 136035 92444 136101 92445
rect 136035 92380 136036 92444
rect 136100 92380 136101 92444
rect 136035 92379 136101 92380
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 91221 151370 94691
rect 151494 92445 151554 94830
rect 151632 94757 151692 95200
rect 151629 94756 151695 94757
rect 151629 94692 151630 94756
rect 151694 94692 151695 94756
rect 151629 94691 151695 94692
rect 151768 94210 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151678 94150 151828 94210
rect 151678 93533 151738 94150
rect 151675 93532 151741 93533
rect 151675 93468 151676 93532
rect 151740 93468 151741 93532
rect 151675 93467 151741 93468
rect 151491 92444 151557 92445
rect 151491 92380 151492 92444
rect 151556 92380 151557 92444
rect 151491 92379 151557 92380
rect 152046 91493 152106 94830
rect 152043 91492 152109 91493
rect 152043 91428 152044 91492
rect 152108 91428 152109 91492
rect 152043 91427 152109 91428
rect 151307 91220 151373 91221
rect 151307 91156 151308 91220
rect 151372 91156 151373 91220
rect 151307 91155 151373 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 88229 166274 96731
rect 166398 92309 166458 99995
rect 166950 95165 167010 175883
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 169155 135556 169221 135557
rect 169155 135492 169156 135556
rect 169220 135492 169221 135556
rect 169155 135491 169221 135492
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 168971 128620 169037 128621
rect 168971 128556 168972 128620
rect 169036 128556 169037 128620
rect 168971 128555 169037 128556
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 166947 95164 167013 95165
rect 166947 95100 166948 95164
rect 167012 95100 167013 95164
rect 166947 95099 167013 95100
rect 166395 92308 166461 92309
rect 166395 92244 166396 92308
rect 166460 92244 166461 92308
rect 166395 92243 166461 92244
rect 166211 88228 166277 88229
rect 166211 88164 166212 88228
rect 166276 88164 166277 88228
rect 166211 88163 166277 88164
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 61174 168134 96618
rect 168974 78573 169034 128555
rect 169158 93669 169218 135491
rect 170259 135420 170325 135421
rect 170259 135356 170260 135420
rect 170324 135356 170325 135420
rect 170259 135355 170325 135356
rect 169155 93668 169221 93669
rect 169155 93604 169156 93668
rect 169220 93604 169221 93668
rect 169155 93603 169221 93604
rect 170262 85509 170322 135355
rect 170443 131204 170509 131205
rect 170443 131140 170444 131204
rect 170508 131140 170509 131204
rect 170443 131139 170509 131140
rect 170259 85508 170325 85509
rect 170259 85444 170260 85508
rect 170324 85444 170325 85508
rect 170259 85443 170325 85444
rect 170446 81429 170506 131139
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 170443 81428 170509 81429
rect 170443 81364 170444 81428
rect 170508 81364 170509 81428
rect 170443 81363 170509 81364
rect 168971 78572 169037 78573
rect 168971 78508 168972 78572
rect 169036 78508 169037 78572
rect 168971 78507 169037 78508
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 64894 171854 100338
rect 173022 84829 173082 359347
rect 174954 356614 175574 392058
rect 177251 385252 177317 385253
rect 177251 385188 177252 385252
rect 177316 385188 177317 385252
rect 177251 385187 177317 385188
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 173019 84828 173085 84829
rect 173019 84764 173020 84828
rect 173084 84764 173085 84828
rect 173019 84763 173085 84764
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 68614 175574 104058
rect 177254 79389 177314 385187
rect 178539 349756 178605 349757
rect 178539 349692 178540 349756
rect 178604 349692 178605 349756
rect 178539 349691 178605 349692
rect 177251 79388 177317 79389
rect 177251 79324 177252 79388
rect 177316 79324 177317 79388
rect 177251 79323 177317 79324
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 178542 3501 178602 349691
rect 180014 227085 180074 405723
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 188291 374644 188357 374645
rect 188291 374580 188292 374644
rect 188356 374580 188357 374644
rect 188291 374579 188357 374580
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 184059 363628 184125 363629
rect 184059 363564 184060 363628
rect 184124 363564 184125 363628
rect 184059 363563 184125 363564
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 180011 227084 180077 227085
rect 180011 227020 180012 227084
rect 180076 227020 180077 227084
rect 180011 227019 180077 227020
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 184062 40629 184122 363563
rect 185514 331174 186134 366618
rect 186819 348532 186885 348533
rect 186819 348468 186820 348532
rect 186884 348468 186885 348532
rect 186819 348467 186885 348468
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 186822 43485 186882 348467
rect 186819 43484 186885 43485
rect 186819 43420 186820 43484
rect 186884 43420 186885 43484
rect 186819 43419 186885 43420
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 184059 40628 184125 40629
rect 184059 40564 184060 40628
rect 184124 40564 184125 40628
rect 184059 40563 184125 40564
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 178539 3500 178605 3501
rect 178539 3436 178540 3500
rect 178604 3436 178605 3500
rect 178539 3435 178605 3436
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 42618
rect 188294 20637 188354 374579
rect 189234 370894 189854 406338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 191235 388380 191301 388381
rect 191235 388316 191236 388380
rect 191300 388316 191301 388380
rect 191235 388315 191301 388316
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 191051 351116 191117 351117
rect 191051 351052 191052 351116
rect 191116 351052 191117 351116
rect 191051 351051 191117 351052
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 188475 331260 188541 331261
rect 188475 331196 188476 331260
rect 188540 331196 188541 331260
rect 188475 331195 188541 331196
rect 188478 237965 188538 331195
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 188475 237964 188541 237965
rect 188475 237900 188476 237964
rect 188540 237900 188541 237964
rect 188475 237899 188541 237900
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 188291 20636 188357 20637
rect 188291 20572 188292 20636
rect 188356 20572 188357 20636
rect 188291 20571 188357 20572
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 46338
rect 191054 29613 191114 351051
rect 191238 81429 191298 388315
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192339 348396 192405 348397
rect 192339 348332 192340 348396
rect 192404 348332 192405 348396
rect 192339 348331 192405 348332
rect 191235 81428 191301 81429
rect 191235 81364 191236 81428
rect 191300 81364 191301 81428
rect 191235 81363 191301 81364
rect 191051 29612 191117 29613
rect 191051 29548 191052 29612
rect 191116 29548 191117 29612
rect 191051 29547 191117 29548
rect 192342 26213 192402 348331
rect 192954 338614 193574 374058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 198595 364580 198661 364581
rect 198595 364516 198596 364580
rect 198660 364516 198661 364580
rect 198595 364515 198661 364516
rect 196571 363220 196637 363221
rect 196571 363156 196572 363220
rect 196636 363156 196637 363220
rect 196571 363155 196637 363156
rect 195099 362404 195165 362405
rect 195099 362340 195100 362404
rect 195164 362340 195165 362404
rect 195099 362339 195165 362340
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 195102 333301 195162 362339
rect 195099 333300 195165 333301
rect 195099 333236 195100 333300
rect 195164 333236 195165 333300
rect 195099 333235 195165 333236
rect 193811 315348 193877 315349
rect 193811 315284 193812 315348
rect 193876 315284 193877 315348
rect 193811 315283 193877 315284
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192339 26212 192405 26213
rect 192339 26148 192340 26212
rect 192404 26148 192405 26212
rect 192339 26147 192405 26148
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 193814 4045 193874 315283
rect 195099 305692 195165 305693
rect 195099 305628 195100 305692
rect 195164 305628 195165 305692
rect 195099 305627 195165 305628
rect 193811 4044 193877 4045
rect 193811 3980 193812 4044
rect 193876 3980 193877 4044
rect 193811 3979 193877 3980
rect 195102 3365 195162 305627
rect 196574 294541 196634 363155
rect 196571 294540 196637 294541
rect 196571 294476 196572 294540
rect 196636 294476 196637 294540
rect 196571 294475 196637 294476
rect 196571 284884 196637 284885
rect 196571 284820 196572 284884
rect 196636 284820 196637 284884
rect 196571 284819 196637 284820
rect 196574 267750 196634 284819
rect 196574 267690 197186 267750
rect 195835 250884 195901 250885
rect 195835 250820 195836 250884
rect 195900 250820 195901 250884
rect 195835 250819 195901 250820
rect 195838 250477 195898 250819
rect 195835 250476 195901 250477
rect 195835 250412 195836 250476
rect 195900 250412 195901 250476
rect 195835 250411 195901 250412
rect 195838 218653 195898 250411
rect 197126 244085 197186 267690
rect 197123 244084 197189 244085
rect 197123 244020 197124 244084
rect 197188 244020 197189 244084
rect 197123 244019 197189 244020
rect 196019 242180 196085 242181
rect 196019 242116 196020 242180
rect 196084 242116 196085 242180
rect 196019 242115 196085 242116
rect 196022 238781 196082 242115
rect 196019 238780 196085 238781
rect 196019 238716 196020 238780
rect 196084 238716 196085 238780
rect 196019 238715 196085 238716
rect 195835 218652 195901 218653
rect 195835 218588 195836 218652
rect 195900 218588 195901 218652
rect 195835 218587 195901 218588
rect 197126 211853 197186 244019
rect 198598 228989 198658 364515
rect 199331 362268 199397 362269
rect 199331 362204 199332 362268
rect 199396 362204 199397 362268
rect 199331 362203 199397 362204
rect 198779 358868 198845 358869
rect 198779 358804 198780 358868
rect 198844 358804 198845 358868
rect 198779 358803 198845 358804
rect 198782 349757 198842 358803
rect 198779 349756 198845 349757
rect 198779 349692 198780 349756
rect 198844 349692 198845 349756
rect 198779 349691 198845 349692
rect 199334 339421 199394 362203
rect 199794 362000 200414 380898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 362000 204134 384618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 362000 207854 388338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 362000 211574 392058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 362000 218414 362898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 362000 222134 366618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 362000 225854 370338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 362000 229574 374058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 362000 236414 380898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 362000 240134 384618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 362000 243854 388338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 362000 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 362000 254414 362898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 362000 258134 366618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 362000 261854 370338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 362000 265574 374058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 362000 272414 380898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 362000 276134 384618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 362000 279854 388338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 362000 283574 392058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 362000 290414 362898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 362000 294134 366618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 362000 297854 370338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 362000 301574 374058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 362000 308414 380898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 362000 312134 384618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 362000 315854 388338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 362000 319574 392058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 324267 371380 324333 371381
rect 324267 371316 324268 371380
rect 324332 371316 324333 371380
rect 324267 371315 324333 371316
rect 200619 361724 200685 361725
rect 200619 361660 200620 361724
rect 200684 361660 200685 361724
rect 200619 361659 200685 361660
rect 200622 346357 200682 361659
rect 320219 360500 320285 360501
rect 320219 360436 320220 360500
rect 320284 360436 320285 360500
rect 320219 360435 320285 360436
rect 320035 358868 320101 358869
rect 320035 358804 320036 358868
rect 320100 358804 320101 358868
rect 320035 358803 320101 358804
rect 320038 356693 320098 358803
rect 320035 356692 320101 356693
rect 320035 356628 320036 356692
rect 320100 356628 320101 356692
rect 320035 356627 320101 356628
rect 200619 346356 200685 346357
rect 200619 346292 200620 346356
rect 200684 346292 200685 346356
rect 200619 346291 200685 346292
rect 219568 345454 219888 345486
rect 219568 345218 219610 345454
rect 219846 345218 219888 345454
rect 219568 345134 219888 345218
rect 219568 344898 219610 345134
rect 219846 344898 219888 345134
rect 219568 344866 219888 344898
rect 250288 345454 250608 345486
rect 250288 345218 250330 345454
rect 250566 345218 250608 345454
rect 250288 345134 250608 345218
rect 250288 344898 250330 345134
rect 250566 344898 250608 345134
rect 250288 344866 250608 344898
rect 281008 345454 281328 345486
rect 281008 345218 281050 345454
rect 281286 345218 281328 345454
rect 281008 345134 281328 345218
rect 281008 344898 281050 345134
rect 281286 344898 281328 345134
rect 281008 344866 281328 344898
rect 311728 345454 312048 345486
rect 311728 345218 311770 345454
rect 312006 345218 312048 345454
rect 311728 345134 312048 345218
rect 311728 344898 311770 345134
rect 312006 344898 312048 345134
rect 311728 344866 312048 344898
rect 199331 339420 199397 339421
rect 199331 339356 199332 339420
rect 199396 339356 199397 339420
rect 199331 339355 199397 339356
rect 204208 327454 204528 327486
rect 204208 327218 204250 327454
rect 204486 327218 204528 327454
rect 204208 327134 204528 327218
rect 204208 326898 204250 327134
rect 204486 326898 204528 327134
rect 204208 326866 204528 326898
rect 234928 327454 235248 327486
rect 234928 327218 234970 327454
rect 235206 327218 235248 327454
rect 234928 327134 235248 327218
rect 234928 326898 234970 327134
rect 235206 326898 235248 327134
rect 234928 326866 235248 326898
rect 265648 327454 265968 327486
rect 265648 327218 265690 327454
rect 265926 327218 265968 327454
rect 265648 327134 265968 327218
rect 265648 326898 265690 327134
rect 265926 326898 265968 327134
rect 265648 326866 265968 326898
rect 296368 327454 296688 327486
rect 296368 327218 296410 327454
rect 296646 327218 296688 327454
rect 296368 327134 296688 327218
rect 296368 326898 296410 327134
rect 296646 326898 296688 327134
rect 296368 326866 296688 326898
rect 219568 309454 219888 309486
rect 219568 309218 219610 309454
rect 219846 309218 219888 309454
rect 219568 309134 219888 309218
rect 219568 308898 219610 309134
rect 219846 308898 219888 309134
rect 219568 308866 219888 308898
rect 250288 309454 250608 309486
rect 250288 309218 250330 309454
rect 250566 309218 250608 309454
rect 250288 309134 250608 309218
rect 250288 308898 250330 309134
rect 250566 308898 250608 309134
rect 250288 308866 250608 308898
rect 281008 309454 281328 309486
rect 281008 309218 281050 309454
rect 281286 309218 281328 309454
rect 281008 309134 281328 309218
rect 281008 308898 281050 309134
rect 281286 308898 281328 309134
rect 281008 308866 281328 308898
rect 311728 309454 312048 309486
rect 311728 309218 311770 309454
rect 312006 309218 312048 309454
rect 311728 309134 312048 309218
rect 311728 308898 311770 309134
rect 312006 308898 312048 309134
rect 311728 308866 312048 308898
rect 204208 291454 204528 291486
rect 204208 291218 204250 291454
rect 204486 291218 204528 291454
rect 204208 291134 204528 291218
rect 204208 290898 204250 291134
rect 204486 290898 204528 291134
rect 204208 290866 204528 290898
rect 234928 291454 235248 291486
rect 234928 291218 234970 291454
rect 235206 291218 235248 291454
rect 234928 291134 235248 291218
rect 234928 290898 234970 291134
rect 235206 290898 235248 291134
rect 234928 290866 235248 290898
rect 265648 291454 265968 291486
rect 265648 291218 265690 291454
rect 265926 291218 265968 291454
rect 265648 291134 265968 291218
rect 265648 290898 265690 291134
rect 265926 290898 265968 291134
rect 265648 290866 265968 290898
rect 296368 291454 296688 291486
rect 296368 291218 296410 291454
rect 296646 291218 296688 291454
rect 296368 291134 296688 291218
rect 296368 290898 296410 291134
rect 296646 290898 296688 291134
rect 296368 290866 296688 290898
rect 219568 273454 219888 273486
rect 219568 273218 219610 273454
rect 219846 273218 219888 273454
rect 219568 273134 219888 273218
rect 219568 272898 219610 273134
rect 219846 272898 219888 273134
rect 219568 272866 219888 272898
rect 250288 273454 250608 273486
rect 250288 273218 250330 273454
rect 250566 273218 250608 273454
rect 250288 273134 250608 273218
rect 250288 272898 250330 273134
rect 250566 272898 250608 273134
rect 250288 272866 250608 272898
rect 281008 273454 281328 273486
rect 281008 273218 281050 273454
rect 281286 273218 281328 273454
rect 281008 273134 281328 273218
rect 281008 272898 281050 273134
rect 281286 272898 281328 273134
rect 281008 272866 281328 272898
rect 311728 273454 312048 273486
rect 311728 273218 311770 273454
rect 312006 273218 312048 273454
rect 311728 273134 312048 273218
rect 311728 272898 311770 273134
rect 312006 272898 312048 273134
rect 311728 272866 312048 272898
rect 204208 255454 204528 255486
rect 204208 255218 204250 255454
rect 204486 255218 204528 255454
rect 204208 255134 204528 255218
rect 204208 254898 204250 255134
rect 204486 254898 204528 255134
rect 204208 254866 204528 254898
rect 234928 255454 235248 255486
rect 234928 255218 234970 255454
rect 235206 255218 235248 255454
rect 234928 255134 235248 255218
rect 234928 254898 234970 255134
rect 235206 254898 235248 255134
rect 234928 254866 235248 254898
rect 265648 255454 265968 255486
rect 265648 255218 265690 255454
rect 265926 255218 265968 255454
rect 265648 255134 265968 255218
rect 265648 254898 265690 255134
rect 265926 254898 265968 255134
rect 265648 254866 265968 254898
rect 296368 255454 296688 255486
rect 296368 255218 296410 255454
rect 296646 255218 296688 255454
rect 296368 255134 296688 255218
rect 296368 254898 296410 255134
rect 296646 254898 296688 255134
rect 296368 254866 296688 254898
rect 319299 253060 319365 253061
rect 319299 252996 319300 253060
rect 319364 252996 319365 253060
rect 319299 252995 319365 252996
rect 200619 240820 200685 240821
rect 200619 240756 200620 240820
rect 200684 240756 200685 240820
rect 200619 240755 200685 240756
rect 199794 237454 200414 238000
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 198595 228988 198661 228989
rect 198595 228924 198596 228988
rect 198660 228924 198661 228988
rect 198595 228923 198661 228924
rect 198598 228309 198658 228923
rect 198595 228308 198661 228309
rect 198595 228244 198596 228308
rect 198660 228244 198661 228308
rect 198595 228243 198661 228244
rect 197123 211852 197189 211853
rect 197123 211788 197124 211852
rect 197188 211788 197189 211852
rect 197123 211787 197189 211788
rect 199794 201454 200414 236898
rect 200622 234293 200682 240755
rect 319302 238770 319362 252995
rect 318750 238710 319362 238770
rect 200619 234292 200685 234293
rect 200619 234228 200620 234292
rect 200684 234228 200685 234292
rect 200619 234227 200685 234228
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 195099 3364 195165 3365
rect 195099 3300 195100 3364
rect 195164 3300 195165 3364
rect 195099 3299 195165 3300
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 205174 204134 238000
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 208894 207854 238000
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 212614 211574 238000
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 219454 218414 238000
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 223174 222134 238000
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 226894 225854 238000
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 228954 230614 229574 238000
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 178000 229574 194058
rect 235794 237454 236414 238000
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 178000 236414 200898
rect 239514 205174 240134 238000
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 178000 240134 204618
rect 243234 208894 243854 238000
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 178000 243854 208338
rect 246954 212614 247574 238000
rect 252507 226948 252573 226949
rect 252507 226884 252508 226948
rect 252572 226884 252573 226948
rect 252507 226883 252573 226884
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 178000 247574 212058
rect 249379 186964 249445 186965
rect 249379 186900 249380 186964
rect 249444 186900 249445 186964
rect 249379 186899 249445 186900
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 249195 175948 249261 175949
rect 249195 175884 249196 175948
rect 249260 175884 249261 175948
rect 249195 175883 249261 175884
rect 249198 173365 249258 175883
rect 249382 174317 249442 186899
rect 249379 174316 249445 174317
rect 249379 174252 249380 174316
rect 249444 174252 249445 174316
rect 249379 174251 249445 174252
rect 249195 173364 249261 173365
rect 249195 173300 249196 173364
rect 249260 173300 249261 173364
rect 249195 173299 249261 173300
rect 227874 165454 228194 165486
rect 227874 165218 227916 165454
rect 228152 165218 228194 165454
rect 227874 165134 228194 165218
rect 227874 164898 227916 165134
rect 228152 164898 228194 165134
rect 227874 164866 228194 164898
rect 237805 165454 238125 165486
rect 237805 165218 237847 165454
rect 238083 165218 238125 165454
rect 237805 165134 238125 165218
rect 237805 164898 237847 165134
rect 238083 164898 238125 165134
rect 237805 164866 238125 164898
rect 252510 158813 252570 226883
rect 253794 219454 254414 238000
rect 255267 236604 255333 236605
rect 255267 236540 255268 236604
rect 255332 236540 255333 236604
rect 255267 236539 255333 236540
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 252507 158812 252573 158813
rect 252507 158748 252508 158812
rect 252572 158748 252573 158812
rect 252507 158747 252573 158748
rect 251771 149700 251837 149701
rect 251771 149636 251772 149700
rect 251836 149636 251837 149700
rect 251771 149635 251837 149636
rect 222910 147454 223230 147486
rect 222910 147218 222952 147454
rect 223188 147218 223230 147454
rect 222910 147134 223230 147218
rect 222910 146898 222952 147134
rect 223188 146898 223230 147134
rect 222910 146866 223230 146898
rect 232840 147454 233160 147486
rect 232840 147218 232882 147454
rect 233118 147218 233160 147454
rect 232840 147134 233160 147218
rect 232840 146898 232882 147134
rect 233118 146898 233160 147134
rect 232840 146866 233160 146898
rect 242771 147454 243091 147486
rect 242771 147218 242813 147454
rect 243049 147218 243091 147454
rect 242771 147134 243091 147218
rect 242771 146898 242813 147134
rect 243049 146898 243091 147134
rect 242771 146866 243091 146898
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 250299 134196 250365 134197
rect 250299 134132 250300 134196
rect 250364 134132 250365 134196
rect 250299 134131 250365 134132
rect 227874 129454 228194 129486
rect 227874 129218 227916 129454
rect 228152 129218 228194 129454
rect 227874 129134 228194 129218
rect 227874 128898 227916 129134
rect 228152 128898 228194 129134
rect 227874 128866 228194 128898
rect 237805 129454 238125 129486
rect 237805 129218 237847 129454
rect 238083 129218 238125 129454
rect 237805 129134 238125 129218
rect 237805 128898 237847 129134
rect 238083 128898 238125 129134
rect 237805 128866 238125 128898
rect 222910 111454 223230 111486
rect 222910 111218 222952 111454
rect 223188 111218 223230 111454
rect 222910 111134 223230 111218
rect 222910 110898 222952 111134
rect 223188 110898 223230 111134
rect 222910 110866 223230 110898
rect 232840 111454 233160 111486
rect 232840 111218 232882 111454
rect 233118 111218 233160 111454
rect 232840 111134 233160 111218
rect 232840 110898 232882 111134
rect 233118 110898 233160 111134
rect 232840 110866 233160 110898
rect 242771 111454 243091 111486
rect 242771 111218 242813 111454
rect 243049 111218 243091 111454
rect 242771 111134 243091 111218
rect 242771 110898 242813 111134
rect 243049 110898 243091 111134
rect 242771 110866 243091 110898
rect 214603 105228 214669 105229
rect 214603 105164 214604 105228
rect 214668 105164 214669 105228
rect 214603 105163 214669 105164
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 214419 103868 214485 103869
rect 214419 103804 214420 103868
rect 214484 103804 214485 103868
rect 214419 103803 214485 103804
rect 214422 91085 214482 103803
rect 214606 94893 214666 105163
rect 249195 97068 249261 97069
rect 249195 97004 249196 97068
rect 249260 97004 249261 97068
rect 249195 97003 249261 97004
rect 214603 94892 214669 94893
rect 214603 94828 214604 94892
rect 214668 94828 214669 94892
rect 214603 94827 214669 94828
rect 214419 91084 214485 91085
rect 214419 91020 214420 91084
rect 214484 91020 214485 91084
rect 214419 91019 214485 91020
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 93454 236414 94000
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 61174 240134 94000
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 64894 243854 94000
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 68614 247574 94000
rect 249198 84210 249258 97003
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 248462 84150 249258 84210
rect 248462 16557 248522 84150
rect 250302 26893 250362 134131
rect 251774 114477 251834 149635
rect 253794 147454 254414 182898
rect 254531 148340 254597 148341
rect 254531 148276 254532 148340
rect 254596 148276 254597 148340
rect 254531 148275 254597 148276
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253611 137188 253677 137189
rect 253611 137124 253612 137188
rect 253676 137124 253677 137188
rect 253611 137123 253677 137124
rect 251955 123316 252021 123317
rect 251955 123252 251956 123316
rect 252020 123252 252021 123316
rect 251955 123251 252021 123252
rect 251771 114476 251837 114477
rect 251771 114412 251772 114476
rect 251836 114412 251837 114476
rect 251771 114411 251837 114412
rect 251958 97069 252018 123251
rect 253614 122850 253674 137123
rect 253062 122790 253674 122850
rect 251955 97068 252021 97069
rect 251955 97004 251956 97068
rect 252020 97004 252021 97068
rect 251955 97003 252021 97004
rect 250299 26892 250365 26893
rect 250299 26828 250300 26892
rect 250364 26828 250365 26892
rect 250299 26827 250365 26828
rect 253062 25533 253122 122790
rect 253794 111454 254414 146898
rect 254534 146029 254594 148275
rect 255270 147933 255330 236539
rect 257514 223174 258134 238000
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 261234 226894 261854 238000
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 259499 199340 259565 199341
rect 259499 199276 259500 199340
rect 259564 199276 259565 199340
rect 259499 199275 259565 199276
rect 258579 192676 258645 192677
rect 258579 192612 258580 192676
rect 258644 192612 258645 192676
rect 258579 192611 258645 192612
rect 258395 192540 258461 192541
rect 258395 192476 258396 192540
rect 258460 192476 258461 192540
rect 258395 192475 258461 192476
rect 258398 190470 258458 192475
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 255451 178940 255517 178941
rect 255451 178876 255452 178940
rect 255516 178876 255517 178940
rect 255451 178875 255517 178876
rect 255267 147932 255333 147933
rect 255267 147868 255268 147932
rect 255332 147868 255333 147932
rect 255267 147867 255333 147868
rect 254531 146028 254597 146029
rect 254531 145964 254532 146028
rect 254596 145964 254597 146028
rect 254531 145963 254597 145964
rect 255454 140453 255514 178875
rect 256739 178804 256805 178805
rect 256739 178740 256740 178804
rect 256804 178740 256805 178804
rect 256739 178739 256805 178740
rect 256742 161125 256802 178739
rect 256739 161124 256805 161125
rect 256739 161060 256740 161124
rect 256804 161060 256805 161124
rect 256739 161059 256805 161060
rect 257514 151174 258134 186618
rect 258214 190410 258458 190470
rect 258214 151830 258274 190410
rect 258582 180810 258642 192611
rect 258398 180750 258642 180810
rect 258398 168469 258458 180750
rect 258395 168468 258461 168469
rect 258395 168404 258396 168468
rect 258460 168404 258461 168468
rect 258395 168403 258461 168404
rect 258214 151770 258458 151830
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 255451 140452 255517 140453
rect 255451 140388 255452 140452
rect 255516 140388 255517 140452
rect 255451 140387 255517 140388
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253059 25532 253125 25533
rect 253059 25468 253060 25532
rect 253124 25468 253125 25532
rect 253059 25467 253125 25468
rect 248459 16556 248525 16557
rect 248459 16492 248460 16556
rect 248524 16492 248525 16556
rect 248459 16491 248525 16492
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 115174 258134 150618
rect 258398 140997 258458 151770
rect 259502 144397 259562 199275
rect 261234 190894 261854 226338
rect 264954 230614 265574 238000
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 263547 210356 263613 210357
rect 263547 210292 263548 210356
rect 263612 210292 263613 210356
rect 263547 210291 263613 210292
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 259683 189684 259749 189685
rect 259683 189620 259684 189684
rect 259748 189620 259749 189684
rect 259683 189619 259749 189620
rect 259499 144396 259565 144397
rect 259499 144332 259500 144396
rect 259564 144332 259565 144396
rect 259499 144331 259565 144332
rect 259686 141133 259746 189619
rect 260971 180164 261037 180165
rect 260971 180100 260972 180164
rect 261036 180100 261037 180164
rect 260971 180099 261037 180100
rect 260974 167381 261034 180099
rect 260971 167380 261037 167381
rect 260971 167316 260972 167380
rect 261036 167316 261037 167380
rect 260971 167315 261037 167316
rect 261234 154894 261854 190338
rect 262259 185604 262325 185605
rect 262259 185540 262260 185604
rect 262324 185540 262325 185604
rect 262259 185539 262325 185540
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 259683 141132 259749 141133
rect 259683 141068 259684 141132
rect 259748 141068 259749 141132
rect 259683 141067 259749 141068
rect 258395 140996 258461 140997
rect 258395 140932 258396 140996
rect 258460 140932 258461 140996
rect 258395 140931 258461 140932
rect 260051 130116 260117 130117
rect 260051 130052 260052 130116
rect 260116 130052 260117 130116
rect 260051 130051 260117 130052
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 260054 61573 260114 130051
rect 261234 118894 261854 154338
rect 262262 138685 262322 185539
rect 262443 178668 262509 178669
rect 262443 178604 262444 178668
rect 262508 178604 262509 178668
rect 262443 178603 262509 178604
rect 262446 163165 262506 178603
rect 262443 163164 262509 163165
rect 262443 163100 262444 163164
rect 262508 163100 262509 163164
rect 262443 163099 262509 163100
rect 262259 138684 262325 138685
rect 262259 138620 262260 138684
rect 262324 138620 262325 138684
rect 262259 138619 262325 138620
rect 263550 137053 263610 210291
rect 263731 200700 263797 200701
rect 263731 200636 263732 200700
rect 263796 200636 263797 200700
rect 263731 200635 263797 200636
rect 263734 142221 263794 200635
rect 264954 194614 265574 230058
rect 271794 237454 272414 238000
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271091 222868 271157 222869
rect 271091 222804 271092 222868
rect 271156 222804 271157 222868
rect 271091 222803 271157 222804
rect 268331 210492 268397 210493
rect 268331 210428 268332 210492
rect 268396 210428 268397 210492
rect 268331 210427 268397 210428
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 266307 188324 266373 188325
rect 266307 188260 266308 188324
rect 266372 188260 266373 188324
rect 266307 188259 266373 188260
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 263731 142220 263797 142221
rect 263731 142156 263732 142220
rect 263796 142156 263797 142220
rect 263731 142155 263797 142156
rect 263547 137052 263613 137053
rect 263547 136988 263548 137052
rect 263612 136988 263613 137052
rect 263547 136987 263613 136988
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 260051 61572 260117 61573
rect 260051 61508 260052 61572
rect 260116 61508 260117 61572
rect 260051 61507 260117 61508
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 122614 265574 158058
rect 266310 153509 266370 188259
rect 266307 153508 266373 153509
rect 266307 153444 266308 153508
rect 266372 153444 266373 153508
rect 266307 153443 266373 153444
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 268334 44845 268394 210427
rect 269067 180028 269133 180029
rect 269067 179964 269068 180028
rect 269132 179964 269133 180028
rect 269067 179963 269133 179964
rect 269070 136917 269130 179963
rect 269067 136916 269133 136917
rect 269067 136852 269068 136916
rect 269132 136852 269133 136916
rect 269067 136851 269133 136852
rect 271094 61573 271154 222803
rect 271794 201454 272414 236898
rect 275514 205174 276134 238000
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 273851 204916 273917 204917
rect 273851 204852 273852 204916
rect 273916 204852 273917 204916
rect 273851 204851 273917 204852
rect 275514 204854 276134 204938
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271091 61572 271157 61573
rect 271091 61508 271092 61572
rect 271156 61508 271157 61572
rect 271091 61507 271157 61508
rect 271794 57454 272414 92898
rect 273854 76669 273914 204851
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 273851 76668 273917 76669
rect 273851 76604 273852 76668
rect 273916 76604 273917 76668
rect 273851 76603 273917 76604
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 268331 44844 268397 44845
rect 268331 44780 268332 44844
rect 268396 44780 268397 44844
rect 268331 44779 268397 44780
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 208894 279854 238000
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 212614 283574 238000
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 219454 290414 238000
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 223174 294134 238000
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 226894 297854 238000
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 230614 301574 238000
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 307794 237454 308414 238000
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 178000 308414 200898
rect 311514 205174 312134 238000
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 178000 312134 204618
rect 315234 208894 315854 238000
rect 318750 231709 318810 238710
rect 318747 231708 318813 231709
rect 318747 231644 318748 231708
rect 318812 231644 318813 231708
rect 318747 231643 318813 231644
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 178000 315854 208338
rect 318954 212614 319574 238000
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 178000 319574 212058
rect 320222 175813 320282 360435
rect 321507 359140 321573 359141
rect 321507 359076 321508 359140
rect 321572 359076 321573 359140
rect 321507 359075 321573 359076
rect 321323 184244 321389 184245
rect 321323 184180 321324 184244
rect 321388 184180 321389 184244
rect 321323 184179 321389 184180
rect 320219 175812 320285 175813
rect 320219 175748 320220 175812
rect 320284 175748 320285 175812
rect 320219 175747 320285 175748
rect 306971 175676 307037 175677
rect 306971 175612 306972 175676
rect 307036 175612 307037 175676
rect 306971 175611 307037 175612
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 306974 145621 307034 175611
rect 321326 170645 321386 184179
rect 321323 170644 321389 170645
rect 321323 170580 321324 170644
rect 321388 170580 321389 170644
rect 321323 170579 321389 170580
rect 314208 165454 314528 165486
rect 314208 165218 314250 165454
rect 314486 165218 314528 165454
rect 314208 165134 314528 165218
rect 314208 164898 314250 165134
rect 314486 164898 314528 165134
rect 314208 164866 314528 164898
rect 317472 165454 317792 165486
rect 317472 165218 317514 165454
rect 317750 165218 317792 165454
rect 317472 165134 317792 165218
rect 317472 164898 317514 165134
rect 317750 164898 317792 165134
rect 317472 164866 317792 164898
rect 312576 147454 312896 147486
rect 312576 147218 312618 147454
rect 312854 147218 312896 147454
rect 312576 147134 312896 147218
rect 312576 146898 312618 147134
rect 312854 146898 312896 147134
rect 312576 146866 312896 146898
rect 315840 147454 316160 147486
rect 315840 147218 315882 147454
rect 316118 147218 316160 147454
rect 315840 147134 316160 147218
rect 315840 146898 315882 147134
rect 316118 146898 316160 147134
rect 315840 146866 316160 146898
rect 319104 147454 319424 147486
rect 319104 147218 319146 147454
rect 319382 147218 319424 147454
rect 319104 147134 319424 147218
rect 319104 146898 319146 147134
rect 319382 146898 319424 147134
rect 319104 146866 319424 146898
rect 306971 145620 307037 145621
rect 306971 145556 306972 145620
rect 307036 145556 307037 145620
rect 306971 145555 307037 145556
rect 307707 145076 307773 145077
rect 307707 145012 307708 145076
rect 307772 145012 307773 145076
rect 307707 145011 307773 145012
rect 307710 143989 307770 145011
rect 307707 143988 307773 143989
rect 307707 143924 307708 143988
rect 307772 143924 307773 143988
rect 307707 143923 307773 143924
rect 321510 132157 321570 359075
rect 324270 311813 324330 371315
rect 325794 363454 326414 398898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 331259 406332 331325 406333
rect 331259 406268 331260 406332
rect 331324 406268 331325 406332
rect 331259 406267 331325 406268
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 326659 365804 326725 365805
rect 326659 365740 326660 365804
rect 326724 365740 326725 365804
rect 326659 365739 326725 365740
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 324267 311812 324333 311813
rect 324267 311748 324268 311812
rect 324332 311748 324333 311812
rect 324267 311747 324333 311748
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 324267 258364 324333 258365
rect 324267 258300 324268 258364
rect 324332 258300 324333 258364
rect 324267 258299 324333 258300
rect 324270 230485 324330 258299
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 324267 230484 324333 230485
rect 324267 230420 324268 230484
rect 324332 230420 324333 230484
rect 324267 230419 324333 230420
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 321691 177444 321757 177445
rect 321691 177380 321692 177444
rect 321756 177380 321757 177444
rect 321691 177379 321757 177380
rect 321694 166837 321754 177379
rect 321691 166836 321757 166837
rect 321691 166772 321692 166836
rect 321756 166772 321757 166836
rect 321691 166771 321757 166772
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 321507 132156 321573 132157
rect 321507 132092 321508 132156
rect 321572 132092 321573 132156
rect 321507 132091 321573 132092
rect 314208 129454 314528 129486
rect 314208 129218 314250 129454
rect 314486 129218 314528 129454
rect 314208 129134 314528 129218
rect 314208 128898 314250 129134
rect 314486 128898 314528 129134
rect 314208 128866 314528 128898
rect 317472 129454 317792 129486
rect 317472 129218 317514 129454
rect 317750 129218 317792 129454
rect 317472 129134 317792 129218
rect 317472 128898 317514 129134
rect 317750 128898 317792 129134
rect 317472 128866 317792 128898
rect 307155 127668 307221 127669
rect 307155 127604 307156 127668
rect 307220 127604 307221 127668
rect 307155 127603 307221 127604
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 302739 118148 302805 118149
rect 302739 118084 302740 118148
rect 302804 118084 302805 118148
rect 302739 118083 302805 118084
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 302742 57221 302802 118083
rect 305499 102916 305565 102917
rect 305499 102852 305500 102916
rect 305564 102852 305565 102916
rect 305499 102851 305565 102852
rect 304211 96932 304277 96933
rect 304211 96868 304212 96932
rect 304276 96868 304277 96932
rect 304211 96867 304277 96868
rect 304214 76533 304274 96867
rect 304763 77892 304829 77893
rect 304763 77828 304764 77892
rect 304828 77828 304829 77892
rect 304763 77827 304829 77828
rect 304211 76532 304277 76533
rect 304211 76468 304212 76532
rect 304276 76468 304277 76532
rect 304211 76467 304277 76468
rect 302739 57220 302805 57221
rect 302739 57156 302740 57220
rect 302804 57156 302805 57220
rect 302739 57155 302805 57156
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 304766 3501 304826 77827
rect 305502 13021 305562 102851
rect 306971 96796 307037 96797
rect 306971 96732 306972 96796
rect 307036 96732 307037 96796
rect 306971 96731 307037 96732
rect 306974 51781 307034 96731
rect 307158 82109 307218 127603
rect 312576 111454 312896 111486
rect 312576 111218 312618 111454
rect 312854 111218 312896 111454
rect 312576 111134 312896 111218
rect 312576 110898 312618 111134
rect 312854 110898 312896 111134
rect 312576 110866 312896 110898
rect 315840 111454 316160 111486
rect 315840 111218 315882 111454
rect 316118 111218 316160 111454
rect 315840 111134 316160 111218
rect 315840 110898 315882 111134
rect 316118 110898 316160 111134
rect 315840 110866 316160 110898
rect 319104 111454 319424 111486
rect 319104 111218 319146 111454
rect 319382 111218 319424 111454
rect 319104 111134 319424 111218
rect 319104 110898 319146 111134
rect 319382 110898 319424 111134
rect 319104 110866 319424 110898
rect 325794 111454 326414 146898
rect 326662 140181 326722 365739
rect 328499 363084 328565 363085
rect 328499 363020 328500 363084
rect 328564 363020 328565 363084
rect 328499 363019 328565 363020
rect 327027 353428 327093 353429
rect 327027 353364 327028 353428
rect 327092 353364 327093 353428
rect 327027 353363 327093 353364
rect 326659 140180 326725 140181
rect 326659 140116 326660 140180
rect 326724 140116 326725 140180
rect 326659 140115 326725 140116
rect 327030 139365 327090 353363
rect 327211 240004 327277 240005
rect 327211 239940 327212 240004
rect 327276 239940 327277 240004
rect 327211 239939 327277 239940
rect 327214 143989 327274 239939
rect 327211 143988 327277 143989
rect 327211 143924 327212 143988
rect 327276 143924 327277 143988
rect 327211 143923 327277 143924
rect 327027 139364 327093 139365
rect 327027 139300 327028 139364
rect 327092 139300 327093 139364
rect 327027 139299 327093 139300
rect 328502 134061 328562 363019
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 330339 240140 330405 240141
rect 330339 240076 330340 240140
rect 330404 240076 330405 240140
rect 330339 240075 330405 240076
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 330342 154869 330402 240075
rect 330339 154868 330405 154869
rect 330339 154804 330340 154868
rect 330404 154804 330405 154868
rect 330339 154803 330405 154804
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 328499 134060 328565 134061
rect 328499 133996 328500 134060
rect 328564 133996 328565 134060
rect 328499 133995 328565 133996
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 324267 98564 324333 98565
rect 324267 98500 324268 98564
rect 324332 98500 324333 98564
rect 324267 98499 324333 98500
rect 307794 93454 308414 94000
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307155 82108 307221 82109
rect 307155 82044 307156 82108
rect 307220 82044 307221 82108
rect 307155 82043 307221 82044
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 306971 51780 307037 51781
rect 306971 51716 306972 51780
rect 307036 51716 307037 51780
rect 306971 51715 307037 51716
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 305499 13020 305565 13021
rect 305499 12956 305500 13020
rect 305564 12956 305565 13020
rect 305499 12955 305565 12956
rect 304763 3500 304829 3501
rect 304763 3436 304764 3500
rect 304828 3436 304829 3500
rect 304763 3435 304829 3436
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 61174 312134 94000
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 64894 315854 94000
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 68614 319574 94000
rect 324270 93805 324330 98499
rect 324267 93804 324333 93805
rect 324267 93740 324268 93804
rect 324332 93740 324333 93804
rect 324267 93739 324333 93740
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 115174 330134 150618
rect 331262 147797 331322 406267
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 332547 364444 332613 364445
rect 332547 364380 332548 364444
rect 332612 364380 332613 364444
rect 332547 364379 332613 364380
rect 331443 181524 331509 181525
rect 331443 181460 331444 181524
rect 331508 181460 331509 181524
rect 331443 181459 331509 181460
rect 331446 171189 331506 181459
rect 331443 171188 331509 171189
rect 331443 171124 331444 171188
rect 331508 171124 331509 171188
rect 331443 171123 331509 171124
rect 331259 147796 331325 147797
rect 331259 147732 331260 147796
rect 331324 147732 331325 147796
rect 331259 147731 331325 147732
rect 332550 133925 332610 364379
rect 333234 334894 333854 370338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 338251 407148 338317 407149
rect 338251 407084 338252 407148
rect 338316 407084 338317 407148
rect 338251 407083 338317 407084
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 334019 363220 334085 363221
rect 334019 363156 334020 363220
rect 334084 363156 334085 363220
rect 334019 363155 334085 363156
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 334022 156501 334082 363155
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 335859 215932 335925 215933
rect 335859 215868 335860 215932
rect 335924 215868 335925 215932
rect 335859 215867 335925 215868
rect 334571 172548 334637 172549
rect 334571 172484 334572 172548
rect 334636 172484 334637 172548
rect 334571 172483 334637 172484
rect 334019 156500 334085 156501
rect 334019 156436 334020 156500
rect 334084 156436 334085 156500
rect 334019 156435 334085 156436
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 332547 133924 332613 133925
rect 332547 133860 332548 133924
rect 332612 133860 332613 133924
rect 332547 133859 332613 133860
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 334574 82245 334634 172483
rect 335862 96389 335922 215867
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336043 169828 336109 169829
rect 336043 169764 336044 169828
rect 336108 169764 336109 169828
rect 336043 169763 336109 169764
rect 335859 96388 335925 96389
rect 335859 96324 335860 96388
rect 335924 96324 335925 96388
rect 335859 96323 335925 96324
rect 334571 82244 334637 82245
rect 334571 82180 334572 82244
rect 334636 82180 334637 82244
rect 334571 82179 334637 82180
rect 336046 62117 336106 169763
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336043 62116 336109 62117
rect 336043 62052 336044 62116
rect 336108 62052 336109 62116
rect 336043 62051 336109 62052
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 86058
rect 338254 77893 338314 407083
rect 342299 404428 342365 404429
rect 342299 404364 342300 404428
rect 342364 404364 342365 404428
rect 342299 404363 342365 404364
rect 339539 401708 339605 401709
rect 339539 401644 339540 401708
rect 339604 401644 339605 401708
rect 339539 401643 339605 401644
rect 338619 157452 338685 157453
rect 338619 157388 338620 157452
rect 338684 157388 338685 157452
rect 338619 157387 338685 157388
rect 338251 77892 338317 77893
rect 338251 77828 338252 77892
rect 338316 77828 338317 77892
rect 338251 77827 338317 77828
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 338622 46885 338682 157387
rect 338619 46884 338685 46885
rect 338619 46820 338620 46884
rect 338684 46820 338685 46884
rect 338619 46819 338685 46820
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 339542 8261 339602 401643
rect 340827 385660 340893 385661
rect 340827 385596 340828 385660
rect 340892 385596 340893 385660
rect 340827 385595 340893 385596
rect 340830 47565 340890 385595
rect 340827 47564 340893 47565
rect 340827 47500 340828 47564
rect 340892 47500 340893 47564
rect 340827 47499 340893 47500
rect 340830 11797 340890 47499
rect 342302 41309 342362 404363
rect 343794 381454 344414 416898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 345059 397492 345125 397493
rect 345059 397428 345060 397492
rect 345124 397428 345125 397492
rect 345059 397427 345125 397428
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 345062 81429 345122 397427
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 349107 379540 349173 379541
rect 349107 379476 349108 379540
rect 349172 379476 349173 379540
rect 349107 379475 349173 379476
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 349110 167109 349170 379475
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 349107 167108 349173 167109
rect 349107 167044 349108 167108
rect 349172 167044 349173 167108
rect 349107 167043 349173 167044
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 345059 81428 345125 81429
rect 345059 81364 345060 81428
rect 345124 81364 345125 81428
rect 345059 81363 345125 81364
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 342299 41308 342365 41309
rect 342299 41244 342300 41308
rect 342364 41244 342365 41308
rect 342299 41243 342365 41244
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 340827 11796 340893 11797
rect 340827 11732 340828 11796
rect 340892 11732 340893 11796
rect 340827 11731 340893 11732
rect 339539 8260 339605 8261
rect 339539 8196 339540 8260
rect 339604 8196 339605 8260
rect 339539 8195 339605 8196
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 181600 420134 204618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 181600 423854 208338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 181600 427574 212058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 181600 434414 182898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 181600 438134 186618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 181600 441854 190338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 181600 445574 194058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 181600 452414 200898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 181600 456134 204618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 181600 459854 208338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 181600 463574 212058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 181600 470414 182898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 181600 474134 186618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 181600 477854 190338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 181600 481574 194058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 181600 488414 200898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 494099 356692 494165 356693
rect 494099 356628 494100 356692
rect 494164 356628 494165 356692
rect 494099 356627 494165 356628
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 181600 492134 204618
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 439568 165454 439888 165486
rect 439568 165218 439610 165454
rect 439846 165218 439888 165454
rect 439568 165134 439888 165218
rect 439568 164898 439610 165134
rect 439846 164898 439888 165134
rect 439568 164866 439888 164898
rect 470288 165454 470608 165486
rect 470288 165218 470330 165454
rect 470566 165218 470608 165454
rect 470288 165134 470608 165218
rect 470288 164898 470330 165134
rect 470566 164898 470608 165134
rect 470288 164866 470608 164898
rect 424208 147454 424528 147486
rect 424208 147218 424250 147454
rect 424486 147218 424528 147454
rect 424208 147134 424528 147218
rect 424208 146898 424250 147134
rect 424486 146898 424528 147134
rect 424208 146866 424528 146898
rect 454928 147454 455248 147486
rect 454928 147218 454970 147454
rect 455206 147218 455248 147454
rect 454928 147134 455248 147218
rect 454928 146898 454970 147134
rect 455206 146898 455248 147134
rect 454928 146866 455248 146898
rect 485648 147454 485968 147486
rect 485648 147218 485690 147454
rect 485926 147218 485968 147454
rect 485648 147134 485968 147218
rect 485648 146898 485690 147134
rect 485926 146898 485968 147134
rect 485648 146866 485968 146898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 439568 129454 439888 129486
rect 439568 129218 439610 129454
rect 439846 129218 439888 129454
rect 439568 129134 439888 129218
rect 439568 128898 439610 129134
rect 439846 128898 439888 129134
rect 439568 128866 439888 128898
rect 470288 129454 470608 129486
rect 470288 129218 470330 129454
rect 470566 129218 470608 129454
rect 470288 129134 470608 129218
rect 470288 128898 470330 129134
rect 470566 128898 470608 129134
rect 494102 129029 494162 356627
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 181600 495854 208338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 503667 191044 503733 191045
rect 503667 190980 503668 191044
rect 503732 190980 503733 191044
rect 503667 190979 503733 190980
rect 502379 178668 502445 178669
rect 502379 178604 502380 178668
rect 502444 178604 502445 178668
rect 502379 178603 502445 178604
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 496859 174452 496925 174453
rect 496859 174388 496860 174452
rect 496924 174388 496925 174452
rect 496859 174387 496925 174388
rect 495939 172276 496005 172277
rect 495939 172212 495940 172276
rect 496004 172212 496005 172276
rect 495939 172211 496005 172212
rect 494283 169828 494349 169829
rect 494283 169764 494284 169828
rect 494348 169764 494349 169828
rect 494283 169763 494349 169764
rect 494099 129028 494165 129029
rect 494099 128964 494100 129028
rect 494164 128964 494165 129028
rect 494099 128963 494165 128964
rect 470288 128866 470608 128898
rect 424208 111454 424528 111486
rect 424208 111218 424250 111454
rect 424486 111218 424528 111454
rect 424208 111134 424528 111218
rect 424208 110898 424250 111134
rect 424486 110898 424528 111134
rect 424208 110866 424528 110898
rect 454928 111454 455248 111486
rect 454928 111218 454970 111454
rect 455206 111218 455248 111454
rect 454928 111134 455248 111218
rect 454928 110898 454970 111134
rect 455206 110898 455248 111134
rect 454928 110866 455248 110898
rect 485648 111454 485968 111486
rect 485648 111218 485690 111454
rect 485926 111218 485968 111454
rect 485648 111134 485968 111218
rect 485648 110898 485690 111134
rect 485926 110898 485968 111134
rect 485648 110866 485968 110898
rect 493915 102236 493981 102237
rect 493915 102172 493916 102236
rect 493980 102172 493981 102236
rect 493915 102171 493981 102172
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 97174 420134 98000
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 64894 423854 98000
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 68614 427574 98000
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 75454 434414 98000
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 79174 438134 98000
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 82894 441854 98000
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 86614 445574 98000
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 93454 452414 98000
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 97174 456134 98000
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 64894 459854 98000
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 68614 463574 98000
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 75454 470414 98000
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 79174 474134 98000
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 82894 477854 98000
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 86614 481574 98000
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 93454 488414 98000
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 97174 492134 98000
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 493918 95165 493978 102171
rect 494286 99381 494346 169763
rect 494283 99380 494349 99381
rect 494283 99316 494284 99380
rect 494348 99316 494349 99380
rect 494283 99315 494349 99316
rect 493915 95164 493981 95165
rect 493915 95100 493916 95164
rect 493980 95100 493981 95164
rect 493915 95099 493981 95100
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 64894 495854 98000
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495942 44845 496002 172211
rect 496862 46885 496922 174387
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 502382 133925 502442 178603
rect 503670 166973 503730 190979
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 503667 166972 503733 166973
rect 503667 166908 503668 166972
rect 503732 166908 503733 166972
rect 503667 166907 503733 166908
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 502379 133924 502445 133925
rect 502379 133860 502380 133924
rect 502444 133860 502445 133924
rect 502379 133859 502445 133860
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 496859 46884 496925 46885
rect 496859 46820 496860 46884
rect 496924 46820 496925 46884
rect 496859 46819 496925 46820
rect 495939 44844 496005 44845
rect 495939 44780 495940 44844
rect 496004 44780 496005 44844
rect 495939 44779 496005 44780
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 74250 651218 74486 651454
rect 74250 650898 74486 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 89610 669218 89846 669454
rect 89610 668898 89846 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 104970 651218 105206 651454
rect 104970 650898 105206 651134
rect 76618 579218 76854 579454
rect 76618 578898 76854 579134
rect 87882 579218 88118 579454
rect 87882 578898 88118 579134
rect 99146 579218 99382 579454
rect 99146 578898 99382 579134
rect 82250 561218 82486 561454
rect 82250 560898 82486 561134
rect 93514 561218 93750 561454
rect 93514 560898 93750 561134
rect 76618 543218 76854 543454
rect 76618 542898 76854 543134
rect 87882 543218 88118 543454
rect 87882 542898 88118 543134
rect 99146 543218 99382 543454
rect 99146 542898 99382 543134
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 75618 471218 75854 471454
rect 75618 470898 75854 471134
rect 84882 471218 85118 471454
rect 84882 470898 85118 471134
rect 94146 471218 94382 471454
rect 94146 470898 94382 471134
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 80250 453218 80486 453454
rect 80250 452898 80486 453134
rect 89514 453218 89750 453454
rect 89514 452898 89750 453134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 89610 381218 89846 381454
rect 89610 380898 89846 381134
rect 74250 363218 74486 363454
rect 74250 362898 74486 363134
rect 104970 363218 105206 363454
rect 104970 362898 105206 363134
rect 89610 345218 89846 345454
rect 89610 344898 89846 345134
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 89610 273218 89846 273454
rect 89610 272898 89846 273134
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 74250 255218 74486 255454
rect 74250 254898 74486 255134
rect 104970 255218 105206 255454
rect 104970 254898 105206 255134
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 219610 345218 219846 345454
rect 219610 344898 219846 345134
rect 250330 345218 250566 345454
rect 250330 344898 250566 345134
rect 281050 345218 281286 345454
rect 281050 344898 281286 345134
rect 311770 345218 312006 345454
rect 311770 344898 312006 345134
rect 204250 327218 204486 327454
rect 204250 326898 204486 327134
rect 234970 327218 235206 327454
rect 234970 326898 235206 327134
rect 265690 327218 265926 327454
rect 265690 326898 265926 327134
rect 296410 327218 296646 327454
rect 296410 326898 296646 327134
rect 219610 309218 219846 309454
rect 219610 308898 219846 309134
rect 250330 309218 250566 309454
rect 250330 308898 250566 309134
rect 281050 309218 281286 309454
rect 281050 308898 281286 309134
rect 311770 309218 312006 309454
rect 311770 308898 312006 309134
rect 204250 291218 204486 291454
rect 204250 290898 204486 291134
rect 234970 291218 235206 291454
rect 234970 290898 235206 291134
rect 265690 291218 265926 291454
rect 265690 290898 265926 291134
rect 296410 291218 296646 291454
rect 296410 290898 296646 291134
rect 219610 273218 219846 273454
rect 219610 272898 219846 273134
rect 250330 273218 250566 273454
rect 250330 272898 250566 273134
rect 281050 273218 281286 273454
rect 281050 272898 281286 273134
rect 311770 273218 312006 273454
rect 311770 272898 312006 273134
rect 204250 255218 204486 255454
rect 204250 254898 204486 255134
rect 234970 255218 235206 255454
rect 234970 254898 235206 255134
rect 265690 255218 265926 255454
rect 265690 254898 265926 255134
rect 296410 255218 296646 255454
rect 296410 254898 296646 255134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 227916 165218 228152 165454
rect 227916 164898 228152 165134
rect 237847 165218 238083 165454
rect 237847 164898 238083 165134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 222952 147218 223188 147454
rect 222952 146898 223188 147134
rect 232882 147218 233118 147454
rect 232882 146898 233118 147134
rect 242813 147218 243049 147454
rect 242813 146898 243049 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 227916 129218 228152 129454
rect 227916 128898 228152 129134
rect 237847 129218 238083 129454
rect 237847 128898 238083 129134
rect 222952 111218 223188 111454
rect 222952 110898 223188 111134
rect 232882 111218 233118 111454
rect 232882 110898 233118 111134
rect 242813 111218 243049 111454
rect 242813 110898 243049 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 314250 165218 314486 165454
rect 314250 164898 314486 165134
rect 317514 165218 317750 165454
rect 317514 164898 317750 165134
rect 312618 147218 312854 147454
rect 312618 146898 312854 147134
rect 315882 147218 316118 147454
rect 315882 146898 316118 147134
rect 319146 147218 319382 147454
rect 319146 146898 319382 147134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 314250 129218 314486 129454
rect 314250 128898 314486 129134
rect 317514 129218 317750 129454
rect 317514 128898 317750 129134
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 312618 111218 312854 111454
rect 312618 110898 312854 111134
rect 315882 111218 316118 111454
rect 315882 110898 316118 111134
rect 319146 111218 319382 111454
rect 319146 110898 319382 111134
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 439610 165218 439846 165454
rect 439610 164898 439846 165134
rect 470330 165218 470566 165454
rect 470330 164898 470566 165134
rect 424250 147218 424486 147454
rect 424250 146898 424486 147134
rect 454970 147218 455206 147454
rect 454970 146898 455206 147134
rect 485690 147218 485926 147454
rect 485690 146898 485926 147134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 439610 129218 439846 129454
rect 439610 128898 439846 129134
rect 470330 129218 470566 129454
rect 470330 128898 470566 129134
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 424250 111218 424486 111454
rect 424250 110898 424486 111134
rect 454970 111218 455206 111454
rect 454970 110898 455206 111134
rect 485690 111218 485926 111454
rect 485690 110898 485926 111134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 89610 669454
rect 89846 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 89610 669134
rect 89846 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 74250 651454
rect 74486 651218 104970 651454
rect 105206 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 74250 651134
rect 74486 650898 104970 651134
rect 105206 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 76618 579454
rect 76854 579218 87882 579454
rect 88118 579218 99146 579454
rect 99382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 76618 579134
rect 76854 578898 87882 579134
rect 88118 578898 99146 579134
rect 99382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 82250 561454
rect 82486 561218 93514 561454
rect 93750 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 82250 561134
rect 82486 560898 93514 561134
rect 93750 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 76618 543454
rect 76854 543218 87882 543454
rect 88118 543218 99146 543454
rect 99382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 76618 543134
rect 76854 542898 87882 543134
rect 88118 542898 99146 543134
rect 99382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 75618 471454
rect 75854 471218 84882 471454
rect 85118 471218 94146 471454
rect 94382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 75618 471134
rect 75854 470898 84882 471134
rect 85118 470898 94146 471134
rect 94382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 80250 453454
rect 80486 453218 89514 453454
rect 89750 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 80250 453134
rect 80486 452898 89514 453134
rect 89750 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 89610 381454
rect 89846 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 89610 381134
rect 89846 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 74250 363454
rect 74486 363218 104970 363454
rect 105206 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 74250 363134
rect 74486 362898 104970 363134
rect 105206 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 89610 345454
rect 89846 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 219610 345454
rect 219846 345218 250330 345454
rect 250566 345218 281050 345454
rect 281286 345218 311770 345454
rect 312006 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 89610 345134
rect 89846 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 219610 345134
rect 219846 344898 250330 345134
rect 250566 344898 281050 345134
rect 281286 344898 311770 345134
rect 312006 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 204250 327454
rect 204486 327218 234970 327454
rect 235206 327218 265690 327454
rect 265926 327218 296410 327454
rect 296646 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 204250 327134
rect 204486 326898 234970 327134
rect 235206 326898 265690 327134
rect 265926 326898 296410 327134
rect 296646 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 219610 309454
rect 219846 309218 250330 309454
rect 250566 309218 281050 309454
rect 281286 309218 311770 309454
rect 312006 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 219610 309134
rect 219846 308898 250330 309134
rect 250566 308898 281050 309134
rect 281286 308898 311770 309134
rect 312006 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 204250 291454
rect 204486 291218 234970 291454
rect 235206 291218 265690 291454
rect 265926 291218 296410 291454
rect 296646 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 204250 291134
rect 204486 290898 234970 291134
rect 235206 290898 265690 291134
rect 265926 290898 296410 291134
rect 296646 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 89610 273454
rect 89846 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219610 273454
rect 219846 273218 250330 273454
rect 250566 273218 281050 273454
rect 281286 273218 311770 273454
rect 312006 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 89610 273134
rect 89846 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219610 273134
rect 219846 272898 250330 273134
rect 250566 272898 281050 273134
rect 281286 272898 311770 273134
rect 312006 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 74250 255454
rect 74486 255218 104970 255454
rect 105206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204250 255454
rect 204486 255218 234970 255454
rect 235206 255218 265690 255454
rect 265926 255218 296410 255454
rect 296646 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 74250 255134
rect 74486 254898 104970 255134
rect 105206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204250 255134
rect 204486 254898 234970 255134
rect 235206 254898 265690 255134
rect 265926 254898 296410 255134
rect 296646 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 227916 165454
rect 228152 165218 237847 165454
rect 238083 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 314250 165454
rect 314486 165218 317514 165454
rect 317750 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 439610 165454
rect 439846 165218 470330 165454
rect 470566 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 227916 165134
rect 228152 164898 237847 165134
rect 238083 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 314250 165134
rect 314486 164898 317514 165134
rect 317750 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 439610 165134
rect 439846 164898 470330 165134
rect 470566 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 222952 147454
rect 223188 147218 232882 147454
rect 233118 147218 242813 147454
rect 243049 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 312618 147454
rect 312854 147218 315882 147454
rect 316118 147218 319146 147454
rect 319382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 424250 147454
rect 424486 147218 454970 147454
rect 455206 147218 485690 147454
rect 485926 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 222952 147134
rect 223188 146898 232882 147134
rect 233118 146898 242813 147134
rect 243049 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 312618 147134
rect 312854 146898 315882 147134
rect 316118 146898 319146 147134
rect 319382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 424250 147134
rect 424486 146898 454970 147134
rect 455206 146898 485690 147134
rect 485926 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 227916 129454
rect 228152 129218 237847 129454
rect 238083 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 314250 129454
rect 314486 129218 317514 129454
rect 317750 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 439610 129454
rect 439846 129218 470330 129454
rect 470566 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 227916 129134
rect 228152 128898 237847 129134
rect 238083 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 314250 129134
rect 314486 128898 317514 129134
rect 317750 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 439610 129134
rect 439846 128898 470330 129134
rect 470566 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 222952 111454
rect 223188 111218 232882 111454
rect 233118 111218 242813 111454
rect 243049 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 312618 111454
rect 312854 111218 315882 111454
rect 316118 111218 319146 111454
rect 319382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 424250 111454
rect 424486 111218 454970 111454
rect 455206 111218 485690 111454
rect 485926 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 222952 111134
rect 223188 110898 232882 111134
rect 233118 110898 242813 111134
rect 243049 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 312618 111134
rect 312854 110898 315882 111134
rect 316118 110898 319146 111134
rect 319382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 424250 111134
rect 424486 110898 454970 111134
rect 455206 110898 485690 111134
rect 485926 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 0
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
use wb_bridge_2way  wb_bridge_2way
timestamp 0
transform 1 0 310000 0 1 96000
box 0 144 12000 80000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 0
transform 1 0 217000 0 1 96000
box 0 144 32000 79688
use wrapped_alu74181  wrapped_alu74181_7
timestamp 0
transform 1 0 70000 0 1 640000
box -10 -52 40000 40000
use wrapped_frequency_counter  wrapped_frequency_counter_2
timestamp 0
transform 1 0 70000 0 1 440000
box -10 -52 30000 50000
use wrapped_function_generator  wrapped_function_generator_0
timestamp 0
transform 1 0 70000 0 1 240000
box 0 0 50000 52000
use wrapped_hack_soc_dffram  wrapped_hack_soc_dffram_11
timestamp 0
transform 1 0 420000 0 1 100000
box 0 0 74470 79600
use wrapped_rgb_mixer  wrapped_rgb_mixer_3
timestamp 0
transform 1 0 70000 0 1 540000
box -10 -52 36000 42000
use wrapped_teras  wrapped_teras_13
timestamp 0
transform 1 0 200000 0 1 240000
box -10 -52 120000 120000
use wrapped_vga_clock  wrapped_vga_clock_1
timestamp 0
transform 1 0 70000 0 1 340000
box -10 -52 46000 46000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 98000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 238000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 294000 74414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 294000 110414 338000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 388000 74414 438000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 492000 74414 538000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 584000 74414 638000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 388000 110414 638000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 682000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 682000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 362000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 362000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 362000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 181600 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 181600 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 98000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 238000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 294000 78134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 294000 114134 338000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 388000 78134 438000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 492000 78134 538000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 584000 78134 638000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 682000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 388000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 362000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 362000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 362000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 181600 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 181600 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 98000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 238000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 294000 81854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 294000 117854 338000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 388000 81854 438000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 492000 81854 538000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 584000 81854 638000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 682000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 388000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 362000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 362000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 362000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 181600 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 181600 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 98000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 238000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 294000 85574 338000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 388000 85574 438000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 492000 85574 538000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 584000 85574 638000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 682000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 294000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 362000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 362000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 362000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 181600 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 181600 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 98000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 178000 243854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 178000 315854 238000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 294000 99854 338000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 388000 99854 438000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 492000 99854 538000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 584000 99854 638000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 682000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 362000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 362000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 362000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 362000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 181600 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 181600 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 181600 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 94000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 98000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 178000 247574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 178000 319574 238000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 294000 103574 338000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 388000 103574 538000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 584000 103574 638000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 682000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 362000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 362000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 362000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 362000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 181600 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 181600 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 98000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 178000 236414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 178000 308414 238000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 294000 92414 338000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 388000 92414 438000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 492000 92414 538000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 584000 92414 638000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 682000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 362000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 362000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 362000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 362000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 181600 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 181600 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 98000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 178000 240134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 178000 312134 238000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 294000 96134 338000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 388000 96134 438000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 492000 96134 538000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 584000 96134 638000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 682000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 362000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 362000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 362000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 362000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 181600 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 181600 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 181600 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
